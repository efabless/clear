* NGSPICE file created from bottom_right_tile.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

.subckt bottom_right_tile VGND VPWR ccff_head ccff_head_1 ccff_tail ccff_tail_0 chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[20] chanx_left_in[21] chanx_left_in[22] chanx_left_in[23]
+ chanx_left_in[24] chanx_left_in[25] chanx_left_in[26] chanx_left_in[27] chanx_left_in[28]
+ chanx_left_in[29] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[20] chanx_left_out[21] chanx_left_out[22] chanx_left_out[23]
+ chanx_left_out[24] chanx_left_out[25] chanx_left_out[26] chanx_left_out[27] chanx_left_out[28]
+ chanx_left_out[29] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chany_top_in[0]
+ chany_top_in[10] chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14]
+ chany_top_in[15] chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19]
+ chany_top_in[1] chany_top_in[20] chany_top_in[21] chany_top_in[22] chany_top_in[23]
+ chany_top_in[24] chany_top_in[25] chany_top_in[26] chany_top_in[27] chany_top_in[28]
+ chany_top_in[29] chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5]
+ chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0]
+ chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14]
+ chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19]
+ chany_top_out[1] chany_top_out[20] chany_top_out[21] chany_top_out[22] chany_top_out[23]
+ chany_top_out[24] chany_top_out[25] chany_top_out[26] chany_top_out[27] chany_top_out[28]
+ chany_top_out[29] chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5]
+ chany_top_out[6] chany_top_out[7] chany_top_out[8] chany_top_out[9] gfpga_pad_io_soc_dir[0]
+ gfpga_pad_io_soc_dir[1] gfpga_pad_io_soc_dir[2] gfpga_pad_io_soc_dir[3] gfpga_pad_io_soc_in[0]
+ gfpga_pad_io_soc_in[1] gfpga_pad_io_soc_in[2] gfpga_pad_io_soc_in[3] gfpga_pad_io_soc_out[0]
+ gfpga_pad_io_soc_out[1] gfpga_pad_io_soc_out[2] gfpga_pad_io_soc_out[3] isol_n prog_clk
+ prog_reset reset test_enable top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
+ top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_ top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_ top_width_0_height_0_subtile_0__pin_inpad_0_
+ top_width_0_height_0_subtile_1__pin_inpad_0_ top_width_0_height_0_subtile_2__pin_inpad_0_
+ top_width_0_height_0_subtile_3__pin_inpad_0_
XFILLER_27_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_top_track_6.mux_l2_in_1_ net190 net25 sb_8__0_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__0_.mux_top_track_0.mux_l2_in_1__A1 net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout149 net68 VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_4
Xsb_8__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_46.out sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold181 sb_8__0_.mem_left_track_5.mem_out\[0\] VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold192 net240 VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold170 net229 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_37_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk net390
+ net148 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_22.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__124__A sb_8__0_.mux_left_track_3.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_top_track_22.mux_l2_in_0__174 VGND VGND VPWR VPWR net174 sb_8__0_.mux_top_track_22.mux_l2_in_0__174/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_20_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk net358
+ net147 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_15.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_23_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_131_ sb_8__0_.mux_top_track_48.out VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input55_A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__119__A sb_8__0_.mux_left_track_13.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk net301
+ net144 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_4.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_114_ net34 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk net402
+ net143 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_28.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold74 net453 VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold41 net407 VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold30 net393 VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold63 net435 VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold52 net401 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold85 net483 VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input18_A chanx_left_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold96 net495 VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_31_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_left_track_11.mux_l1_in_0__S sb_8__0_.mem_left_track_11.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_5 net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__132__A sb_8__0_.mux_top_track_46.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output86_A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_49.mux_l2_in_0_ net161 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_49.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output124_A net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput86 net86 VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_12
Xoutput97 net97 VGND VGND VPWR VPWR chanx_left_out[26] sky130_fd_sc_hd__buf_12
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__S cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__127__A net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk net408
+ net149 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_9.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_51.mux_l2_in_0_ net163 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X
+ cbx_8__0_.cbx_8__0_.ccff_head VGND VGND VPWR VPWR sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__0_.mux_top_track_6.mux_l2_in_0_ sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_22_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net151 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_left_track_35.mux_l1_in_0__A0 top_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold182 net234 VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_1__A0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
Xhold193 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
+ VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold160 net220 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold171 sb_8__0_.mem_top_track_28.ccff_tail VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_37_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_left_track_5.mux_l2_in_0__A0 net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_0__A0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_6_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_6_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_top_track_6.mux_l1_in_1_ top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ net73 sb_8__0_.mem_top_track_6.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_130_ sb_8__0_.mux_top_track_50.out VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_2
Xsb_8__0_.mux_left_track_49.mux_l2_in_0__161 VGND VGND VPWR VPWR net161 sb_8__0_.mux_left_track_49.mux_l2_in_0__161/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_2_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input48_A chany_top_in[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_ net195 net51 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk net294
+ net144 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_4.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_113_ net35 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A0 net43 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__S cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk net398
+ net143 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_28.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xhold31 net375 VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold86 net486 VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold53 net467 VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold64 net437 VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold20 net359 VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold42 net421 VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold75 net463 VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold97 net500 VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_31_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_6 net168 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_ net45 net31 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output79_A net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net149 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold312_A cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xoutput87 net87 VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_12
Xoutput98 net98 VGND VGND VPWR VPWR chanx_left_out[27] sky130_fd_sc_hd__buf_12
XFILLER_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input30_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output117_A net117 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk net460
+ net146 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_40.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X net78 VGND VGND VPWR
+ VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X sky130_fd_sc_hd__mux2_1
XFILLER_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout148_A net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold320 net322 VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk net448
+ net150 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_33.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mux_top_track_18.mux_l2_in_0_ sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_18.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xsb_8__0_.mux_top_track_34.mux_l2_in_0__180 VGND VGND VPWR VPWR net180 sb_8__0_.mux_top_track_34.mux_l2_in_0__180/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_20.mux_l2_in_0_ net173 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_20.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_left_track_49.mux_l1_in_0_ top_width_0_height_0_subtile_2__pin_inpad_0_
+ net48 sb_8__0_.mem_left_track_49.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
Xhold161 sb_8__0_.mem_top_track_46.ccff_tail VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_1__A1 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_16.mux_l1_in_1__170 VGND VGND VPWR VPWR net170 sb_8__0_.mux_top_track_16.mux_l1_in_1__170/LO
+ sky130_fd_sc_hd__conb_1
Xhold194 net230 VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold172 net226 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold183 sb_8__0_.mem_top_track_34.mem_out\[0\] VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold150 net219 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_0__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_51.mux_l1_in_0_ top_width_0_height_0_subtile_3__pin_inpad_0_
+ net49 sb_8__0_.mem_left_track_51.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_6.mux_l1_in_0_ net70 net75 sb_8__0_.mem_top_track_6.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net152 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_left_track_9.mux_l1_in_0__S sb_8__0_.mem_left_track_9.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_18.mux_l1_in_1_ net171 net31 sb_8__0_.mem_top_track_18.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__151__A sb_8__0_.mux_top_track_8.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_ net25 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_hold175_A sb_8__0_.mem_left_track_15.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk net336
+ net152 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_4.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_34_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_112_ net36 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input60_A chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A1 net32 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__D net340 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__146__A sb_8__0_.mux_top_track_18.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_left_track_5.mux_l2_in_0_ net162 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_5.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold65 net455 VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold21 net357 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold76 net473 VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold43 net387 VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold54 net389 VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold87 net487 VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_16_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold32 net377 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_2
Xhold10 net335 VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold98 net496 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_31_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net151 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_7 net173 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_ sb_8__0_.mux_left_track_31.out net8
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_left_track_51.mux_l1_in_0__A0 top_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__0_.mux_top_track_34.mux_l1_in_0__A0 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out[1] sky130_fd_sc_hd__ebufn_8
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__A1 net50 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold305_A sb_8__0_.mem_top_track_46.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput88 net88 VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_12
Xoutput77 net77 VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_12
Xsb_8__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_7.out sky130_fd_sc_hd__clkbuf_2
Xoutput99 net99 VGND VGND VPWR VPWR chanx_left_out[28] sky130_fd_sc_hd__buf_12
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A0 sb_8__0_.mux_left_track_3.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input23_A chanx_left_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_4_0_prog_clk net366
+ net146 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_40.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output91_A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold310 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR net510
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold321 net1 VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk net462
+ net150 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_33.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__0_.mux_top_track_26.mux_l1_in_0__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_left_track_15.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_15.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold31_A net375 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold140 net209 VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold162 net218 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 sb_8__0_.mem_top_track_40.ccff_tail VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_12_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xhold184 net237 VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold173 sb_8__0_.mem_top_track_18.ccff_tail VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold195 sb_8__0_.mem_top_track_32.ccff_tail VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__149__A sb_8__0_.mux_top_track_12.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__CLK clknet_4_15_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk net305
+ net147 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_46.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_4_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_18.mux_l1_in_0_ top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ net70 sb_8__0_.mem_top_track_18.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__0_.mux_left_track_9.mux_l1_in_0__A0 top_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_20.mux_l1_in_0_ net32 net71 sb_8__0_.mem_top_track_20.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_32.mux_l2_in_0_ net179 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_32.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_111_ sb_8__0_.mux_left_track_29.out VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input53_A chany_top_in[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_top_track_42.mux_l1_in_0__A0 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_0__A0 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold285_A cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xhold22 net355 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold11 net333 VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold55 net441 VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold66 net447 VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold77 net457 VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold44 net411 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold88 net489 VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold33 net379 VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold99 net499 VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_8 net173 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_ sb_8__0_.mux_left_track_19.out net15
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_34.mux_l1_in_0__A1 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput89 net89 VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_12
Xoutput78 net78 VGND VGND VPWR VPWR ccff_tail_0 sky130_fd_sc_hd__buf_12
Xsb_8__0_.mux_left_track_5.mux_l1_in_0_ top_width_0_height_0_subtile_2__pin_inpad_0_
+ net44 sb_8__0_.mem_left_track_5.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A1 net23 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_16_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input16_A chanx_left_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1__S cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_9_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold322 ccff_head_1 VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold300 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR net500
+ sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold311 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR VPWR net511
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input8_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output122_A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_32_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net63 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR top_width_0_height_0_subtile_3__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
Xsb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk net308
+ net144 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_14.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_35_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold130 net207 VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold152 net217 VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold141 sb_8__0_.mem_top_track_12.ccff_tail VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold163 sb_8__0_.mem_top_track_16.ccff_tail VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold185 sb_8__0_.mem_top_track_20.mem_out\[0\] VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_12_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold174 net227 VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__D net418 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold196 net246 VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_26_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_8.out sky130_fd_sc_hd__clkbuf_1
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk net418
+ net147 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_46.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold113_A net516 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__CLK clknet_4_15_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_left_track_9.mux_l1_in_0__A1 net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_0__A0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_5_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_5_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_28_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_left_track_5.mux_l1_in_0__S sb_8__0_.mem_left_track_5.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_110_ sb_8__0_.mux_left_track_31.out VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input46_A chany_top_in[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__0_.mux_top_track_42.mux_l1_in_0__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_0__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold34 net381 VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold12 net347 VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold56 net451 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold23 net353 VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold45 net413 VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold78 net471 VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold89 net488 VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold67 net439 VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk net478
+ net151 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_16_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_top_track_32.mux_l1_in_0_ net9 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ sb_8__0_.mem_top_track_32.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_ sb_8__0_.mux_left_track_7.out net21
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_19.mux_l2_in_0_ net153 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_19.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__0_.mux_top_track_44.mux_l2_in_0_ sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_44.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_38_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput79 net79 VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_12
XFILLER_0_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output77_A net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold323 net317 VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_1_0_prog_clk
+ net296 net143 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xhold301 sb_8__0_.mem_top_track_12.mem_out\[0\] VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold312 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR net512
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_26_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output115_A net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_44.mux_l1_in_1_ net186 net16 sb_8__0_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_40_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk net342
+ net144 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_14.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__0_.mux_top_track_6.mux_l2_in_1__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__0_.mux_top_track_22.mux_l1_in_0__S sb_8__0_.mem_top_track_22.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout146_A net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold175 sb_8__0_.mem_left_track_15.mem_out\[0\] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkbuf_2
Xhold120 net202 VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold131 sb_8__0_.mem_left_track_29.mem_out\[0\] VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold153 sb_8__0_.mem_top_track_6.ccff_tail VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold186 net248 VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold164 net225 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold142 net213 VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold197 sb_8__0_.mem_top_track_26.ccff_tail VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_37_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input76_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_0__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_20.out sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net66 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR top_width_0_height_0_subtile_0__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_9_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1__A0 sb_8__0_.mux_left_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input39_A chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold79 net481 VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold35 net403 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 net395 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold57 net425 VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold24 net365 VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold13 net341 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold68 net431 VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk net452
+ net151 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_51.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_14.out sky130_fd_sc_hd__clkbuf_1
XFILLER_12_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_ sb_8__0_.mux_left_track_1.out net24
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__0_.mux_top_track_36.mux_l2_in_0__A0 net181 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A0 net36 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1__S cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold290_A sb_8__0_.mem_top_track_6.mem_out\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_1_0_prog_clk
+ net299 net143 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold324 net201 VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold313 sb_8__0_.mem_top_track_0.mem_out\[0\] VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold302 sb_8__0_.mem_top_track_8.mem_out\[1\] VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_left_track_11.mux_l2_in_0__A0 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_19.mux_l1_in_0_ top_width_0_height_0_subtile_3__pin_inpad_0_
+ net61 sb_8__0_.mem_left_track_19.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input21_A chanx_left_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_44.mux_l1_in_0_ top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ net71 sb_8__0_.mem_top_track_44.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_4.mux_l2_in_1__183 VGND VGND VPWR VPWR net183 sb_8__0_.mux_top_track_4.mux_l2_in_1__183/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_35_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold110 net509 VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold176 net231 VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold132 net208 VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold154 net223 VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold121 net517 VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold143 sb_8__0_.mem_top_track_26.mem_out\[0\] VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold165 sb_8__0_.mem_top_track_38.ccff_tail VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold187 sb_8__0_.mem_top_track_48.ccff_tail VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold198 net247 VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold253_A sb_8__0_.mem_left_track_13.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0__CLK clknet_4_15_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_left_track_33.mux_l2_in_0_ net157 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_33.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__0_.mux_left_track_17.mux_l2_in_0__S sb_8__0_.mem_left_track_17.ccff_tail
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input69_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_1__A0 net186 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_20.mux_l2_in_0__173 VGND VGND VPWR VPWR net173 sb_8__0_.mux_top_track_20.mux_l2_in_0__173/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_2.mux_l3_in_0_ sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X sb_8__0_.mem_top_track_2.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_6_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__S cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net152 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_099_ net50 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_2
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_42.out sky130_fd_sc_hd__clkbuf_1
Xsb_8__0_.mux_top_track_2.mux_l2_in_1_ net172 net3 sb_8__0_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
Xhold58 net423 VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold14 net337 VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold69 net443 VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold25 net363 VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold47 net397 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold36 net399 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__097__A net52 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input51_A chany_top_in[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output138_A net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A1 net10 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_30_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk net370
+ net145 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_32.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_38_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_36.out sky130_fd_sc_hd__clkbuf_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk
+ net314 net145 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold325 net318 VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold303 sb_8__0_.mem_top_track_18.mem_out\[0\] VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold314 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR VPWR net514
+ sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_26_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input14_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_left_track_49.mux_l1_in_0__A0 top_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold122 net519 VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold144 net215 VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold133 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
+ VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold111 net510 VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold100 net502 VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold188 net243 VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold177 sb_8__0_.mem_top_track_42.ccff_tail VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input6_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold166 net224 VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold155 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold199 sb_8__0_.mem_top_track_24.mem_out\[0\] VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_37_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__195 VGND VGND VPWR VPWR net195 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__195/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_1__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output120_A net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout151_A net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_1__A0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_left_track_47.mux_l2_in_0__160 VGND VGND VPWR VPWR net160 sb_8__0_.mux_left_track_47.mux_l2_in_0__160/LO
+ sky130_fd_sc_hd__conb_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_top_track_48.mux_l1_in_1__188 VGND VGND VPWR VPWR net188 sb_8__0_.mux_top_track_48.mux_l1_in_1__188/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_14_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_top_track_46.mux_l2_in_0__S sb_8__0_.mem_top_track_46.ccff_tail
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_left_track_33.mux_l1_in_0_ top_width_0_height_0_subtile_2__pin_inpad_0_
+ net39 sb_8__0_.mem_left_track_33.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_45.mux_l2_in_0_ net159 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_45.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_2
XFILLER_19_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_098_ net51 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__D net472 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_2.mux_l2_in_0_ sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_2.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_0_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold26 net371 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold15 net343 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold59 net405 VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold48 net385 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold37 net383 VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_12_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input44_A chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_4_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_4_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk net406
+ net145 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_32.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_2.mux_l1_in_1_ top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ net74 sb_8__0_.mem_top_track_2.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold326 net2 VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold304 sb_8__0_.mem_top_track_0.mem_out\[1\] VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__clkdlybuf4s25_1
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_1_0_prog_clk
+ net414 net143 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold315 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR net515
+ sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_10_0_prog_clk net334 net152 VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold167 sb_8__0_.mem_left_track_1.ccff_head VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold156 net222 VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold123 net521 VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold134 net211 VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold101 net498 VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold112 net511 VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold145 sb_8__0_.mem_top_track_22.ccff_tail VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold178 net232 VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold189 sb_8__0_.mem_top_track_20.ccff_tail VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_sb_8__0_.mux_left_track_15.mux_l1_in_0__A0 top_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk net450
+ net146 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_38.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_26_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output113_A net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout144_A net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_1__A1 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input74_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A0 net45 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_22_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__0_.mux_left_track_13.mux_l2_in_0__S sb_8__0_.mem_left_track_13.ccff_tail
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__S cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_097_ net52 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold82_A net465 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold38 net409 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold27 net373 VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold16 net345 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold49 net415 VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__A0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold221_A sb_8__0_.mem_top_track_22.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_top_track_14.mux_l2_in_0_ sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_14.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_3_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input37_A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_149_ sb_8__0_.mux_top_track_12.out VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_0__S sb_8__0_.mem_top_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_left_track_45.mux_l1_in_0_ top_width_0_height_0_subtile_0__pin_inpad_0_
+ net46 sb_8__0_.mem_left_track_45.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__0_.mux_top_track_6.mux_l2_in_0__S sb_8__0_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_2.mux_l1_in_0_ net71 net76 sb_8__0_.mem_top_track_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold305 sb_8__0_.mem_top_track_46.mem_out\[0\] VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold316 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR net516
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_7_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_14.mux_l1_in_1_ net169 net29 sb_8__0_.mem_top_track_14.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_1_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_left_track_51.mux_l2_in_0__163 VGND VGND VPWR VPWR net163 sb_8__0_.mux_left_track_51.mux_l2_in_0__163/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_23_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold157 sb_8__0_.mem_left_track_13.ccff_tail VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold168 net228 VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold179 sb_8__0_.mem_top_track_0.ccff_tail VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold146 net216 VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold124 net204 VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold102 net501 VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold113 net516 VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold135 sb_8__0_.mem_top_track_2.ccff_tail VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk net420
+ net145 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_38.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_32_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__0_.mux_left_track_9.mux_l2_in_0__165 VGND VGND VPWR VPWR net165 sb_8__0_.mux_left_track_9.mux_l2_in_0__165/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_40_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_1.mux_l2_in_0_ sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_left_track_1.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net152 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_3.out sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A1 net31 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_input67_A isol_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk net295
+ net148 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_1.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_11.out sky130_fd_sc_hd__dlymetal6s2s_1
Xsb_8__0_.mux_left_track_1.mux_l1_in_1_ net196 top_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_8__0_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_096_ net53 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_35.mux_l2_in_0__158 VGND VGND VPWR VPWR net158 sb_8__0_.mux_left_track_35.mux_l2_in_0__158/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_37_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_top_track_42.mux_l2_in_0__S sb_8__0_.mem_top_track_42.ccff_tail
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold39 net417 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold28 net367 VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold17 net351 VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__A1 net51 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_1__S sb_8__0_.mem_top_track_48.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__A0 sb_8__0_.mux_left_track_5.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_left_track_31.mux_l1_in_0__A0 top_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_1__A0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_148_ sb_8__0_.mux_top_track_14.out VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_14.mux_l1_in_0__A0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output136_A net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A0 sb_8__0_.mux_left_track_13.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net152 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold317 ccff_head VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold306 sb_8__0_.mem_top_track_16.mem_out\[0\] VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_7_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_14.mux_l1_in_0_ top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ net76 sb_8__0_.mem_top_track_14.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_0_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_26.mux_l2_in_0_ net176 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_26.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__103__A sb_8__0_.mux_left_track_45.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold158 net221 VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__clkbuf_1
Xhold125 sb_8__0_.mem_left_track_17.mem_out\[0\] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold147 sb_8__0_.mem_left_track_9.mem_out\[0\] VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold169 sb_8__0_.mem_top_track_32.mem_out\[0\] VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_7_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold103 net503 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold114 net512 VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold136 net210 VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input12_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk net289
+ net147 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_11.ccff_tail sky130_fd_sc_hd__dfrtp_2
XFILLER_1_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__S cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk net388
+ net148 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_50.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_left_track_1.mux_l1_in_1__A1 top_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1__D net376 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_left_track_1.mux_l1_in_0_ top_width_0_height_0_subtile_0__pin_inpad_0_
+ net54 sb_8__0_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_top_track_22.mux_l1_in_0__A0 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_5_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold18 net361 VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold29 net369 VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_24_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__A1 net22 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_4.out sky130_fd_sc_hd__clkbuf_1
XFILLER_30_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__0_.mux_left_track_31.mux_l1_in_0__A1 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_33.out sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_1__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_147_ sb_8__0_.mux_top_track_16.out VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_2
XANTENNA__106__A net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_14.mux_l1_in_0__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold157_A sb_8__0_.mem_left_track_13.ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input42_A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A1 net18 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold318 net321 VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold307 sb_8__0_.mem_top_track_2.mem_out\[1\] VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_38_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk net382
+ net147 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_5.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk net434
+ net151 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_49.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_3_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_3_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_17_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__S cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold126 net205 VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_31_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold104 net504 VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold115 net514 VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold148 net212 VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold137 sb_8__0_.mem_left_track_5.ccff_tail VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold159 sb_8__0_.mem_top_track_30.mem_out\[0\] VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__114__A net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_26.mux_l1_in_0_ net6 net74 sb_8__0_.mem_top_track_26.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__0_.mux_top_track_30.mux_l1_in_0__A0 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk net412
+ net147 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_11.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mux_top_track_38.mux_l2_in_0_ net182 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_38.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output111_A net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__109__A sb_8__0_.mux_left_track_33.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_left_track_15.mux_l2_in_0_ net199 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_15.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_top_track_40.mux_l2_in_0_ net184 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_40.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1__CLK clknet_4_15_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_14_0_prog_clk net304
+ net151 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input72_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_top_track_22.mux_l1_in_0__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold19 net349 VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk net400
+ net148 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_24.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_3_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_146_ sb_8__0_.mux_top_track_18.out VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
XANTENNA__122__A sb_8__0_.mux_left_track_7.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk net326
+ net150 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_17.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_33_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_37_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold317_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input35_A chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__117__A sb_8__0_.mux_left_track_17.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold308 sb_8__0_.mem_top_track_14.mem_out\[0\] VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__0_.mux_left_track_5.mux_l1_in_0__A0 top_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk net340
+ net147 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_5.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk net438
+ net151 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_49.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_129_ net20 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_2
Xhold319 net203 VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_1__S sb_8__0_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold267_A sb_8__0_.mem_top_track_48.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold127 sb_8__0_.mem_left_track_31.mem_out\[0\] VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold138 net214 VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold43_A net387 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold105 net505 VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold116 net515 VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold149 sb_8__0_.mem_top_track_10.ccff_head VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_10.out sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_0__A0 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__193 VGND VGND VPWR VPWR net193 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__193/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_49.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_49.out sky130_fd_sc_hd__clkbuf_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__130__A sb_8__0_.mux_top_track_50.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__0_.mux_top_track_30.mux_l1_in_0__A1 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk net309
+ net151 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_0.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_input65_A gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk net346
+ net148 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_24.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xinput1 net520 VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_38.mux_l1_in_0_ net12 net76 sb_8__0_.mem_top_track_38.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_24_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0_prog_clk prog_clk VGND VGND VPWR VPWR clknet_0_prog_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_3_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_left_track_15.mux_l1_in_0_ top_width_0_height_0_subtile_1__pin_inpad_0_
+ net59 sb_8__0_.mem_left_track_15.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_145_ sb_8__0_.mux_top_track_20.out VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_2
Xsb_8__0_.mux_top_track_40.mux_l1_in_0_ net13 net69 sb_8__0_.mem_top_track_40.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
Xsb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk net466
+ net150 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_17.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_33_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2__A0 net26 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_21_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_7.mux_l1_in_1__164 VGND VGND VPWR VPWR net164 sb_8__0_.mux_left_track_7.mux_l1_in_1__164/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input28_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold309 sb_8__0_.mem_top_track_44.mem_out\[0\] VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_128_ net21 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_9_0_prog_clk net290
+ net148 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_6.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput70 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ VGND VGND VPWR
+ VPWR net70 sky130_fd_sc_hd__buf_2
XANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net152 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1__S cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output134_A net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_2.mux_l2_in_1__172 VGND VGND VPWR VPWR net172 sb_8__0_.mux_top_track_2.mux_l2_in_1__172/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA__128__A net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold117 net522 VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold128 net206 VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold139 sb_8__0_.mem_left_track_3.ccff_tail VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold106 net507 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkdlybuf4s50_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_0__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_32.out sky130_fd_sc_hd__clkbuf_1
Xsb_8__0_.mux_top_track_46.mux_l1_in_1__187 VGND VGND VPWR VPWR net187 sb_8__0_.mux_top_track_46.mux_l1_in_1__187/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_10_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_4_14_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input10_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__141__A sb_8__0_.mux_top_track_28.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net151 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__D net378 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk net320
+ net152 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_0.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input58_A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__A1 net9 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput2 net525 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_24_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_26.out sky130_fd_sc_hd__clkbuf_2
XFILLER_24_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_144_ sb_8__0_.mux_top_track_22.out VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__S cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_left_track_29.mux_l2_in_0__154 VGND VGND VPWR VPWR net154 sb_8__0_.mux_left_track_29.mux_l2_in_0__154/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_37_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk net287
+ net148 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_6.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_output89_A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_127_ net22 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput60 chany_top_in[7] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
Xinput71 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ VGND VGND VPWR
+ VPWR net71 sky130_fd_sc_hd__buf_2
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold322_A ccff_head_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_left_track_29.mux_l1_in_0__A0 top_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input40_A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__144__A sb_8__0_.mux_top_track_22.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_10.mux_l3_in_0_ sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sb_8__0_.mem_top_track_10.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
Xhold118 net524 VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold107 net506 VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkdlybuf4s50_1
Xsb_8__0_.mux_top_track_50.mux_l1_in_1__189 VGND VGND VPWR VPWR net189 sb_8__0_.mux_top_track_50.mux_l1_in_1__189/LO
+ sky130_fd_sc_hd__conb_1
Xhold129 sb_8__0_.mem_top_track_34.ccff_tail VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_39_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk net293
+ net144 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_10.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_22_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_2_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_2_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_8__0_.mux_top_track_8.mux_l3_in_0_ sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X sb_8__0_.mem_top_track_10.ccff_head
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk net436
+ net146 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_42.ccff_tail sky130_fd_sc_hd__dfrtp_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__CLK clknet_4_15_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net151 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__0_.mux_left_track_3.mux_l2_in_0__S sb_8__0_.mem_left_track_3.ccff_tail
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_10.mux_l2_in_1_ net167 net27 sb_8__0_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
+ net152 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk net456
+ net150 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_35.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold235_A sb_8__0_.mem_top_track_42.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold290 sb_8__0_.mem_top_track_6.mem_out\[1\] VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_8.mux_l2_in_1_ net191 net26 sb_8__0_.mem_top_track_8.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XANTENNA__152__A sb_8__0_.mux_top_track_6.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 chanx_left_in[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input70_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_143_ sb_8__0_.mux_top_track_24.out VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_48.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_1__A0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_30 net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_15_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_15_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XFILLER_11_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk net432
+ net148 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_6.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
X_126_ net23 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput72 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_ VGND VGND VPWR
+ VPWR net72 sky130_fd_sc_hd__buf_2
Xinput50 chany_top_in[25] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
Xinput61 chany_top_in[8] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
XFILLER_21_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold315_A cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input33_A chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_40.mux_l2_in_0__A0 net184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_15.mux_l2_in_0__199 VGND VGND VPWR VPWR net199 sb_8__0_.mux_left_track_15.mux_l2_in_0__199/LO
+ sky130_fd_sc_hd__conb_1
Xhold108 net508 VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold119 net526 VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_109_ sb_8__0_.mux_left_track_33.out VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk net298
+ net144 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_10.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hold265_A sb_8__0_.mem_left_track_15.ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_A
+ net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk net352
+ net146 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_42.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ net77 net67 VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XFILLER_38_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_top_track_10.mux_l2_in_0_ sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_10.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk net484
+ net150 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_35.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_ net192 sb_8__0_.mux_left_track_49.out
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold280 net284 VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold291 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\] VGND VGND VPWR VPWR net491
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_left_track_33.mux_l2_in_0__157 VGND VGND VPWR VPWR net157 sb_8__0_.mux_left_track_33.mux_l2_in_0__157/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_1__A1 top_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_8.mux_l2_in_0_ sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_8.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput4 chanx_left_in[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_sb_8__0_.mux_left_track_45.mux_l1_in_0__A0 top_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_top_track_10.mux_l1_in_1_ top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_ sb_8__0_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_10_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hold178_A net232 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_142_ sb_8__0_.mux_top_track_26.out VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk net468
+ net147 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_48.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_ net41 net5 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input63_A gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_20 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_31 net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_1__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_8.mux_l1_in_1_ top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ net74 sb_8__0_.mem_top_track_8.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X cbx_8__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
X_125_ sb_8__0_.mux_left_track_1.out VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_2
XFILLER_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput62 chany_top_in[9] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput73 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ VGND VGND VPWR
+ VPWR net73 sky130_fd_sc_hd__clkbuf_2
Xinput40 chany_top_in[16] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
Xinput51 chany_top_in[26] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
XFILLER_29_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2__S cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input26_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold109 net513 VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_7_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_108_ sb_8__0_.mux_left_track_35.out VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_10_0_prog_clk net350
+ net152 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_10.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__D net305 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__0_.mux_top_track_36.mux_l1_in_0__A0 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_ net28 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net64 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR top_width_0_height_0_subtile_2__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk net307
+ net144 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_16.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold281 sb_8__0_.mem_left_track_1.mem_out\[0\] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold270 net270 VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_clkbuf_0_prog_clk_A prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold292 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\] VGND VGND VPWR VPWR net492
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_33_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_0__S sb_8__0_.mem_top_track_46.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail net67
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
Xinput5 chanx_left_in[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_10.mux_l1_in_0_ net72 net69 sb_8__0_.mem_top_track_10.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_20_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__0_.mux_top_track_28.mux_l1_in_0__A1 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_1_0_prog_clk
+ net291 net143 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk net362
+ net147 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_48.mem_out\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_141_ sb_8__0_.mux_top_track_28.out VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_2
Xsb_8__0_.mux_top_track_22.mux_l2_in_0_ net174 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_22.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input56_A chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_ net35 net11 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_left_track_11.mux_l1_in_0__A0 top_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_21 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_10 net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 net178 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold288_A sb_8__0_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold190_A net254 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_8.mux_l1_in_0_ net71 net76 sb_8__0_.mem_top_track_8.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_124_ sb_8__0_.mux_left_track_3.out VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__D net412 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput74 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_ VGND VGND VPWR
+ VPWR net74 sky130_fd_sc_hd__buf_2
Xinput52 chany_top_in[27] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput41 chany_top_in[17] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
Xinput30 chanx_left_in[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
Xinput63 gfpga_pad_io_soc_in[0] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_40_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input19_A chanx_left_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_107_ net41 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_2
XANTENNA_output87_A net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_0.out sky130_fd_sc_hd__clkbuf_1
Xsb_8__0_.mux_left_track_7.mux_l2_in_0_ sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_left_track_7.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_4_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output125_A net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_0__A0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_1_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0__A cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_36.mux_l1_in_0__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_left_track_7.mux_l1_in_1_ net164 top_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_8__0_.mem_left_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold271 sb_8__0_.mem_left_track_11.ccff_tail VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold260 net272 VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__clkdlybuf4s50_1
Xsb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_2_0_prog_clk net428
+ net144 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_16.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xhold282 net279 VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold293 sb_8__0_.mem_top_track_50.mem_out\[0\] VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__clkbuf_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_1_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_1_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_8__0_.mux_left_track_9.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_9.out sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_8__0_.mux_left_track_13.mux_l1_in_0__S sb_8__0_.mem_left_track_13.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput6 chanx_left_in[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_20_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_1_0_prog_clk
+ net311 net143 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_140_ sb_8__0_.mux_top_track_30.out VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_2
XFILLER_23_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input49_A chany_top_in[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_ sb_8__0_.mux_left_track_13.out net18
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_2_0_prog_clk net394 net144 VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A1 net17 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_17.out sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_22 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_11 net179 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 net389 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput140 net140 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[1] sky130_fd_sc_hd__buf_12
XFILLER_28_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1__CLK clknet_4_15_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_123_ sb_8__0_.mux_left_track_5.out VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_4_6_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__S cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput20 chanx_left_in[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_2
Xinput31 chanx_left_in[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput42 chany_top_in[18] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
Xinput75 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ VGND VGND VPWR VPWR
+ net75 sky130_fd_sc_hd__buf_2
Xinput53 chany_top_in[28] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
Xinput64 gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
Xsb_8__0_.mux_top_track_22.mux_l1_in_0_ net4 net72 sb_8__0_.mem_top_track_22.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_40_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_top_track_34.mux_l2_in_0_ net180 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_34.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_106_ net42 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_left_track_11.mux_l2_in_0_ net197 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_11.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_14_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_14_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_28.mux_l2_in_0__177 VGND VGND VPWR VPWR net177 sb_8__0_.mux_top_track_28.mux_l2_in_0__177/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_0__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input31_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output118_A net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout149_A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_0__A0 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0__S cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_51.out sky130_fd_sc_hd__clkbuf_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_7.mux_l1_in_0_ top_width_0_height_0_subtile_0__pin_inpad_0_
+ net55 sb_8__0_.mem_left_track_7.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold272 net278 VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold283 sb_8__0_.mem_left_track_33.ccff_tail VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold261 sb_8__0_.mem_left_track_31.ccff_tail VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold250 net271 VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold294 sb_8__0_.mem_top_track_4.mem_out\[0\] VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_26_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 chanx_left_in[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net152 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ net316 net145 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_ sb_8__0_.mux_left_track_7.out net21
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_45.out sky130_fd_sc_hd__clkbuf_1
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_8.mux_l2_in_1__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_42.mux_l1_in_0__S sb_8__0_.mem_top_track_42.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 net464 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput130 net130 VGND VGND VPWR VPWR chany_top_out[29] sky130_fd_sc_hd__buf_12
Xoutput141 net141 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[2] sky130_fd_sc_hd__buf_12
XFILLER_28_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__098__A net51 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input61_A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_122_ sb_8__0_.mux_left_track_7.out VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput54 chany_top_in[29] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_1
Xinput43 chany_top_in[19] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
Xinput10 chanx_left_in[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput32 chanx_left_in[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput21 chanx_left_in[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput76 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_ VGND VGND VPWR VPWR
+ net76 sky130_fd_sc_hd__buf_2
Xinput65 gfpga_pad_io_soc_in[2] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
Xsb_8__0_.mux_top_track_32.mux_l2_in_0__179 VGND VGND VPWR VPWR net179 sb_8__0_.mux_top_track_32.mux_l2_in_0__179/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold293_A sb_8__0_.mem_top_track_50.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_105_ net43 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_14.mux_l1_in_1__169 VGND VGND VPWR VPWR net169 sb_8__0_.mux_top_track_14.mux_l1_in_1__169/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_25_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold139_A sb_8__0_.mem_left_track_3.ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_6_0_prog_clk net384
+ net145 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_34.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_21_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input24_A chanx_left_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_top_track_34.mux_l1_in_0_ net10 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ sb_8__0_.mem_top_track_34.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_0__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_44.mux_l1_in_1__186 VGND VGND VPWR VPWR net186 sb_8__0_.mux_top_track_44.mux_l1_in_1__186/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_9_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_top_track_38.mux_l2_in_0__A0 net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_11.mux_l1_in_0_ top_width_0_height_0_subtile_2__pin_inpad_0_
+ net57 sb_8__0_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_46.mux_l2_in_0_ sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_46.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A0 sb_8__0_.mux_left_track_31.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold284 net285 VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold273 sb_8__0_.mem_left_track_45.ccff_tail VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold262 net273 VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold240 net267 VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold251 sb_8__0_.mem_left_track_49.ccff_tail VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold295 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\] VGND VGND VPWR VPWR net495
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_14_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 chanx_left_in[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_left_track_13.mux_l2_in_0__A0 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2__A0 net25 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk
+ net426 net143 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xsb_8__0_.mux_top_track_46.mux_l1_in_1_ net187 net17 sb_8__0_.mem_top_track_46.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ sb_8__0_.mux_left_track_1.out net24
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_13 net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net152 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_35 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_24 net493 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput120 net120 VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_12
Xoutput131 net131 VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_12
XANTENNA_sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__D net454 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput142 net142 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[3] sky130_fd_sc_hd__buf_12
XFILLER_28_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_121_ sb_8__0_.mux_left_track_9.out VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input54_A chany_top_in[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_1__A0 net187 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__S cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput44 chany_top_in[1] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
Xinput55 chany_top_in[2] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
Xinput66 gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
Xinput22 chanx_left_in[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput33 chany_top_in[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput11 chanx_left_in[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_29_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net151 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold286_A sb_8__0_.mem_left_track_17.ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_10_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_104_ net45 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_22.out sky130_fd_sc_hd__clkbuf_1
XFILLER_19_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out[0] sky130_fd_sc_hd__ebufn_8
XANTENNA_sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_6_0_prog_clk net396
+ net145 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_34.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_21_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_5.mux_l2_in_0__162 VGND VGND VPWR VPWR net162 sb_8__0_.mux_left_track_5.mux_l2_in_0__162/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input17_A chanx_left_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input9_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold151_A sb_8__0_.mem_top_track_40.ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A1 net8 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_16.out sky130_fd_sc_hd__clkbuf_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_left_track_1.mux_l1_in_0__A0 top_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold241 sb_8__0_.mem_left_track_45.mem_out\[0\] VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold274 net276 VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold230 net261 VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold252 net256 VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold263 sb_8__0_.mem_top_track_36.mem_out\[0\] VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold285 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\] VGND VGND VPWR VPWR net485
+ sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold296 sb_8__0_.mem_top_track_10.mem_out\[0\] VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__S cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput9 chanx_left_in[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_top_track_46.mux_l1_in_0_ top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ net72 sb_8__0_.mem_top_track_46.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_4_15_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_0__A0 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
Xsb_8__0_.mux_left_track_35.mux_l2_in_0_ net158 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_35.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_14 net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 sb_8__0_.mux_top_track_14.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput121 net121 VGND VGND VPWR VPWR chany_top_out[20] sky130_fd_sc_hd__buf_12
Xoutput110 net110 VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_12
Xoutput132 net132 VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_12
XFILLER_21_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_0_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_0_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_28_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_120_ sb_8__0_.mux_left_track_11.out VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_2
XFILLER_23_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input47_A chany_top_in[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_1__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1__A0 sb_8__0_.mux_left_track_7.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput45 chany_top_in[20] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
Xinput56 chany_top_in[3] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 chany_top_in[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xinput23 chanx_left_in[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
Xinput67 isol_n VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput12 chanx_left_in[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B net151 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_1__S sb_8__0_.mem_top_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_4.mux_l3_in_0_ sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X sb_8__0_.mem_top_track_4.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold181_A sb_8__0_.mem_left_track_5.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_50.out sky130_fd_sc_hd__clkbuf_2
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_103_ sb_8__0_.mux_left_track_45.out VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__0_.mux_top_track_6.mux_l2_in_1__S sb_8__0_.mem_top_track_6.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_left_track_13.mux_l2_in_0__198 VGND VGND VPWR VPWR net198 sb_8__0_.mux_left_track_13.mux_l2_in_0__198/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_30_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_4.mux_l2_in_1_ net183 net14 sb_8__0_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 net523 VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_44.out sky130_fd_sc_hd__clkbuf_1
XFILLER_21_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
+ cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR gfpga_pad_io_soc_out[2] sky130_fd_sc_hd__ebufn_8
XANTENNA_hold311_A cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_13_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_13_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output116_A net116 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold253 sb_8__0_.mem_left_track_13.mem_out\[0\] VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold242 net255 VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold220 net251 VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold231 sb_8__0_.mem_top_track_4.ccff_tail VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold275 sb_8__0_.mem_left_track_35.ccff_tail VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold286 sb_8__0_.mem_left_track_17.ccff_tail VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold297 sb_8__0_.mem_top_track_10.mem_out\[1\] VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold264 net275 VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_31.mux_l2_in_0__156 VGND VGND VPWR VPWR net156 sb_8__0_.mux_left_track_31.mux_l2_in_0__156/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_5_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_38.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_38.out sky130_fd_sc_hd__clkbuf_1
XFILLER_32_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_0__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_15 net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 net171 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput111 net111 VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_12
Xoutput133 net133 VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_12
XANTENNA_sb_8__0_.mux_left_track_17.mux_l1_in_0__A0 top_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput122 net122 VGND VGND VPWR VPWR chany_top_out[21] sky130_fd_sc_hd__buf_12
Xoutput100 net100 VGND VGND VPWR VPWR chanx_left_out[29] sky130_fd_sc_hd__buf_12
XFILLER_36_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1__A1 net21 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xinput13 chanx_left_in[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
Xinput68 prog_reset VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput35 chany_top_in[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput46 chany_top_in[21] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
Xinput57 chany_top_in[4] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
Xinput24 chanx_left_in[29] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk net442
+ net152 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_45.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk net482
+ net151 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_1.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_25_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_1__A1 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_102_ sb_8__0_.mux_left_track_47.out VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_35.mux_l1_in_0_ top_width_0_height_0_subtile_3__pin_inpad_0_
+ net40 sb_8__0_.mem_left_track_35.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_left_track_47.mux_l2_in_0_ net160 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_47.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__104__A net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_top_track_4.mux_l2_in_0_ sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_4.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_39_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2 net319 VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_15_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold137_A sb_8__0_.mem_left_track_5.ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
Xsb_8__0_.mux_top_track_10.mux_l2_in_1__167 VGND VGND VPWR VPWR net167 sb_8__0_.mux_top_track_10.mux_l2_in_1__167/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_13_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input22_A chanx_left_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output109_A net109 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output90_A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold254 net274 VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold276 net283 VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold265 sb_8__0_.mem_left_track_15.ccff_tail VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__clkbuf_2
Xhold221 sb_8__0_.mem_top_track_22.mem_out\[0\] VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold210 net238 VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold243 sb_8__0_.mem_top_track_24.ccff_tail VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold232 net268 VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold287 sb_8__0_.mem_top_track_6.mem_out\[0\] VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold298 sb_8__0_.mem_top_track_4.mem_out\[1\] VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_26_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_top_track_4.mux_l1_in_1_ top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_ sb_8__0_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0__CLK clknet_4_15_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1__S cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk net386
+ net148 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_20.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_2_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_ net193 sb_8__0_.mux_left_track_51.out
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1__CLK clknet_4_15_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__112__A net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk net454
+ net147 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_13.ccff_tail sky130_fd_sc_hd__dfrtp_2
XANTENNA_16 net197 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_27 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput112 net112 VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_12
Xoutput134 net134 VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_12
Xoutput123 net123 VGND VGND VPWR VPWR chany_top_out[22] sky130_fd_sc_hd__buf_12
Xoutput101 net101 VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_12
XFILLER_23_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold217_A sb_8__0_.mem_top_track_44.ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput36 chany_top_in[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_2
XANTENNA__107__A net41 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput14 chanx_left_in[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xinput25 chanx_left_in[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput58 chany_top_in[5] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_1
Xinput69 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_ VGND VGND VPWR
+ VPWR net69 sky130_fd_sc_hd__buf_2
Xinput47 chany_top_in[22] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk net476
+ net152 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_45.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk net368
+ net151 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_1.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_25_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_ net42 net4 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
X_101_ sb_8__0_.mux_left_track_49.out VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input52_A chany_top_in[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X cbx_8__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__S cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__120__A sb_8__0_.mux_left_track_11.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3 net518 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_22_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_16.mux_l2_in_0_ sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_16.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk net288
+ net150 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_7.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input15_A chanx_left_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_left_track_33.mux_l1_in_0__A0 top_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_1__A0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_left_track_47.mux_l1_in_0_ top_width_0_height_0_subtile_1__pin_inpad_0_
+ net47 sb_8__0_.mem_left_track_47.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__115__A net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_16.mux_l1_in_0__A0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold266 net282 VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold255 sb_8__0_.mem_left_track_35.mem_out\[0\] VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold288 sb_8__0_.mem_left_track_11.mem_out\[0\] VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold211 sb_8__0_.mem_left_track_11.ccff_head VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold233 sb_8__0_.mem_left_track_49.mem_out\[0\] VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold277 sb_8__0_.mem_left_track_51.mem_out\[0\] VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold200 net236 VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold244 net269 VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold222 net242 VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold299 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR net499
+ sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_38_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input7_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_4.mux_l1_in_0_ net72 net69 sb_8__0_.mem_top_track_4.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_14_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A0 sb_8__0_.mux_left_track_17.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_16.mux_l1_in_1_ net170 net30 sb_8__0_.mem_top_track_16.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_36_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output121_A net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout152_A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_9_0_prog_clk net374
+ net148 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_20.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_2_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_ net27 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A0 net41 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk net472
+ net147 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_13.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_28 net174 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput124 net124 VGND VGND VPWR VPWR chany_top_out[23] sky130_fd_sc_hd__buf_12
Xoutput113 net113 VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_12
Xoutput135 net135 VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_12
Xoutput102 net102 VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_12
XFILLER_36_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_3.mux_l2_in_0_ net155 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_3.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput48 chany_top_in[23] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
Xinput37 chany_top_in[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xinput59 chany_top_in[6] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
Xinput26 chanx_left_in[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput15 chanx_left_in[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__123__A sb_8__0_.mux_left_track_5.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk net306
+ net144 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_2.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_ net36 net10 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_5.out sky130_fd_sc_hd__dlymetal6s2s_1
X_100_ sb_8__0_.mux_left_track_51.out VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_2
XANTENNA_input45_A chany_top_in[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_2_0_prog_clk net344
+ net143 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_26.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_30_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_26.mux_l2_in_0__176 VGND VGND VPWR VPWR net176 sb_8__0_.mux_top_track_26.mux_l2_in_0__176/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk net424
+ net150 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_19.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_0_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_top_track_24.mux_l1_in_0__A0 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_13.out sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold4 net323 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_left_track_45.mux_l2_in_0__159 VGND VGND VPWR VPWR net159 sb_8__0_.mux_left_track_45.mux_l2_in_0__159/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_12_0_prog_clk net338
+ net147 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_7.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_left_track_33.mux_l1_in_0__A1 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_1__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_top_track_16.mux_l1_in_0__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_17.mux_l2_in_0__200 VGND VGND VPWR VPWR net200 sb_8__0_.mux_left_track_17.mux_l2_in_0__200/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net151 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__131__A sb_8__0_.mux_top_track_48.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold201 sb_8__0_.mem_top_track_28.mem_out\[0\] VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold256 net265 VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold223 sb_8__0_.mem_left_track_19.mem_out\[0\] VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold212 net244 VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold267 sb_8__0_.mem_top_track_48.mem_out\[0\] VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold289 sb_8__0_.mem_left_track_7.mem_out\[0\] VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__clkbuf_1
Xhold234 net260 VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold278 net281 VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold245 sb_8__0_.mem_top_track_2.mem_out\[0\] VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_26_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A1 net16 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_16.mux_l1_in_0_ top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ net69 sb_8__0_.mem_top_track_16.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_output114_A net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_2_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__126__A net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_28.mux_l2_in_0_ net177 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_28.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_12_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_12_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout145_A net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_top_track_30.mux_l2_in_0_ net178 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_30.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input75_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_ VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_18 sb_8__0_.mux_left_track_3.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 net175 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A1 net5 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput125 net125 VGND VGND VPWR VPWR chany_top_out[24] sky130_fd_sc_hd__buf_12
Xoutput114 net114 VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_12
Xoutput103 net103 VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_12
XFILLER_9_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput136 net136 VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_12
XFILLER_36_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput38 chany_top_in[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
Xinput49 chany_top_in[24] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
Xinput16 chanx_left_in[21] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput27 chanx_left_in[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0__D net466 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk net446
+ net152 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_2.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mux_top_track_30.mux_l2_in_0__178 VGND VGND VPWR VPWR net178 sb_8__0_.mux_top_track_30.mux_l2_in_0__178/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_33_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_ sb_8__0_.mux_left_track_15.out net17
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__0_.mux_top_track_32.mux_l1_in_0__A0 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_top_track_0.mux_l2_in_1__166 VGND VGND VPWR VPWR net166 sb_8__0_.mux_top_track_0.mux_l2_in_1__166/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__0_.mux_top_track_8.mux_l2_in_1__191 VGND VGND VPWR VPWR net191 sb_8__0_.mux_top_track_8.mux_l2_in_1__191/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_input38_A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk net444
+ net144 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_26.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net151 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_12.mux_l1_in_1__168 VGND VGND VPWR VPWR net168 sb_8__0_.mux_top_track_12.mux_l1_in_1__168/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_8_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_159_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
XFILLER_38_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_3.mux_l1_in_0_ top_width_0_height_0_subtile_1__pin_inpad_0_
+ net33 sb_8__0_.mem_left_track_3.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk net286
+ net150 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_19.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_7_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_24.mux_l1_in_0__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_left_track_15.mux_l2_in_0__S sb_8__0_.mem_left_track_15.ccff_tail
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__S cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold5 net325 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__129__A net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_8_0_prog_clk net300
+ net152 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_10.ccff_head sky130_fd_sc_hd__dfrtp_1
XFILLER_28_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_6.out sky130_fd_sc_hd__clkbuf_1
XFILLER_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_35.out sky130_fd_sc_hd__clkbuf_1
Xhold224 net258 VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__clkdlybuf4s50_1
Xsb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk net328
+ net150 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_31.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xhold235 sb_8__0_.mem_top_track_42.mem_out\[0\] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold213 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold202 net252 VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold257 sb_8__0_.mem_left_track_19.ccff_tail VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold268 net253 VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold246 net250 VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold279 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
+ VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input20_A chanx_left_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_0__A0 top_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__142__A sb_8__0_.mux_top_track_26.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__D net310 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_29.out sky130_fd_sc_hd__clkbuf_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input68_A prog_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_19 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xoutput126 net126 VGND VGND VPWR VPWR chany_top_out[25] sky130_fd_sc_hd__buf_12
Xoutput115 net115 VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_12
Xoutput137 net137 VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_12
Xoutput104 net104 VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_12
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__0_.mux_top_track_40.mux_l1_in_0__A0 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_0__A0 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput39 chany_top_in[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
Xinput28 chanx_left_in[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_28.mux_l1_in_0_ net7 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ sb_8__0_.mem_top_track_28.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xinput17 chanx_left_in[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dlymetal6s2s_1
Xsb_8__0_.mux_top_track_38.mux_l2_in_0__182 VGND VGND VPWR VPWR net182 sb_8__0_.mux_top_track_38.mux_l2_in_0__182/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_37_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk net380
+ net151 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_2.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_33_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_32.mux_l1_in_0__A1 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_30.mux_l1_in_0_ net8 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ sb_8__0_.mem_top_track_30.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_ sb_8__0_.mux_left_track_9.out net20
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_left_track_17.mux_l2_in_0_ net200 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_17.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xfanout150 net151 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_8
Xsb_8__0_.mux_top_track_42.mux_l2_in_0_ net185 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_42.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_158_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__150__A sb_8__0_.mux_top_track_10.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input50_A chany_top_in[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold6 net327 VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net151 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output137_A net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__145__A sb_8__0_.mux_top_track_20.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_10_0_prog_clk net410
+ net151 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_8.mem_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_28_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_44.mux_l2_in_0__S sb_8__0_.mem_top_track_44.ccff_tail
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk net440
+ net150 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_31.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xhold247 sb_8__0_.mem_left_track_33.mem_out\[0\] VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold258 net277 VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold269 sb_8__0_.mem_left_track_3.mem_out\[0\] VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold203 cbx_8__0_.cbx_8__0_.ccff_head VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold236 net263 VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold225 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold214 net245 VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_26_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input13_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input5_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_7_0_prog_clk net310
+ net146 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_44.ccff_tail sky130_fd_sc_hd__dfrtp_2
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput127 net127 VGND VGND VPWR VPWR chany_top_out[26] sky130_fd_sc_hd__buf_12
Xoutput138 net138 VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_12
Xoutput116 net116 VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_12
Xoutput105 net105 VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_12
XANTENNA_sb_8__0_.mux_top_track_40.mux_l1_in_0__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout150_A net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_0__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_12.out sky130_fd_sc_hd__clkbuf_2
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput18 chanx_left_in[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net149 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput29 chanx_left_in[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_ sb_8__0_.mux_left_track_3.out net23
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout151 net152 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_8
Xsb_8__0_.mux_left_track_11.mux_l2_in_0__197 VGND VGND VPWR VPWR net197 sb_8__0_.mux_left_track_11.mux_l2_in_0__197/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_34_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_1__A1 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_157_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_2
XFILLER_8_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__0_.mux_top_track_26.mux_l2_in_0__A0 net176 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input43_A chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold7 net329 VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_15_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_left_track_17.mux_l1_in_0_ top_width_0_height_0_subtile_2__pin_inpad_0_
+ net60 sb_8__0_.mem_left_track_17.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_9_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_9_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
Xsb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk net354
+ net151 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_8.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_11_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_42.mux_l1_in_0_ net15 net70 sb_8__0_.mem_top_track_42.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_0_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__0_.mux_left_track_29.mux_l2_in_0_ net154 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_29.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_0_0_prog_clk net324 net143 VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_left_track_11.mux_l2_in_0__S sb_8__0_.mem_left_track_11.ccff_tail
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__156__A cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold248 net266 VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold237 sb_8__0_.mem_left_track_47.ccff_tail VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__clkdlybuf4s25_1
Xsb_8__0_.mux_left_track_31.mux_l2_in_0_ net156 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_31.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xhold215 sb_8__0_.mem_left_track_1.ccff_tail VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold204 net235 VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold259 sb_8__0_.mem_top_track_40.mem_out\[0\] VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold226 net257 VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_8_0_prog_clk net302
+ net144 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_12.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0__S cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__194 VGND VGND VPWR VPWR net194 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__194/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__0_.mux_top_track_0.mux_l3_in_0_ sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sb_8__0_.mem_top_track_0.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_top_track_42.mux_l2_in_0__185 VGND VGND VPWR VPWR net185 sb_8__0_.mux_top_track_42.mux_l2_in_0__185/LO
+ sky130_fd_sc_hd__conb_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_7_0_prog_clk net378
+ net146 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_44.mem_out\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output112_A net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A0 sb_8__0_.mux_left_track_9.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput117 net117 VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_12
Xoutput128 net128 VGND VGND VPWR VPWR chany_top_out[27] sky130_fd_sc_hd__buf_12
Xoutput106 net106 VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_12
Xoutput139 net139 VGND VGND VPWR VPWR gfpga_pad_io_soc_dir[0] sky130_fd_sc_hd__buf_12
Xsb_8__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_40.out sky130_fd_sc_hd__clkbuf_1
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout143_A net149 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1__CLK clknet_4_15_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput19 chanx_left_in[24] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_input73_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_11_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__0_.mux_top_track_34.mux_l2_in_0__A0 net180 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_0.mux_l2_in_1_ net166 net24 sb_8__0_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X sky130_fd_sc_hd__mux2_1
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_34.out sky130_fd_sc_hd__clkbuf_1
Xfanout152 net68 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__buf_4
X_156_ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_2
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input36_A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold8 net331 VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__S cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_139_ sb_8__0_.mux_top_track_32.out VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__buf_2
XFILLER_7_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_28.out sky130_fd_sc_hd__clkbuf_2
XFILLER_29_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_0_0_prog_clk
+ net292 net143 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_35_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold238 net264 VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold216 net249 VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold249 sb_8__0_.mem_top_track_38.mem_out\[0\] VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold227 sb_8__0_.mem_top_track_14.ccff_tail VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold205 sb_8__0_.mem_top_track_30.ccff_tail VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_1__A0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_left_track_9.mux_l2_in_0__A0 net165 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_8_0_prog_clk net392
+ net144 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_12.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_40.mux_l2_in_0__S sb_8__0_.mem_top_track_40.ccff_tail
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_left_track_29.mux_l1_in_0_ top_width_0_height_0_subtile_0__pin_inpad_0_
+ net37 sb_8__0_.mem_left_track_29.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_top_track_42.mux_l2_in_0__A0 net185 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_left_track_31.mux_l1_in_0_ top_width_0_height_0_subtile_1__pin_inpad_0_
+ net38 sb_8__0_.mem_left_track_31.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_1__S sb_8__0_.mem_top_track_46.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A1 net20 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_40_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput107 net107 VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_12
XFILLER_13_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput129 net129 VGND VGND VPWR VPWR chany_top_out[28] sky130_fd_sc_hd__buf_12
Xoutput118 net118 VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_12
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
+ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ sky130_fd_sc_hd__inv_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
+ net65 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
+ VGND VGND VPWR VPWR top_width_0_height_0_subtile_1__pin_inpad_0_ sky130_fd_sc_hd__ebufn_8
XFILLER_10_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input66_A gfpga_pad_io_soc_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_0.mux_l2_in_0_ sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_0.mem_out\[1\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0__CLK clknet_4_15_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk net303
+ net148 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_18.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_9_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_left_track_9.mux_l2_in_0__S sb_8__0_.mem_left_track_11.ccff_head
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
+ net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_155_ sb_8__0_.mux_top_track_0.out VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_ clknet_4_5_0_prog_clk
+ net280 net145 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__D net289 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_top_track_0.mux_l1_in_1_ top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ net73 sb_8__0_.mem_top_track_0.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xhold9 net339 VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input29_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_left_track_47.mux_l1_in_0__A0 top_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_138_ sb_8__0_.mux_top_track_34.out VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_0_0_prog_clk
+ net297 net143 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_output135_A net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__S cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold217 sb_8__0_.mem_top_track_44.ccff_tail VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold206 net259 VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold239 sb_8__0_.mem_left_track_29.ccff_tail VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold228 net262 VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_38_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_1__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input11_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput119 net119 VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_12
Xoutput108 net108 VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_12
Xoutput90 net90 VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_12
XFILLER_36_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input3_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_input59_A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_3_0_prog_clk net364
+ net144 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_18.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mux_top_track_12.mux_l2_in_0_ sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_12.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout143 net149 VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_8
XFILLER_27_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_ net194 net50 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_154_ sb_8__0_.mux_top_track_2.out VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_10_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__S cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_ clknet_4_4_0_prog_clk
+ net312 net145 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__0_.mux_top_track_38.mux_l1_in_0__A0 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__0_.mux_top_track_24.mux_l2_in_0__175 VGND VGND VPWR VPWR net175 sb_8__0_.mux_top_track_24.mux_l2_in_0__175/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__0_.mux_top_track_0.mux_l1_in_0_ net70 net75 sb_8__0_.mem_top_track_0.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_3_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_3_0_prog_clk net360
+ net145 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_30.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_12.mux_l1_in_1_ net168 net28 sb_8__0_.mem_top_track_12.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_137_ sb_8__0_.mux_top_track_36.out VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_ net43 net32 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__096__A net53 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_left_track_13.mux_l1_in_0__A0 top_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input41_A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_1_0_prog_clk
+ net313 net145 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A0 sb_8__0_.mux_left_track_19.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold229 sb_8__0_.mem_left_track_47.mem_out\[0\] VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold207 sb_8__0_.mem_left_track_7.ccff_tail VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold218 net239 VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__dlymetal6s2s_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X cbx_8__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_1.out sky130_fd_sc_hd__clkbuf_2
XFILLER_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net151 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1__S cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_8_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_8_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold90 net490 VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A0 net42 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_16_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net151 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput109 net109 VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_12
XANTENNA_sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__D net362 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput91 net91 VGND VGND VPWR VPWR chanx_left_out[20] sky130_fd_sc_hd__buf_12
Xoutput80 net80 VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_12
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__A0 net193 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_0__A0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output110_A net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1__CLK clknet_4_15_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_6.mux_l2_in_1__190 VGND VGND VPWR VPWR net190 sb_8__0_.mux_top_track_6.mux_l2_in_1__190/LO
+ sky130_fd_sc_hd__conb_1
XANTENNA_hold186_A net248 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout144 net149 VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_8
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_ net26 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__099__A net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_153_ sb_8__0_.mux_top_track_4.out VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input71_A top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_ VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_38.mux_l1_in_0__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_4_0_prog_clk
+ net315 net145 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_21_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_left_track_3.mux_l2_in_0__155 VGND VGND VPWR VPWR net155 sb_8__0_.mux_left_track_3.mux_l2_in_0__155/LO
+ sky130_fd_sc_hd__conb_1
Xclkbuf_4_10_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_10_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_sb_8__0_.mux_left_track_5.mux_l2_in_0__S sb_8__0_.mem_left_track_5.ccff_tail
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk net372
+ net143 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_30.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_30_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_12.mux_l1_in_0_ top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ net75 sb_8__0_.mem_top_track_12.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_136_ sb_8__0_.mux_top_track_38.out VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_24.mux_l2_in_0_ net175 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_24.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_ sb_8__0_.mux_left_track_29.out net9
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold316_A cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_11_0_prog_clk
+ net404 net148 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_4_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A1 net15 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_input34_A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold208 net241 VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__clkdlybuf4s50_1
X_119_ sb_8__0_.mux_left_track_13.out VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_2
Xhold219 sb_8__0_.mem_top_track_36.ccff_tail VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A1 net4 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_5_0_prog_clk net464
+ net145 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_36.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold80 net485 VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold91 net492 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_31_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold42_A net421 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B net151 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_14_0_prog_clk net332
+ net150 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_29.ccff_tail sky130_fd_sc_hd__dfrtp_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
+ sky130_fd_sc_hd__mux2_1
Xoutput92 net92 VGND VGND VPWR VPWR chanx_left_out[21] sky130_fd_sc_hd__buf_12
Xoutput81 net81 VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_12
Xsb_8__0_.mux_left_track_9.mux_l2_in_0_ net165 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_11.ccff_head VGND VGND VPWR VPWR sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_2.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_0__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_3_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xsb_8__0_.mux_top_track_36.mux_l2_in_0__181 VGND VGND VPWR VPWR net181 sb_8__0_.mux_top_track_36.mux_l2_in_0__181/LO
+ sky130_fd_sc_hd__conb_1
Xsb_8__0_.mux_left_track_31.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_31.out sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_0__A0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout145 net149 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_8
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1__D net348 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_152_ sb_8__0_.mux_top_track_6.out VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dlymetal6s2s_1
Xsb_8__0_.mux_top_track_18.mux_l1_in_1__171 VGND VGND VPWR VPWR net171 sb_8__0_.mux_top_track_18.mux_l1_in_1__171/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_6_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xcbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_0_0_prog_clk
+ net356 net143 VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_input64_A gfpga_pad_io_soc_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__S cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_135_ sb_8__0_.mux_top_track_40.out VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_ sb_8__0_.mux_left_track_17.out net16
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold309_A sb_8__0_.mem_top_track_44.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold211_A sb_8__0_.mem_left_track_11.ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input27_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_118_ sb_8__0_.mux_left_track_15.out VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_2
Xhold209 sb_8__0_.mem_top_track_8.mem_out\[0\] VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__clkdlybuf4s50_1
Xsb_8__0_.mux_left_track_19.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_19.out sky130_fd_sc_hd__clkbuf_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_8_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hold161_A sb_8__0_.mem_top_track_46.ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold70 net469 VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold81 net477 VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_output133_A net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_24.mux_l1_in_0_ net5 net73 sb_8__0_.mem_top_track_24.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold92 net491 VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_5_0_prog_clk net330
+ net145 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_36.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_1 net157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__192 VGND VGND VPWR VPWR net192 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__192/LO
+ sky130_fd_sc_hd__conb_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_36.mux_l2_in_0_ net181 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_top_track_36.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_left_track_13.mux_l2_in_0_ net198 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
+ sb_8__0_.mem_left_track_13.ccff_tail VGND VGND VPWR VPWR sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_13_0_prog_clk net458
+ net150 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_29.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput82 net82 VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_12
Xoutput93 net93 VGND VGND VPWR VPWR chanx_left_out[22] sky130_fd_sc_hd__buf_12
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__S cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_top_track_20.mux_l1_in_0__A0 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xsb_8__0_.mux_left_track_1.mux_l1_in_1__196 VGND VGND VPWR VPWR net196 sb_8__0_.mux_left_track_1.mux_l1_in_1__196/LO
+ sky130_fd_sc_hd__conb_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A1 net24 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
+ VGND VGND VPWR VPWR cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_36_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_0__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout146 net149 VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__buf_2
XFILLER_27_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
+ VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_151_ sb_8__0_.mux_top_track_8.out VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xsb_8__0_.mux_left_track_9.mux_l1_in_0_ top_width_0_height_0_subtile_1__pin_inpad_0_
+ net56 sb_8__0_.mem_left_track_9.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input57_A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR_A
+ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_134_ sb_8__0_.mux_top_track_42.out VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_2
XFILLER_11_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_ sb_8__0_.mux_left_track_11.out net19
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_left_track_47.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__S sb_8__0_.mem_top_track_48.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_117_ sb_8__0_.mux_left_track_17.out VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_2
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output88_A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_1__A0 net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold82 net465 VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_output126_A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold60 net433 VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold93 net497 VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold71 net449 VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_2 net157 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold28_A net367 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_40.mux_l2_in_0__184 VGND VGND VPWR VPWR net184 sb_8__0_.mux_top_track_40.mux_l2_in_0__184/LO
+ sky130_fd_sc_hd__conb_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold271_A sb_8__0_.mem_left_track_11.ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput83 net83 VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_12
Xoutput94 net94 VGND VGND VPWR VPWR chanx_left_out[23] sky130_fd_sc_hd__buf_12
XFILLER_36_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_top_track_20.mux_l1_in_0__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__CLK clknet_4_15_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_7_0_prog_clk clknet_0_prog_clk VGND VGND VPWR VPWR clknet_4_7_0_prog_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail net67
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
Xsb_8__0_.mux_top_track_36.mux_l1_in_0_ net11 net75 sb_8__0_.mem_top_track_36.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X sky130_fd_sc_hd__mux2_1
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold95_A net493 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_left_track_13.mux_l1_in_0_ top_width_0_height_0_subtile_0__pin_inpad_0_
+ net58 sb_8__0_.mem_left_track_13.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__0_.mux_top_track_48.mux_l2_in_0_ sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_top_track_48.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout147 net148 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_4
X_150_ sb_8__0_.mux_top_track_10.out VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__clkbuf_2
XFILLER_23_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_50.mux_l2_in_0_ sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
+ sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X sb_8__0_.mem_left_track_1.ccff_head
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_2_X sky130_fd_sc_hd__mux2_1
Xhold190 net254 VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_2_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_left_track_3.mux_l1_in_0__A0 top_width_0_height_0_subtile_1__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
+ clknet_4_10_0_prog_clk net480 net152 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dfrtp_4
XANTENNA_sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0__D net358 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_133_ sb_8__0_.mux_top_track_44.out VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_2
XANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1__CLK clknet_4_15_0_prog_clk
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__110__A sb_8__0_.mux_left_track_31.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_48.mux_l1_in_1_ net188 net18 sb_8__0_.mem_top_track_48.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xcbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_ sb_8__0_.mux_left_track_5.out net22
+ cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\] VGND VGND VPWR VPWR cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__0_.mux_top_track_50.mux_l1_in_1_ net189 net19 sb_8__0_.mem_top_track_50.mem_out\[0\]
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X sky130_fd_sc_hd__mux2_1
XANTENNA_sb_8__0_.mux_left_track_15.mux_l1_in_0__S sb_8__0_.mem_left_track_15.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_15_0_prog_clk net430
+ net151 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_47.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_31_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_11_0_prog_clk net470
+ net147 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_3.ccff_tail sky130_fd_sc_hd__dfrtp_1
XANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_0__A0 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_116_ sb_8__0_.mux_left_track_19.out VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_2
XANTENNA__105__A net43 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_hold147_A sb_8__0_.mem_left_track_9.mem_out\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_30.out sky130_fd_sc_hd__clkbuf_1
XANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_1__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold314_A cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\] VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold83 net475 VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_output119_A net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold61 net429 VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1__A0 sb_8__0_.mux_left_track_11.out
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold50 net445 VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input32_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold72 net459 VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold94 net494 VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_3 net164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_12_0_prog_clk_A clknet_0_prog_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0__A sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE_TE_B
+ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput84 net84 VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_12
Xoutput95 net95 VGND VGND VPWR VPWR chanx_left_out[24] sky130_fd_sc_hd__buf_12
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__S cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A0 net35 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_31_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xsb_8__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_24.out sky130_fd_sc_hd__clkbuf_1
XFILLER_39_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mux_left_track_31.mux_l2_in_0__A0 net156 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1__D net436 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__113__A net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_hold88_A net489 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_left_track_19.mux_l2_in_0__153 VGND VGND VPWR VPWR net153 sb_8__0_.mux_left_track_19.mux_l2_in_0__153/LO
+ sky130_fd_sc_hd__conb_1
Xfanout148 net149 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_8
XFILLER_27_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold180 net233 VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2__A0 net28 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_18_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_ sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_18.out sky130_fd_sc_hd__clkbuf_2
Xhold191 sb_8__0_.mem_top_track_10.ccff_tail VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_33_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xsb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_9_0_prog_clk net422
+ net148 VGND VGND VPWR VPWR sb_8__0_.mem_top_track_22.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_sb_8__0_.mux_left_track_3.mux_l1_in_0__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B net151 VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xcbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
+ cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail net67
+ VGND VGND VPWR VPWR cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
+ sky130_fd_sc_hd__or2b_2
XANTENNA_hold177_A sb_8__0_.mem_top_track_42.ccff_tail VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_13_0_prog_clk net376
+ net147 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_15.ccff_tail sky130_fd_sc_hd__dfrtp_1
XFILLER_23_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_132_ sb_8__0_.mux_top_track_46.out VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_2
XANTENNA_input62_A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xsb_8__0_.mux_top_track_48.mux_l1_in_0_ top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
+ net73 sb_8__0_.mem_top_track_48.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xsb_8__0_.mux_top_track_50.mux_l1_in_0_ top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
+ net74 sb_8__0_.mem_top_track_50.mem_out\[0\] VGND VGND VPWR VPWR sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
+ sky130_fd_sc_hd__mux2_1
Xsb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_15_0_prog_clk net474
+ net151 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_47.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
Xsb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_ clknet_4_14_0_prog_clk net416
+ net150 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_3.mem_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_0__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_115_ net62 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_2
XFILLER_7_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__121__A sb_8__0_.mux_left_track_9.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_sb_8__0_.mux_left_track_19.mux_l1_in_0__A0 top_width_0_height_0_subtile_3__pin_inpad_0_
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xsb_8__0_.mux_top_track_6.mux_l3_in_0_ sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
+ sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X sb_8__0_.mem_top_track_6.ccff_tail
+ VGND VGND VPWR VPWR sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X sky130_fd_sc_hd__mux2_1
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1__A1 net19 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold40 net391 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold73 net461 VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold95 net493 VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__clkdlybuf4s50_1
Xhold62 net427 VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__clkdlybuf4s50_1
XANTENNA_input25_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold51 net419 VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold84 net479 VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_31_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__116__A sb_8__0_.mux_left_track_19.out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_4 net164 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_0__S sb_8__0_.mem_top_track_44.mem_out\[0\]
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput85 net85 VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_12
Xoutput96 net96 VGND VGND VPWR VPWR chanx_left_out[25] sky130_fd_sc_hd__buf_12
XANTENNA_output131_A net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A1 net11 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xsb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1_ clknet_4_12_0_prog_clk net348
+ net149 VGND VGND VPWR VPWR sb_8__0_.mem_left_track_11.ccff_head sky130_fd_sc_hd__dfrtp_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

