magic
tech sky130A
magscale 1 2
timestamp 1680902775
<< viali >>
rect 13829 54281 13863 54315
rect 18981 54281 19015 54315
rect 2237 54145 2271 54179
rect 4813 54145 4847 54179
rect 7389 54145 7423 54179
rect 9597 54145 9631 54179
rect 12173 54145 12207 54179
rect 14473 54145 14507 54179
rect 15117 54145 15151 54179
rect 15393 54145 15427 54179
rect 17049 54145 17083 54179
rect 17325 54145 17359 54179
rect 17877 54145 17911 54179
rect 18153 54145 18187 54179
rect 19441 54145 19475 54179
rect 20729 54145 20763 54179
rect 21281 54145 21315 54179
rect 22017 54145 22051 54179
rect 22569 54145 22603 54179
rect 23213 54145 23247 54179
rect 23765 54145 23799 54179
rect 24041 54145 24075 54179
rect 24685 54145 24719 54179
rect 2513 54077 2547 54111
rect 5181 54077 5215 54111
rect 7849 54077 7883 54111
rect 9873 54077 9907 54111
rect 12633 54077 12667 54111
rect 19717 54077 19751 54111
rect 14933 54009 14967 54043
rect 17693 54009 17727 54043
rect 22201 54009 22235 54043
rect 14289 53941 14323 53975
rect 16865 53941 16899 53975
rect 20913 53941 20947 53975
rect 23397 53941 23431 53975
rect 24225 53941 24259 53975
rect 25329 53941 25363 53975
rect 24501 53737 24535 53771
rect 24777 53737 24811 53771
rect 2053 53601 2087 53635
rect 4445 53601 4479 53635
rect 7113 53601 7147 53635
rect 11253 53601 11287 53635
rect 1777 53533 1811 53567
rect 4169 53533 4203 53567
rect 6837 53533 6871 53567
rect 10793 53533 10827 53567
rect 22753 53533 22787 53567
rect 23121 53533 23155 53567
rect 23765 53533 23799 53567
rect 25053 53533 25087 53567
rect 23213 53397 23247 53431
rect 23949 53397 23983 53431
rect 25237 53397 25271 53431
rect 5181 53193 5215 53227
rect 5365 53057 5399 53091
rect 23581 53057 23615 53091
rect 24317 53057 24351 53091
rect 25053 53057 25087 53091
rect 25237 52921 25271 52955
rect 23765 52853 23799 52887
rect 24501 52853 24535 52887
rect 6561 52649 6595 52683
rect 24041 52649 24075 52683
rect 6745 52445 6779 52479
rect 24593 52445 24627 52479
rect 25329 52445 25363 52479
rect 24961 52377 24995 52411
rect 24869 52105 24903 52139
rect 25329 51969 25363 52003
rect 25145 51765 25179 51799
rect 8309 51561 8343 51595
rect 9229 51493 9263 51527
rect 7849 51357 7883 51391
rect 8493 51357 8527 51391
rect 9413 51357 9447 51391
rect 7665 51289 7699 51323
rect 24593 51289 24627 51323
rect 24961 51289 24995 51323
rect 25329 51289 25363 51323
rect 24593 50881 24627 50915
rect 24961 50881 24995 50915
rect 25053 50677 25087 50711
rect 7849 50473 7883 50507
rect 9597 50473 9631 50507
rect 8033 50405 8067 50439
rect 8401 50337 8435 50371
rect 7573 50269 7607 50303
rect 9505 50201 9539 50235
rect 25513 50133 25547 50167
rect 24501 49793 24535 49827
rect 24777 49725 24811 49759
rect 10701 49317 10735 49351
rect 11713 49317 11747 49351
rect 10517 49113 10551 49147
rect 11529 49113 11563 49147
rect 24777 49113 24811 49147
rect 25145 49113 25179 49147
rect 25237 49045 25271 49079
rect 6653 48705 6687 48739
rect 6929 48637 6963 48671
rect 8401 48637 8435 48671
rect 8769 48569 8803 48603
rect 8953 48501 8987 48535
rect 25421 48501 25455 48535
rect 10368 48093 10402 48127
rect 23397 48093 23431 48127
rect 25145 48093 25179 48127
rect 25329 48025 25363 48059
rect 10471 47957 10505 47991
rect 24041 47957 24075 47991
rect 9873 47753 9907 47787
rect 10149 47685 10183 47719
rect 9413 47617 9447 47651
rect 24869 47617 24903 47651
rect 25329 47617 25363 47651
rect 9505 47413 9539 47447
rect 25145 47413 25179 47447
rect 11656 47005 11690 47039
rect 11759 46937 11793 46971
rect 25421 46869 25455 46903
rect 10793 46665 10827 46699
rect 11069 46665 11103 46699
rect 14105 46597 14139 46631
rect 10333 46529 10367 46563
rect 12576 46529 12610 46563
rect 13921 46529 13955 46563
rect 25329 46529 25363 46563
rect 15761 46461 15795 46495
rect 10425 46325 10459 46359
rect 12679 46325 12713 46359
rect 25145 46325 25179 46359
rect 8493 46121 8527 46155
rect 8125 45985 8159 46019
rect 14841 45985 14875 46019
rect 15025 45985 15059 46019
rect 16497 45985 16531 46019
rect 7941 45917 7975 45951
rect 13312 45917 13346 45951
rect 24869 45917 24903 45951
rect 25329 45917 25363 45951
rect 13415 45781 13449 45815
rect 25145 45781 25179 45815
rect 12909 45509 12943 45543
rect 12725 45441 12759 45475
rect 14565 45373 14599 45407
rect 25421 45237 25455 45271
rect 10885 45033 10919 45067
rect 15669 44897 15703 44931
rect 9137 44829 9171 44863
rect 25329 44829 25363 44863
rect 9413 44761 9447 44795
rect 11253 44761 11287 44795
rect 15853 44761 15887 44795
rect 17509 44761 17543 44795
rect 11437 44693 11471 44727
rect 25145 44693 25179 44727
rect 9597 44489 9631 44523
rect 9137 44353 9171 44387
rect 10609 44353 10643 44387
rect 11529 44353 11563 44387
rect 24777 44353 24811 44387
rect 25145 44353 25179 44387
rect 8953 44285 8987 44319
rect 10701 44149 10735 44183
rect 11069 44149 11103 44183
rect 25237 44149 25271 44183
rect 22109 43945 22143 43979
rect 20637 43809 20671 43843
rect 20361 43741 20395 43775
rect 22385 43673 22419 43707
rect 25513 43605 25547 43639
rect 25145 43333 25179 43367
rect 25237 43061 25271 43095
rect 10241 42721 10275 42755
rect 9597 42653 9631 42687
rect 9781 42653 9815 42687
rect 24777 42585 24811 42619
rect 25145 42585 25179 42619
rect 25237 42517 25271 42551
rect 11161 42313 11195 42347
rect 9413 42109 9447 42143
rect 9689 42109 9723 42143
rect 11529 41973 11563 42007
rect 11713 41973 11747 42007
rect 25421 41973 25455 42007
rect 10885 41769 10919 41803
rect 10425 41633 10459 41667
rect 10241 41565 10275 41599
rect 25145 41565 25179 41599
rect 25329 41497 25363 41531
rect 24869 41089 24903 41123
rect 25329 41089 25363 41123
rect 25145 40885 25179 40919
rect 25513 40341 25547 40375
rect 25145 40137 25179 40171
rect 25329 40001 25363 40035
rect 24869 39389 24903 39423
rect 25329 39389 25363 39423
rect 25145 39253 25179 39287
rect 25421 38709 25455 38743
rect 25329 38301 25363 38335
rect 25145 38165 25179 38199
rect 8677 37961 8711 37995
rect 8861 37825 8895 37859
rect 24777 37825 24811 37859
rect 25145 37825 25179 37859
rect 25329 37689 25363 37723
rect 25513 37077 25547 37111
rect 25145 36805 25179 36839
rect 25329 36601 25363 36635
rect 24869 36125 24903 36159
rect 25329 36125 25363 36159
rect 25145 35989 25179 36023
rect 22477 35785 22511 35819
rect 11529 35717 11563 35751
rect 21189 35717 21223 35751
rect 9413 35649 9447 35683
rect 21097 35649 21131 35683
rect 22385 35649 22419 35683
rect 9689 35581 9723 35615
rect 11161 35581 11195 35615
rect 21281 35581 21315 35615
rect 22569 35581 22603 35615
rect 11805 35445 11839 35479
rect 20361 35445 20395 35479
rect 20729 35445 20763 35479
rect 22017 35445 22051 35479
rect 25421 35445 25455 35479
rect 23305 35105 23339 35139
rect 23213 35037 23247 35071
rect 25329 35037 25363 35071
rect 22385 34969 22419 35003
rect 23121 34969 23155 35003
rect 21833 34901 21867 34935
rect 22753 34901 22787 34935
rect 25145 34901 25179 34935
rect 25145 34697 25179 34731
rect 24869 34561 24903 34595
rect 25329 34561 25363 34595
rect 21373 34357 21407 34391
rect 9137 34153 9171 34187
rect 15393 34017 15427 34051
rect 21649 34017 21683 34051
rect 9321 33949 9355 33983
rect 19441 33949 19475 33983
rect 24869 33949 24903 33983
rect 25329 33949 25363 33983
rect 14657 33881 14691 33915
rect 15853 33881 15887 33915
rect 19717 33881 19751 33915
rect 21925 33881 21959 33915
rect 21189 33813 21223 33847
rect 23397 33813 23431 33847
rect 23673 33813 23707 33847
rect 25145 33813 25179 33847
rect 19809 33541 19843 33575
rect 19533 33473 19567 33507
rect 22017 33473 22051 33507
rect 25329 33473 25363 33507
rect 21281 33405 21315 33439
rect 22293 33405 22327 33439
rect 23765 33405 23799 33439
rect 21557 33269 21591 33303
rect 24133 33269 24167 33303
rect 24317 33269 24351 33303
rect 24593 33269 24627 33303
rect 24869 33269 24903 33303
rect 25145 33269 25179 33303
rect 16773 33065 16807 33099
rect 24041 33065 24075 33099
rect 16129 32929 16163 32963
rect 16589 32929 16623 32963
rect 17049 32929 17083 32963
rect 22293 32929 22327 32963
rect 22569 32929 22603 32963
rect 25053 32929 25087 32963
rect 25237 32929 25271 32963
rect 16037 32861 16071 32895
rect 20637 32861 20671 32895
rect 15945 32793 15979 32827
rect 19901 32793 19935 32827
rect 15577 32725 15611 32759
rect 19625 32725 19659 32759
rect 24593 32725 24627 32759
rect 24961 32725 24995 32759
rect 17049 32521 17083 32555
rect 25237 32521 25271 32555
rect 15393 32453 15427 32487
rect 16865 32453 16899 32487
rect 22845 32453 22879 32487
rect 22109 32385 22143 32419
rect 23489 32385 23523 32419
rect 16129 32317 16163 32351
rect 19073 32317 19107 32351
rect 19349 32317 19383 32351
rect 23765 32317 23799 32351
rect 20821 32181 20855 32215
rect 21189 32181 21223 32215
rect 21649 32181 21683 32215
rect 17036 31977 17070 32011
rect 22661 31977 22695 32011
rect 15577 31909 15611 31943
rect 23029 31909 23063 31943
rect 25145 31909 25179 31943
rect 16129 31841 16163 31875
rect 18521 31841 18555 31875
rect 19717 31841 19751 31875
rect 22109 31841 22143 31875
rect 22201 31841 22235 31875
rect 23489 31841 23523 31875
rect 23581 31841 23615 31875
rect 16037 31773 16071 31807
rect 16773 31773 16807 31807
rect 19441 31773 19475 31807
rect 24869 31773 24903 31807
rect 25329 31773 25363 31807
rect 23397 31705 23431 31739
rect 15945 31637 15979 31671
rect 18889 31637 18923 31671
rect 21189 31637 21223 31671
rect 21649 31637 21683 31671
rect 22017 31637 22051 31671
rect 24685 31637 24719 31671
rect 15761 31433 15795 31467
rect 19165 31433 19199 31467
rect 21373 31433 21407 31467
rect 21557 31433 21591 31467
rect 24225 31433 24259 31467
rect 19533 31365 19567 31399
rect 22753 31365 22787 31399
rect 17417 31297 17451 31331
rect 20453 31297 20487 31331
rect 20545 31297 20579 31331
rect 22477 31297 22511 31331
rect 25329 31297 25363 31331
rect 13369 31229 13403 31263
rect 13645 31229 13679 31263
rect 15485 31229 15519 31263
rect 16405 31229 16439 31263
rect 17693 31229 17727 31263
rect 20637 31229 20671 31263
rect 20085 31161 20119 31195
rect 15117 31093 15151 31127
rect 16773 31093 16807 31127
rect 19809 31093 19843 31127
rect 24593 31093 24627 31127
rect 25145 31093 25179 31127
rect 9137 30889 9171 30923
rect 15577 30889 15611 30923
rect 15761 30889 15795 30923
rect 18521 30889 18555 30923
rect 18889 30889 18923 30923
rect 22477 30889 22511 30923
rect 22845 30889 22879 30923
rect 25513 30889 25547 30923
rect 16773 30753 16807 30787
rect 20729 30753 20763 30787
rect 9321 30685 9355 30719
rect 14381 30685 14415 30719
rect 15117 30617 15151 30651
rect 17049 30617 17083 30651
rect 21005 30617 21039 30651
rect 24593 30617 24627 30651
rect 20085 30549 20119 30583
rect 15945 30345 15979 30379
rect 16773 30345 16807 30379
rect 18981 30345 19015 30379
rect 20269 30345 20303 30379
rect 14105 30277 14139 30311
rect 20361 30277 20395 30311
rect 22477 30277 22511 30311
rect 9137 30209 9171 30243
rect 11805 30209 11839 30243
rect 15853 30209 15887 30243
rect 16865 30209 16899 30243
rect 21281 30209 21315 30243
rect 22385 30209 22419 30243
rect 12081 30141 12115 30175
rect 14841 30141 14875 30175
rect 16037 30141 16071 30175
rect 20545 30141 20579 30175
rect 22661 30141 22695 30175
rect 23305 30141 23339 30175
rect 23581 30141 23615 30175
rect 25053 30141 25087 30175
rect 8953 30073 8987 30107
rect 13553 30005 13587 30039
rect 15485 30005 15519 30039
rect 19901 30005 19935 30039
rect 22017 30005 22051 30039
rect 25329 30005 25363 30039
rect 13461 29801 13495 29835
rect 16313 29801 16347 29835
rect 23857 29801 23891 29835
rect 12909 29733 12943 29767
rect 16497 29733 16531 29767
rect 20177 29733 20211 29767
rect 25145 29733 25179 29767
rect 11161 29665 11195 29699
rect 15853 29665 15887 29699
rect 17049 29665 17083 29699
rect 20729 29665 20763 29699
rect 15577 29597 15611 29631
rect 20637 29597 20671 29631
rect 23397 29597 23431 29631
rect 24041 29597 24075 29631
rect 25329 29597 25363 29631
rect 11437 29529 11471 29563
rect 17325 29529 17359 29563
rect 22937 29529 22971 29563
rect 13277 29461 13311 29495
rect 13737 29461 13771 29495
rect 15209 29461 15243 29495
rect 15669 29461 15703 29495
rect 18797 29461 18831 29495
rect 19441 29461 19475 29495
rect 20545 29461 20579 29495
rect 23213 29461 23247 29495
rect 24501 29461 24535 29495
rect 24777 29461 24811 29495
rect 9505 29257 9539 29291
rect 9873 29257 9907 29291
rect 12541 29257 12575 29291
rect 12633 29257 12667 29291
rect 15117 29257 15151 29291
rect 16037 29257 16071 29291
rect 17233 29257 17267 29291
rect 18061 29257 18095 29291
rect 19165 29257 19199 29291
rect 19257 29257 19291 29291
rect 23949 29257 23983 29291
rect 25421 29257 25455 29291
rect 15945 29189 15979 29223
rect 17325 29189 17359 29223
rect 17969 29189 18003 29223
rect 19993 29189 20027 29223
rect 13369 29121 13403 29155
rect 22201 29121 22235 29155
rect 24041 29121 24075 29155
rect 25329 29121 25363 29155
rect 9965 29053 9999 29087
rect 10057 29053 10091 29087
rect 12817 29053 12851 29087
rect 16129 29053 16163 29087
rect 17509 29053 17543 29087
rect 19441 29053 19475 29087
rect 22937 29053 22971 29087
rect 24133 29053 24167 29087
rect 24777 29053 24811 29087
rect 12173 28985 12207 29019
rect 15577 28985 15611 29019
rect 16865 28985 16899 29019
rect 18797 28985 18831 29019
rect 21833 28985 21867 29019
rect 23581 28985 23615 29019
rect 13632 28917 13666 28951
rect 10885 28713 10919 28747
rect 13553 28713 13587 28747
rect 15853 28713 15887 28747
rect 18889 28713 18923 28747
rect 22385 28713 22419 28747
rect 22845 28645 22879 28679
rect 9137 28577 9171 28611
rect 11437 28577 11471 28611
rect 13185 28577 13219 28611
rect 15301 28577 15335 28611
rect 15393 28577 15427 28611
rect 17417 28577 17451 28611
rect 20085 28577 20119 28611
rect 23397 28577 23431 28611
rect 25053 28577 25087 28611
rect 25237 28577 25271 28611
rect 17141 28509 17175 28543
rect 20637 28509 20671 28543
rect 23213 28509 23247 28543
rect 24041 28509 24075 28543
rect 24961 28509 24995 28543
rect 9413 28441 9447 28475
rect 11713 28441 11747 28475
rect 15209 28441 15243 28475
rect 20913 28441 20947 28475
rect 23305 28441 23339 28475
rect 14841 28373 14875 28407
rect 16037 28373 16071 28407
rect 16221 28373 16255 28407
rect 19441 28373 19475 28407
rect 19809 28373 19843 28407
rect 19901 28373 19935 28407
rect 23949 28373 23983 28407
rect 24593 28373 24627 28407
rect 11069 28169 11103 28203
rect 13737 28169 13771 28203
rect 15577 28169 15611 28203
rect 16405 28169 16439 28203
rect 18981 28169 19015 28203
rect 19717 28169 19751 28203
rect 21557 28169 21591 28203
rect 22385 28169 22419 28203
rect 22477 28169 22511 28203
rect 11989 28101 12023 28135
rect 21097 28101 21131 28135
rect 15669 28033 15703 28067
rect 17233 28033 17267 28067
rect 20361 28033 20395 28067
rect 11713 27965 11747 27999
rect 15761 27965 15795 27999
rect 17325 27965 17359 27999
rect 17417 27965 17451 27999
rect 18061 27965 18095 27999
rect 22569 27965 22603 27999
rect 23213 27965 23247 27999
rect 23489 27965 23523 27999
rect 19349 27897 19383 27931
rect 22017 27897 22051 27931
rect 13461 27829 13495 27863
rect 15209 27829 15243 27863
rect 16313 27829 16347 27863
rect 16865 27829 16899 27863
rect 18521 27829 18555 27863
rect 18797 27829 18831 27863
rect 24961 27829 24995 27863
rect 25237 27829 25271 27863
rect 25421 27829 25455 27863
rect 12633 27625 12667 27659
rect 20164 27625 20198 27659
rect 23857 27625 23891 27659
rect 17509 27557 17543 27591
rect 10517 27489 10551 27523
rect 10793 27489 10827 27523
rect 13553 27489 13587 27523
rect 15761 27489 15795 27523
rect 18061 27489 18095 27523
rect 19901 27489 19935 27523
rect 22109 27489 22143 27523
rect 24133 27489 24167 27523
rect 25053 27489 25087 27523
rect 25145 27489 25179 27523
rect 13461 27421 13495 27455
rect 17877 27421 17911 27455
rect 24961 27421 24995 27455
rect 13369 27353 13403 27387
rect 16221 27353 16255 27387
rect 22385 27353 22419 27387
rect 12265 27285 12299 27319
rect 13001 27285 13035 27319
rect 15209 27285 15243 27319
rect 15577 27285 15611 27319
rect 15669 27285 15703 27319
rect 16497 27285 16531 27319
rect 17969 27285 18003 27319
rect 21649 27285 21683 27319
rect 24593 27285 24627 27319
rect 15669 27081 15703 27115
rect 19993 27081 20027 27115
rect 22845 27081 22879 27115
rect 25329 27081 25363 27115
rect 11621 27013 11655 27047
rect 13369 27013 13403 27047
rect 15761 27013 15795 27047
rect 9321 26945 9355 26979
rect 13093 26945 13127 26979
rect 17969 26945 18003 26979
rect 22753 26945 22787 26979
rect 23581 26945 23615 26979
rect 9597 26877 9631 26911
rect 11069 26877 11103 26911
rect 15853 26877 15887 26911
rect 18245 26877 18279 26911
rect 23029 26877 23063 26911
rect 23857 26877 23891 26911
rect 14841 26741 14875 26775
rect 15301 26741 15335 26775
rect 19717 26741 19751 26775
rect 21833 26741 21867 26775
rect 22385 26741 22419 26775
rect 11161 26537 11195 26571
rect 15669 26537 15703 26571
rect 17233 26537 17267 26571
rect 21189 26537 21223 26571
rect 22293 26537 22327 26571
rect 23857 26537 23891 26571
rect 14289 26469 14323 26503
rect 21465 26469 21499 26503
rect 22661 26469 22695 26503
rect 24593 26469 24627 26503
rect 9137 26401 9171 26435
rect 10885 26401 10919 26435
rect 14933 26401 14967 26435
rect 15301 26401 15335 26435
rect 16221 26401 16255 26435
rect 16681 26401 16715 26435
rect 19441 26401 19475 26435
rect 19717 26401 19751 26435
rect 23213 26401 23247 26435
rect 25237 26401 25271 26435
rect 16865 26333 16899 26367
rect 17141 26333 17175 26367
rect 23029 26333 23063 26367
rect 23121 26333 23155 26367
rect 24041 26333 24075 26367
rect 24961 26333 24995 26367
rect 25053 26333 25087 26367
rect 9413 26265 9447 26299
rect 11345 26265 11379 26299
rect 14657 26265 14691 26299
rect 14749 26265 14783 26299
rect 16037 26265 16071 26299
rect 16129 26265 16163 26299
rect 18245 26197 18279 26231
rect 12633 25993 12667 26027
rect 14013 25993 14047 26027
rect 14841 25993 14875 26027
rect 15301 25993 15335 26027
rect 17785 25993 17819 26027
rect 18153 25993 18187 26027
rect 19165 25993 19199 26027
rect 22477 25993 22511 26027
rect 13921 25925 13955 25959
rect 17417 25925 17451 25959
rect 18245 25925 18279 25959
rect 12541 25857 12575 25891
rect 15209 25857 15243 25891
rect 16037 25857 16071 25891
rect 17049 25857 17083 25891
rect 22385 25857 22419 25891
rect 23489 25857 23523 25891
rect 23949 25857 23983 25891
rect 12725 25789 12759 25823
rect 14105 25789 14139 25823
rect 15393 25789 15427 25823
rect 18429 25789 18463 25823
rect 22661 25789 22695 25823
rect 25145 25789 25179 25823
rect 13553 25721 13587 25755
rect 12173 25653 12207 25687
rect 16865 25653 16899 25687
rect 21557 25653 21591 25687
rect 22017 25653 22051 25687
rect 23305 25653 23339 25687
rect 14289 25449 14323 25483
rect 18337 25449 18371 25483
rect 20269 25449 20303 25483
rect 21557 25449 21591 25483
rect 24593 25449 24627 25483
rect 12909 25381 12943 25415
rect 16957 25381 16991 25415
rect 24501 25381 24535 25415
rect 25145 25381 25179 25415
rect 10885 25313 10919 25347
rect 11161 25313 11195 25347
rect 14749 25313 14783 25347
rect 14841 25313 14875 25347
rect 16313 25313 16347 25347
rect 17141 25245 17175 25279
rect 17785 25245 17819 25279
rect 18153 25245 18187 25279
rect 19809 25245 19843 25279
rect 21005 25245 21039 25279
rect 21741 25245 21775 25279
rect 22661 25245 22695 25279
rect 25329 25245 25363 25279
rect 15301 25177 15335 25211
rect 16129 25177 16163 25211
rect 19349 25177 19383 25211
rect 23857 25177 23891 25211
rect 24869 25177 24903 25211
rect 12633 25109 12667 25143
rect 14657 25109 14691 25143
rect 15761 25109 15795 25143
rect 16221 25109 16255 25143
rect 17601 25109 17635 25143
rect 18705 25109 18739 25143
rect 19901 25109 19935 25143
rect 20821 25109 20855 25143
rect 15117 24905 15151 24939
rect 18429 24905 18463 24939
rect 12081 24837 12115 24871
rect 15393 24837 15427 24871
rect 17233 24837 17267 24871
rect 18521 24837 18555 24871
rect 22477 24837 22511 24871
rect 12173 24769 12207 24803
rect 13001 24769 13035 24803
rect 17325 24769 17359 24803
rect 19073 24769 19107 24803
rect 19717 24769 19751 24803
rect 23581 24769 23615 24803
rect 9413 24701 9447 24735
rect 9689 24701 9723 24735
rect 12265 24701 12299 24735
rect 13277 24701 13311 24735
rect 14749 24701 14783 24735
rect 17417 24701 17451 24735
rect 18613 24701 18647 24735
rect 19993 24701 20027 24735
rect 21465 24701 21499 24735
rect 22569 24701 22603 24735
rect 22661 24701 22695 24735
rect 23857 24701 23891 24735
rect 11161 24565 11195 24599
rect 11713 24565 11747 24599
rect 15485 24565 15519 24599
rect 16865 24565 16899 24599
rect 18061 24565 18095 24599
rect 19349 24565 19383 24599
rect 22109 24565 22143 24599
rect 25329 24565 25363 24599
rect 14197 24361 14231 24395
rect 21189 24361 21223 24395
rect 25329 24361 25363 24395
rect 25513 24361 25547 24395
rect 18153 24293 18187 24327
rect 21557 24293 21591 24327
rect 25145 24293 25179 24327
rect 9413 24225 9447 24259
rect 11989 24225 12023 24259
rect 18797 24225 18831 24259
rect 19441 24225 19475 24259
rect 21925 24225 21959 24259
rect 24593 24225 24627 24259
rect 9137 24157 9171 24191
rect 17693 24157 17727 24191
rect 18521 24157 18555 24191
rect 18613 24157 18647 24191
rect 11253 24089 11287 24123
rect 11437 24089 11471 24123
rect 12265 24089 12299 24123
rect 15945 24089 15979 24123
rect 19717 24089 19751 24123
rect 22201 24089 22235 24123
rect 10885 24021 10919 24055
rect 13737 24021 13771 24055
rect 23673 24021 23707 24055
rect 24041 24021 24075 24055
rect 9781 23817 9815 23851
rect 10425 23817 10459 23851
rect 10793 23817 10827 23851
rect 14933 23817 14967 23851
rect 17233 23817 17267 23851
rect 17325 23817 17359 23851
rect 18061 23817 18095 23851
rect 18613 23817 18647 23851
rect 18889 23817 18923 23851
rect 24961 23817 24995 23851
rect 25421 23817 25455 23851
rect 13645 23749 13679 23783
rect 13737 23749 13771 23783
rect 25329 23749 25363 23783
rect 8033 23681 8067 23715
rect 14841 23681 14875 23715
rect 18245 23681 18279 23715
rect 19625 23681 19659 23715
rect 19717 23681 19751 23715
rect 20821 23681 20855 23715
rect 20913 23681 20947 23715
rect 21465 23681 21499 23715
rect 22385 23681 22419 23715
rect 23213 23681 23247 23715
rect 8309 23613 8343 23647
rect 10885 23613 10919 23647
rect 10977 23613 11011 23647
rect 13829 23613 13863 23647
rect 15025 23613 15059 23647
rect 15669 23613 15703 23647
rect 17417 23613 17451 23647
rect 19901 23613 19935 23647
rect 21005 23613 21039 23647
rect 23489 23613 23523 23647
rect 14473 23545 14507 23579
rect 10057 23477 10091 23511
rect 13277 23477 13311 23511
rect 16865 23477 16899 23511
rect 18797 23477 18831 23511
rect 19257 23477 19291 23511
rect 20453 23477 20487 23511
rect 22201 23477 22235 23511
rect 9137 23273 9171 23307
rect 15853 23273 15887 23307
rect 18981 23273 19015 23307
rect 14749 23205 14783 23239
rect 17877 23205 17911 23239
rect 9689 23137 9723 23171
rect 10241 23137 10275 23171
rect 11713 23137 11747 23171
rect 11805 23137 11839 23171
rect 13553 23137 13587 23171
rect 15301 23137 15335 23171
rect 18429 23137 18463 23171
rect 20177 23137 20211 23171
rect 20729 23137 20763 23171
rect 25053 23137 25087 23171
rect 25237 23137 25271 23171
rect 9597 23069 9631 23103
rect 11621 23069 11655 23103
rect 13369 23069 13403 23103
rect 15117 23069 15151 23103
rect 18245 23069 18279 23103
rect 19901 23069 19935 23103
rect 19993 23069 20027 23103
rect 21833 23069 21867 23103
rect 22845 23069 22879 23103
rect 24961 23069 24995 23103
rect 9505 23001 9539 23035
rect 14473 23001 14507 23035
rect 15209 23001 15243 23035
rect 23857 23001 23891 23035
rect 11253 22933 11287 22967
rect 13001 22933 13035 22967
rect 13461 22933 13495 22967
rect 14197 22933 14231 22967
rect 18337 22933 18371 22967
rect 19533 22933 19567 22967
rect 21649 22933 21683 22967
rect 24593 22933 24627 22967
rect 14473 22729 14507 22763
rect 16865 22729 16899 22763
rect 18705 22729 18739 22763
rect 19717 22729 19751 22763
rect 21189 22729 21223 22763
rect 14565 22661 14599 22695
rect 8125 22593 8159 22627
rect 10149 22593 10183 22627
rect 12357 22593 12391 22627
rect 17049 22593 17083 22627
rect 18889 22593 18923 22627
rect 21097 22593 21131 22627
rect 22109 22593 22143 22627
rect 23949 22593 23983 22627
rect 8401 22525 8435 22559
rect 12633 22525 12667 22559
rect 21281 22525 21315 22559
rect 23305 22525 23339 22559
rect 24777 22525 24811 22559
rect 20361 22457 20395 22491
rect 9873 22389 9907 22423
rect 14105 22389 14139 22423
rect 20729 22389 20763 22423
rect 11989 22185 12023 22219
rect 23305 22185 23339 22219
rect 23765 22185 23799 22219
rect 11345 22049 11379 22083
rect 12633 22049 12667 22083
rect 15301 22049 15335 22083
rect 15485 22049 15519 22083
rect 18153 22049 18187 22083
rect 20361 22049 20395 22083
rect 21557 22049 21591 22083
rect 25053 22049 25087 22083
rect 25237 22049 25271 22083
rect 12449 21981 12483 22015
rect 16129 21981 16163 22015
rect 23949 21981 23983 22015
rect 24961 21981 24995 22015
rect 11161 21913 11195 21947
rect 16405 21913 16439 21947
rect 21833 21913 21867 21947
rect 8953 21845 8987 21879
rect 10333 21845 10367 21879
rect 10701 21845 10735 21879
rect 11069 21845 11103 21879
rect 12357 21845 12391 21879
rect 14841 21845 14875 21879
rect 15209 21845 15243 21879
rect 17877 21845 17911 21879
rect 19717 21845 19751 21879
rect 20085 21845 20119 21879
rect 20177 21845 20211 21879
rect 20913 21845 20947 21879
rect 24593 21845 24627 21879
rect 10425 21641 10459 21675
rect 11713 21641 11747 21675
rect 21373 21641 21407 21675
rect 21557 21641 21591 21675
rect 22477 21641 22511 21675
rect 25329 21641 25363 21675
rect 9689 21573 9723 21607
rect 10885 21573 10919 21607
rect 15669 21573 15703 21607
rect 21189 21573 21223 21607
rect 9597 21505 9631 21539
rect 10793 21505 10827 21539
rect 18889 21505 18923 21539
rect 19901 21505 19935 21539
rect 20729 21505 20763 21539
rect 22385 21505 22419 21539
rect 23305 21505 23339 21539
rect 6929 21437 6963 21471
rect 7205 21437 7239 21471
rect 9781 21437 9815 21471
rect 10977 21437 11011 21471
rect 13093 21437 13127 21471
rect 13369 21437 13403 21471
rect 19993 21437 20027 21471
rect 20177 21437 20211 21471
rect 22661 21437 22695 21471
rect 23581 21437 23615 21471
rect 9229 21369 9263 21403
rect 15853 21369 15887 21403
rect 18705 21369 18739 21403
rect 8677 21301 8711 21335
rect 14841 21301 14875 21335
rect 15117 21301 15151 21335
rect 19165 21301 19199 21335
rect 19533 21301 19567 21335
rect 22017 21301 22051 21335
rect 25053 21301 25087 21335
rect 21465 21097 21499 21131
rect 12449 21029 12483 21063
rect 20821 21029 20855 21063
rect 9965 20961 9999 20995
rect 15209 20961 15243 20995
rect 19993 20961 20027 20995
rect 22017 20961 22051 20995
rect 23857 20961 23891 20995
rect 25053 20961 25087 20995
rect 25145 20961 25179 20995
rect 10701 20893 10735 20927
rect 19901 20893 19935 20927
rect 21005 20893 21039 20927
rect 22661 20893 22695 20927
rect 10977 20825 11011 20859
rect 12725 20825 12759 20859
rect 14565 20825 14599 20859
rect 15485 20825 15519 20859
rect 19809 20825 19843 20859
rect 21281 20825 21315 20859
rect 9045 20757 9079 20791
rect 16957 20757 16991 20791
rect 17233 20757 17267 20791
rect 18705 20757 18739 20791
rect 19441 20757 19475 20791
rect 20453 20757 20487 20791
rect 24593 20757 24627 20791
rect 24961 20757 24995 20791
rect 10425 20553 10459 20587
rect 10793 20553 10827 20587
rect 15393 20553 15427 20587
rect 15485 20553 15519 20587
rect 20821 20553 20855 20587
rect 20913 20553 20947 20587
rect 25329 20553 25363 20587
rect 8033 20485 8067 20519
rect 17141 20485 17175 20519
rect 21465 20485 21499 20519
rect 16865 20417 16899 20451
rect 19257 20417 19291 20451
rect 19901 20417 19935 20451
rect 22201 20417 22235 20451
rect 22937 20417 22971 20451
rect 7757 20349 7791 20383
rect 9781 20349 9815 20383
rect 10885 20349 10919 20383
rect 10977 20349 11011 20383
rect 12725 20349 12759 20383
rect 13001 20349 13035 20383
rect 15577 20349 15611 20383
rect 21097 20349 21131 20383
rect 23581 20349 23615 20383
rect 23857 20349 23891 20383
rect 22017 20281 22051 20315
rect 10149 20213 10183 20247
rect 14473 20213 14507 20247
rect 15025 20213 15059 20247
rect 18613 20213 18647 20247
rect 19073 20213 19107 20247
rect 19717 20213 19751 20247
rect 20453 20213 20487 20247
rect 22753 20213 22787 20247
rect 8493 20009 8527 20043
rect 11345 20009 11379 20043
rect 16037 20009 16071 20043
rect 16497 20009 16531 20043
rect 23857 20009 23891 20043
rect 9137 19873 9171 19907
rect 11989 19873 12023 19907
rect 14565 19873 14599 19907
rect 17969 19873 18003 19907
rect 18061 19873 18095 19907
rect 19901 19873 19935 19907
rect 22109 19873 22143 19907
rect 14289 19805 14323 19839
rect 16681 19805 16715 19839
rect 18889 19805 18923 19839
rect 9413 19737 9447 19771
rect 11805 19737 11839 19771
rect 17877 19737 17911 19771
rect 20177 19737 20211 19771
rect 22385 19737 22419 19771
rect 24133 19737 24167 19771
rect 25421 19737 25455 19771
rect 10885 19669 10919 19703
rect 11713 19669 11747 19703
rect 16957 19669 16991 19703
rect 17509 19669 17543 19703
rect 18705 19669 18739 19703
rect 21649 19669 21683 19703
rect 24409 19669 24443 19703
rect 8769 19465 8803 19499
rect 11713 19465 11747 19499
rect 16865 19465 16899 19499
rect 17325 19465 17359 19499
rect 18981 19465 19015 19499
rect 20453 19465 20487 19499
rect 20545 19465 20579 19499
rect 22661 19465 22695 19499
rect 25145 19465 25179 19499
rect 25421 19465 25455 19499
rect 23673 19397 23707 19431
rect 9137 19329 9171 19363
rect 9229 19329 9263 19363
rect 15209 19329 15243 19363
rect 16129 19329 16163 19363
rect 17233 19329 17267 19363
rect 19165 19329 19199 19363
rect 21281 19329 21315 19363
rect 22569 19329 22603 19363
rect 23397 19329 23431 19363
rect 6561 19261 6595 19295
rect 6837 19261 6871 19295
rect 9321 19261 9355 19295
rect 11161 19261 11195 19295
rect 12541 19261 12575 19295
rect 12817 19261 12851 19295
rect 17417 19261 17451 19295
rect 20729 19261 20763 19295
rect 22753 19261 22787 19295
rect 11069 19193 11103 19227
rect 15945 19193 15979 19227
rect 20085 19193 20119 19227
rect 21833 19193 21867 19227
rect 22201 19193 22235 19227
rect 8309 19125 8343 19159
rect 14289 19125 14323 19159
rect 14657 19125 14691 19159
rect 15025 19125 15059 19159
rect 10057 18921 10091 18955
rect 12725 18921 12759 18955
rect 25237 18921 25271 18955
rect 11529 18853 11563 18887
rect 6929 18785 6963 18819
rect 10609 18785 10643 18819
rect 12081 18785 12115 18819
rect 13277 18785 13311 18819
rect 17509 18785 17543 18819
rect 23857 18785 23891 18819
rect 6653 18717 6687 18751
rect 9689 18717 9723 18751
rect 10425 18717 10459 18751
rect 11069 18717 11103 18751
rect 11989 18717 12023 18751
rect 17233 18717 17267 18751
rect 17877 18717 17911 18751
rect 21465 18717 21499 18751
rect 22201 18717 22235 18751
rect 22753 18717 22787 18751
rect 24685 18717 24719 18751
rect 8769 18649 8803 18683
rect 24869 18649 24903 18683
rect 8401 18581 8435 18615
rect 10517 18581 10551 18615
rect 11897 18581 11931 18615
rect 13093 18581 13127 18615
rect 13185 18581 13219 18615
rect 13829 18581 13863 18615
rect 14289 18581 14323 18615
rect 16865 18581 16899 18615
rect 17325 18581 17359 18615
rect 18061 18581 18095 18615
rect 21281 18581 21315 18615
rect 22017 18581 22051 18615
rect 9505 18377 9539 18411
rect 9965 18377 9999 18411
rect 10425 18377 10459 18411
rect 14289 18377 14323 18411
rect 14933 18377 14967 18411
rect 14197 18309 14231 18343
rect 23305 18309 23339 18343
rect 10333 18241 10367 18275
rect 11253 18241 11287 18275
rect 12449 18241 12483 18275
rect 16865 18241 16899 18275
rect 21281 18241 21315 18275
rect 22109 18241 22143 18275
rect 23949 18241 23983 18275
rect 7757 18173 7791 18207
rect 8033 18173 8067 18207
rect 10609 18173 10643 18207
rect 13185 18173 13219 18207
rect 14381 18173 14415 18207
rect 17141 18173 17175 18207
rect 24685 18173 24719 18207
rect 13829 18105 13863 18139
rect 18981 18105 19015 18139
rect 11069 18037 11103 18071
rect 18613 18037 18647 18071
rect 21097 18037 21131 18071
rect 7849 17833 7883 17867
rect 12265 17833 12299 17867
rect 20637 17765 20671 17799
rect 8401 17697 8435 17731
rect 11805 17697 11839 17731
rect 12725 17697 12759 17731
rect 12909 17697 12943 17731
rect 16129 17697 16163 17731
rect 17969 17697 18003 17731
rect 19901 17697 19935 17731
rect 19993 17697 20027 17731
rect 23857 17697 23891 17731
rect 25053 17697 25087 17731
rect 25145 17697 25179 17731
rect 9781 17629 9815 17663
rect 12633 17629 12667 17663
rect 16405 17629 16439 17663
rect 18429 17629 18463 17663
rect 20821 17629 20855 17663
rect 21465 17629 21499 17663
rect 22845 17629 22879 17663
rect 8217 17561 8251 17595
rect 10057 17561 10091 17595
rect 14197 17561 14231 17595
rect 17785 17561 17819 17595
rect 18797 17561 18831 17595
rect 22017 17561 22051 17595
rect 22201 17561 22235 17595
rect 7205 17493 7239 17527
rect 8309 17493 8343 17527
rect 9137 17493 9171 17527
rect 13461 17493 13495 17527
rect 15485 17493 15519 17527
rect 17417 17493 17451 17527
rect 17877 17493 17911 17527
rect 18705 17493 18739 17527
rect 19441 17493 19475 17527
rect 19809 17493 19843 17527
rect 21281 17493 21315 17527
rect 24593 17493 24627 17527
rect 24961 17493 24995 17527
rect 8033 17289 8067 17323
rect 9045 17289 9079 17323
rect 9413 17289 9447 17323
rect 17509 17289 17543 17323
rect 20361 17289 20395 17323
rect 22017 17289 22051 17323
rect 22753 17289 22787 17323
rect 10977 17221 11011 17255
rect 13185 17221 13219 17255
rect 16957 17221 16991 17255
rect 17969 17221 18003 17255
rect 20729 17221 20763 17255
rect 23765 17221 23799 17255
rect 10241 17153 10275 17187
rect 14565 17153 14599 17187
rect 21281 17153 21315 17187
rect 22661 17153 22695 17187
rect 23489 17153 23523 17187
rect 8125 17085 8159 17119
rect 8309 17085 8343 17119
rect 8769 17085 8803 17119
rect 9505 17085 9539 17119
rect 9597 17085 9631 17119
rect 11897 17085 11931 17119
rect 12541 17085 12575 17119
rect 13277 17085 13311 17119
rect 13461 17085 13495 17119
rect 14841 17085 14875 17119
rect 16313 17085 16347 17119
rect 18613 17085 18647 17119
rect 18889 17085 18923 17119
rect 22845 17085 22879 17119
rect 25237 17085 25271 17119
rect 7665 17017 7699 17051
rect 12817 17017 12851 17051
rect 18153 17017 18187 17051
rect 22293 17017 22327 17051
rect 7297 16949 7331 16983
rect 11529 16949 11563 16983
rect 12081 16949 12115 16983
rect 17049 16949 17083 16983
rect 8585 16745 8619 16779
rect 11345 16745 11379 16779
rect 13921 16745 13955 16779
rect 22293 16745 22327 16779
rect 16865 16677 16899 16711
rect 10701 16609 10735 16643
rect 10885 16609 10919 16643
rect 11805 16609 11839 16643
rect 15117 16609 15151 16643
rect 16313 16609 16347 16643
rect 17969 16609 18003 16643
rect 20269 16609 20303 16643
rect 16129 16541 16163 16575
rect 18889 16541 18923 16575
rect 19809 16541 19843 16575
rect 22661 16541 22695 16575
rect 23581 16541 23615 16575
rect 24777 16541 24811 16575
rect 10609 16473 10643 16507
rect 12081 16473 12115 16507
rect 14933 16473 14967 16507
rect 17233 16473 17267 16507
rect 20545 16473 20579 16507
rect 25421 16473 25455 16507
rect 9873 16405 9907 16439
rect 10241 16405 10275 16439
rect 13553 16405 13587 16439
rect 14289 16405 14323 16439
rect 14565 16405 14599 16439
rect 15025 16405 15059 16439
rect 15761 16405 15795 16439
rect 16221 16405 16255 16439
rect 18705 16405 18739 16439
rect 19257 16405 19291 16439
rect 19625 16405 19659 16439
rect 22017 16405 22051 16439
rect 24593 16405 24627 16439
rect 8309 16201 8343 16235
rect 13369 16201 13403 16235
rect 14565 16201 14599 16235
rect 15761 16201 15795 16235
rect 16221 16201 16255 16235
rect 16865 16201 16899 16235
rect 8585 16133 8619 16167
rect 11805 16133 11839 16167
rect 13829 16133 13863 16167
rect 17233 16133 17267 16167
rect 20085 16133 20119 16167
rect 6561 16065 6595 16099
rect 12541 16065 12575 16099
rect 12633 16065 12667 16099
rect 13737 16065 13771 16099
rect 14933 16065 14967 16099
rect 18061 16065 18095 16099
rect 18705 16065 18739 16099
rect 19257 16065 19291 16099
rect 21097 16065 21131 16099
rect 22017 16065 22051 16099
rect 24777 16065 24811 16099
rect 6837 15997 6871 16031
rect 12725 15997 12759 16031
rect 14013 15997 14047 16031
rect 15025 15997 15059 16031
rect 15117 15997 15151 16031
rect 21189 15997 21223 16031
rect 21373 15997 21407 16031
rect 22293 15997 22327 16031
rect 24501 15997 24535 16031
rect 12173 15929 12207 15963
rect 17325 15861 17359 15895
rect 17877 15861 17911 15895
rect 18521 15861 18555 15895
rect 20729 15861 20763 15895
rect 23765 15861 23799 15895
rect 24133 15861 24167 15895
rect 9137 15657 9171 15691
rect 11621 15657 11655 15691
rect 15485 15657 15519 15691
rect 18521 15657 18555 15691
rect 21189 15657 21223 15691
rect 13185 15589 13219 15623
rect 9689 15521 9723 15555
rect 12265 15521 12299 15555
rect 12633 15521 12667 15555
rect 16405 15521 16439 15555
rect 16681 15521 16715 15555
rect 19441 15521 19475 15555
rect 22293 15521 22327 15555
rect 22569 15521 22603 15555
rect 24041 15521 24075 15555
rect 24593 15521 24627 15555
rect 10149 15453 10183 15487
rect 12081 15453 12115 15487
rect 21833 15453 21867 15487
rect 9597 15385 9631 15419
rect 11989 15385 12023 15419
rect 19717 15385 19751 15419
rect 9505 15317 9539 15351
rect 14289 15317 14323 15351
rect 14749 15317 14783 15351
rect 15761 15317 15795 15351
rect 18153 15317 18187 15351
rect 21649 15317 21683 15351
rect 25053 15317 25087 15351
rect 10149 15113 10183 15147
rect 13737 15113 13771 15147
rect 14105 15113 14139 15147
rect 15945 15113 15979 15147
rect 17509 15113 17543 15147
rect 20085 15113 20119 15147
rect 10517 15045 10551 15079
rect 18705 15045 18739 15079
rect 23305 15045 23339 15079
rect 25145 15045 25179 15079
rect 19993 14977 20027 15011
rect 21005 14977 21039 15011
rect 21373 14977 21407 15011
rect 22109 14977 22143 15011
rect 24133 14977 24167 15011
rect 7665 14909 7699 14943
rect 7941 14909 7975 14943
rect 9689 14909 9723 14943
rect 10609 14909 10643 14943
rect 10701 14909 10735 14943
rect 13461 14909 13495 14943
rect 14197 14909 14231 14943
rect 14381 14909 14415 14943
rect 16037 14909 16071 14943
rect 16221 14909 16255 14943
rect 20269 14909 20303 14943
rect 12173 14841 12207 14875
rect 15577 14841 15611 14875
rect 19625 14841 19659 14875
rect 20821 14841 20855 14875
rect 11345 14773 11379 14807
rect 12541 14773 12575 14807
rect 15301 14773 15335 14807
rect 18797 14773 18831 14807
rect 8217 14569 8251 14603
rect 8585 14569 8619 14603
rect 12449 14569 12483 14603
rect 15393 14569 15427 14603
rect 21465 14569 21499 14603
rect 9597 14501 9631 14535
rect 6469 14433 6503 14467
rect 10241 14433 10275 14467
rect 11989 14433 12023 14467
rect 13001 14433 13035 14467
rect 14933 14433 14967 14467
rect 16957 14433 16991 14467
rect 17141 14433 17175 14467
rect 21925 14433 21959 14467
rect 22109 14433 22143 14467
rect 23857 14433 23891 14467
rect 9965 14365 9999 14399
rect 13461 14365 13495 14399
rect 20453 14365 20487 14399
rect 22845 14365 22879 14399
rect 25053 14365 25087 14399
rect 6745 14297 6779 14331
rect 12909 14297 12943 14331
rect 14749 14297 14783 14331
rect 16865 14297 16899 14331
rect 17693 14297 17727 14331
rect 12817 14229 12851 14263
rect 13921 14229 13955 14263
rect 14289 14229 14323 14263
rect 14657 14229 14691 14263
rect 16497 14229 16531 14263
rect 20269 14229 20303 14263
rect 21833 14229 21867 14263
rect 24869 14229 24903 14263
rect 12265 14025 12299 14059
rect 13001 14025 13035 14059
rect 15577 14025 15611 14059
rect 8033 13957 8067 13991
rect 10241 13957 10275 13991
rect 19165 13957 19199 13991
rect 19533 13957 19567 13991
rect 19717 13957 19751 13991
rect 7757 13889 7791 13923
rect 10977 13889 11011 13923
rect 18981 13889 19015 13923
rect 20361 13889 20395 13923
rect 21097 13889 21131 13923
rect 22201 13889 22235 13923
rect 25237 13889 25271 13923
rect 9781 13821 9815 13855
rect 11713 13821 11747 13855
rect 13093 13821 13127 13855
rect 13185 13821 13219 13855
rect 13829 13821 13863 13855
rect 15945 13821 15979 13855
rect 16865 13821 16899 13855
rect 17141 13821 17175 13855
rect 18613 13821 18647 13855
rect 22845 13821 22879 13855
rect 23121 13821 23155 13855
rect 24593 13821 24627 13855
rect 20177 13753 20211 13787
rect 22017 13753 22051 13787
rect 12633 13685 12667 13719
rect 14092 13685 14126 13719
rect 20913 13685 20947 13719
rect 25053 13685 25087 13719
rect 8309 13481 8343 13515
rect 8677 13481 8711 13515
rect 9229 13481 9263 13515
rect 10688 13481 10722 13515
rect 21097 13481 21131 13515
rect 24593 13481 24627 13515
rect 6561 13345 6595 13379
rect 6837 13345 6871 13379
rect 9781 13345 9815 13379
rect 10425 13345 10459 13379
rect 13461 13345 13495 13379
rect 15761 13345 15795 13379
rect 16313 13345 16347 13379
rect 20269 13345 20303 13379
rect 23765 13345 23799 13379
rect 12633 13277 12667 13311
rect 14933 13277 14967 13311
rect 15669 13277 15703 13311
rect 17509 13277 17543 13311
rect 17877 13277 17911 13311
rect 18613 13277 18647 13311
rect 19441 13277 19475 13311
rect 20821 13277 20855 13311
rect 21373 13277 21407 13311
rect 21649 13277 21683 13311
rect 22753 13277 22787 13311
rect 24777 13277 24811 13311
rect 9597 13209 9631 13243
rect 15577 13209 15611 13243
rect 18061 13209 18095 13243
rect 18797 13209 18831 13243
rect 20729 13209 20763 13243
rect 9689 13141 9723 13175
rect 12173 13141 12207 13175
rect 13921 13141 13955 13175
rect 14657 13141 14691 13175
rect 15209 13141 15243 13175
rect 25053 13141 25087 13175
rect 7849 12937 7883 12971
rect 9045 12937 9079 12971
rect 9413 12937 9447 12971
rect 10425 12937 10459 12971
rect 10793 12937 10827 12971
rect 11621 12937 11655 12971
rect 11897 12937 11931 12971
rect 12081 12937 12115 12971
rect 12265 12937 12299 12971
rect 17325 12937 17359 12971
rect 18061 12937 18095 12971
rect 18797 12937 18831 12971
rect 22477 12937 22511 12971
rect 25145 12937 25179 12971
rect 9505 12869 9539 12903
rect 13093 12869 13127 12903
rect 14197 12869 14231 12903
rect 21189 12869 21223 12903
rect 23397 12869 23431 12903
rect 7021 12801 7055 12835
rect 7113 12801 7147 12835
rect 8217 12801 8251 12835
rect 10885 12801 10919 12835
rect 13001 12801 13035 12835
rect 14289 12801 14323 12835
rect 15393 12801 15427 12835
rect 15485 12801 15519 12835
rect 17233 12801 17267 12835
rect 18245 12801 18279 12835
rect 19165 12801 19199 12835
rect 20177 12801 20211 12835
rect 21097 12801 21131 12835
rect 22201 12801 22235 12835
rect 23121 12801 23155 12835
rect 7205 12733 7239 12767
rect 8309 12733 8343 12767
rect 8493 12733 8527 12767
rect 9689 12733 9723 12767
rect 10977 12733 11011 12767
rect 13185 12733 13219 12767
rect 14381 12733 14415 12767
rect 15577 12733 15611 12767
rect 17509 12733 17543 12767
rect 19257 12733 19291 12767
rect 19441 12733 19475 12767
rect 21373 12733 21407 12767
rect 6653 12665 6687 12699
rect 16865 12665 16899 12699
rect 22017 12665 22051 12699
rect 11713 12597 11747 12631
rect 12633 12597 12667 12631
rect 13829 12597 13863 12631
rect 15025 12597 15059 12631
rect 16129 12597 16163 12631
rect 19993 12597 20027 12631
rect 20729 12597 20763 12631
rect 22661 12597 22695 12631
rect 24869 12597 24903 12631
rect 10241 12393 10275 12427
rect 11437 12393 11471 12427
rect 12633 12393 12667 12427
rect 16313 12393 16347 12427
rect 22201 12393 22235 12427
rect 24593 12393 24627 12427
rect 14289 12325 14323 12359
rect 15301 12325 15335 12359
rect 7389 12257 7423 12291
rect 8217 12257 8251 12291
rect 10793 12257 10827 12291
rect 11989 12257 12023 12291
rect 13277 12257 13311 12291
rect 14841 12257 14875 12291
rect 15577 12257 15611 12291
rect 18705 12257 18739 12291
rect 19993 12257 20027 12291
rect 20453 12257 20487 12291
rect 20729 12257 20763 12291
rect 11805 12189 11839 12223
rect 13093 12189 13127 12223
rect 13645 12189 13679 12223
rect 13921 12189 13955 12223
rect 14749 12189 14783 12223
rect 17325 12189 17359 12223
rect 19533 12189 19567 12223
rect 22845 12189 22879 12223
rect 24777 12189 24811 12223
rect 10701 12121 10735 12155
rect 18061 12121 18095 12155
rect 23857 12121 23891 12155
rect 8953 12053 8987 12087
rect 10609 12053 10643 12087
rect 11897 12053 11931 12087
rect 13001 12053 13035 12087
rect 14657 12053 14691 12087
rect 15669 12053 15703 12087
rect 16681 12053 16715 12087
rect 19625 12053 19659 12087
rect 9045 11849 9079 11883
rect 9873 11849 9907 11883
rect 10241 11849 10275 11883
rect 11897 11849 11931 11883
rect 13093 11849 13127 11883
rect 13461 11849 13495 11883
rect 13553 11849 13587 11883
rect 14289 11849 14323 11883
rect 14749 11849 14783 11883
rect 17325 11849 17359 11883
rect 18061 11849 18095 11883
rect 18429 11849 18463 11883
rect 21189 11849 21223 11883
rect 9597 11781 9631 11815
rect 10333 11781 10367 11815
rect 21373 11781 21407 11815
rect 23305 11781 23339 11815
rect 11253 11713 11287 11747
rect 11621 11713 11655 11747
rect 12265 11713 12299 11747
rect 14657 11713 14691 11747
rect 15393 11713 15427 11747
rect 15577 11713 15611 11747
rect 17233 11713 17267 11747
rect 19349 11713 19383 11747
rect 20085 11713 20119 11747
rect 22293 11713 22327 11747
rect 24133 11713 24167 11747
rect 7297 11645 7331 11679
rect 7573 11645 7607 11679
rect 10425 11645 10459 11679
rect 12357 11645 12391 11679
rect 12449 11645 12483 11679
rect 13737 11645 13771 11679
rect 14841 11645 14875 11679
rect 17417 11645 17451 11679
rect 18521 11645 18555 11679
rect 18705 11645 18739 11679
rect 20729 11645 20763 11679
rect 21649 11645 21683 11679
rect 24777 11645 24811 11679
rect 16865 11577 16899 11611
rect 9413 11509 9447 11543
rect 19441 11509 19475 11543
rect 20177 11509 20211 11543
rect 12633 11305 12667 11339
rect 17233 11305 17267 11339
rect 22109 11305 22143 11339
rect 25053 11305 25087 11339
rect 11437 11237 11471 11271
rect 16681 11237 16715 11271
rect 17877 11237 17911 11271
rect 18153 11237 18187 11271
rect 21557 11237 21591 11271
rect 9413 11169 9447 11203
rect 12081 11169 12115 11203
rect 13277 11169 13311 11203
rect 14933 11169 14967 11203
rect 18613 11169 18647 11203
rect 18797 11169 18831 11203
rect 20269 11169 20303 11203
rect 23305 11169 23339 11203
rect 9137 11101 9171 11135
rect 13001 11101 13035 11135
rect 13645 11101 13679 11135
rect 17049 11101 17083 11135
rect 19257 11101 19291 11135
rect 19993 11101 20027 11135
rect 20913 11101 20947 11135
rect 21741 11101 21775 11135
rect 22845 11101 22879 11135
rect 25237 11101 25271 11135
rect 13093 11033 13127 11067
rect 13921 11033 13955 11067
rect 15209 11033 15243 11067
rect 17601 11033 17635 11067
rect 18521 11033 18555 11067
rect 21097 11033 21131 11067
rect 10885 10965 10919 10999
rect 11805 10965 11839 10999
rect 11897 10965 11931 10999
rect 14289 10965 14323 10999
rect 19625 10965 19659 10999
rect 20085 10965 20119 10999
rect 9965 10761 9999 10795
rect 12357 10761 12391 10795
rect 12725 10761 12759 10795
rect 14197 10761 14231 10795
rect 15945 10761 15979 10795
rect 19901 10761 19935 10795
rect 20729 10761 20763 10795
rect 8493 10693 8527 10727
rect 17601 10693 17635 10727
rect 22477 10693 22511 10727
rect 23397 10693 23431 10727
rect 12817 10625 12851 10659
rect 17049 10625 17083 10659
rect 18429 10625 18463 10659
rect 19073 10625 19107 10659
rect 19993 10625 20027 10659
rect 21097 10625 21131 10659
rect 22201 10625 22235 10659
rect 23121 10625 23155 10659
rect 8217 10557 8251 10591
rect 11713 10557 11747 10591
rect 12909 10557 12943 10591
rect 14289 10557 14323 10591
rect 14473 10557 14507 10591
rect 15301 10557 15335 10591
rect 16037 10557 16071 10591
rect 16221 10557 16255 10591
rect 20177 10557 20211 10591
rect 21189 10557 21223 10591
rect 21281 10557 21315 10591
rect 10425 10489 10459 10523
rect 11069 10489 11103 10523
rect 13829 10489 13863 10523
rect 15577 10489 15611 10523
rect 16865 10489 16899 10523
rect 18245 10489 18279 10523
rect 25145 10489 25179 10523
rect 7849 10421 7883 10455
rect 11253 10421 11287 10455
rect 13461 10421 13495 10455
rect 17693 10421 17727 10455
rect 18889 10421 18923 10455
rect 19533 10421 19567 10455
rect 22017 10421 22051 10455
rect 22661 10421 22695 10455
rect 24869 10421 24903 10455
rect 11069 10217 11103 10251
rect 11621 10217 11655 10251
rect 12817 10217 12851 10251
rect 14565 10217 14599 10251
rect 15669 10217 15703 10251
rect 22293 10217 22327 10251
rect 24593 10217 24627 10251
rect 17969 10149 18003 10183
rect 9597 10081 9631 10115
rect 12173 10081 12207 10115
rect 13461 10081 13495 10115
rect 13921 10081 13955 10115
rect 15025 10081 15059 10115
rect 15117 10081 15151 10115
rect 18613 10081 18647 10115
rect 23305 10081 23339 10115
rect 23397 10081 23431 10115
rect 9321 10013 9355 10047
rect 13185 10013 13219 10047
rect 14289 10013 14323 10047
rect 20545 10013 20579 10047
rect 24777 10013 24811 10047
rect 11989 9945 12023 9979
rect 14933 9945 14967 9979
rect 16865 9945 16899 9979
rect 19533 9945 19567 9979
rect 20821 9945 20855 9979
rect 12081 9877 12115 9911
rect 13277 9877 13311 9911
rect 15853 9877 15887 9911
rect 16037 9877 16071 9911
rect 16129 9877 16163 9911
rect 16957 9877 16991 9911
rect 18337 9877 18371 9911
rect 18429 9877 18463 9911
rect 18981 9877 19015 9911
rect 19625 9877 19659 9911
rect 19993 9877 20027 9911
rect 20177 9877 20211 9911
rect 22845 9877 22879 9911
rect 23213 9877 23247 9911
rect 11345 9673 11379 9707
rect 22017 9673 22051 9707
rect 15485 9605 15519 9639
rect 11713 9537 11747 9571
rect 14289 9537 14323 9571
rect 20269 9537 20303 9571
rect 22661 9537 22695 9571
rect 25053 9537 25087 9571
rect 14381 9469 14415 9503
rect 14565 9469 14599 9503
rect 15577 9469 15611 9503
rect 15761 9469 15795 9503
rect 17325 9469 17359 9503
rect 21189 9469 21223 9503
rect 22937 9469 22971 9503
rect 25329 9469 25363 9503
rect 13461 9401 13495 9435
rect 13921 9401 13955 9435
rect 16129 9401 16163 9435
rect 16405 9401 16439 9435
rect 11976 9333 12010 9367
rect 15117 9333 15151 9367
rect 16865 9333 16899 9367
rect 17049 9333 17083 9367
rect 17588 9333 17622 9367
rect 19073 9333 19107 9367
rect 19441 9333 19475 9367
rect 24409 9333 24443 9367
rect 24869 9333 24903 9367
rect 11161 9129 11195 9163
rect 12633 9129 12667 9163
rect 14289 9129 14323 9163
rect 18245 9129 18279 9163
rect 21373 9129 21407 9163
rect 13001 9061 13035 9095
rect 15485 9061 15519 9095
rect 9137 8993 9171 9027
rect 13553 8993 13587 9027
rect 14841 8993 14875 9027
rect 16497 8993 16531 9027
rect 17785 8993 17819 9027
rect 13461 8925 13495 8959
rect 16405 8925 16439 8959
rect 17601 8925 17635 8959
rect 19625 8925 19659 8959
rect 22017 8925 22051 8959
rect 22661 8925 22695 8959
rect 24777 8925 24811 8959
rect 9413 8857 9447 8891
rect 13369 8857 13403 8891
rect 17509 8857 17543 8891
rect 18705 8857 18739 8891
rect 18889 8857 18923 8891
rect 19901 8857 19935 8891
rect 23857 8857 23891 8891
rect 10885 8789 10919 8823
rect 14657 8789 14691 8823
rect 14749 8789 14783 8823
rect 15393 8789 15427 8823
rect 15945 8789 15979 8823
rect 16313 8789 16347 8823
rect 17141 8789 17175 8823
rect 21833 8789 21867 8823
rect 22385 8789 22419 8823
rect 24593 8789 24627 8823
rect 12817 8585 12851 8619
rect 14473 8585 14507 8619
rect 15071 8585 15105 8619
rect 13921 8517 13955 8551
rect 14105 8517 14139 8551
rect 14841 8449 14875 8483
rect 16129 8449 16163 8483
rect 17233 8449 17267 8483
rect 17325 8449 17359 8483
rect 17969 8449 18003 8483
rect 18429 8449 18463 8483
rect 20269 8449 20303 8483
rect 22201 8449 22235 8483
rect 23949 8449 23983 8483
rect 11713 8381 11747 8415
rect 13185 8381 13219 8415
rect 17417 8381 17451 8415
rect 19441 8381 19475 8415
rect 21281 8381 21315 8415
rect 22569 8381 22603 8415
rect 24777 8381 24811 8415
rect 16865 8313 16899 8347
rect 11069 8041 11103 8075
rect 13001 8041 13035 8075
rect 14289 8041 14323 8075
rect 15853 8041 15887 8075
rect 24869 7973 24903 8007
rect 11713 7905 11747 7939
rect 13645 7905 13679 7939
rect 14841 7905 14875 7939
rect 16405 7905 16439 7939
rect 18705 7905 18739 7939
rect 22385 7905 22419 7939
rect 11437 7837 11471 7871
rect 13369 7837 13403 7871
rect 14657 7837 14691 7871
rect 17693 7837 17727 7871
rect 20453 7837 20487 7871
rect 22109 7837 22143 7871
rect 11529 7769 11563 7803
rect 13461 7769 13495 7803
rect 14749 7769 14783 7803
rect 15393 7769 15427 7803
rect 16221 7769 16255 7803
rect 21465 7769 21499 7803
rect 24685 7769 24719 7803
rect 12357 7701 12391 7735
rect 16313 7701 16347 7735
rect 19441 7701 19475 7735
rect 19901 7701 19935 7735
rect 23857 7701 23891 7735
rect 24225 7701 24259 7735
rect 11989 7497 12023 7531
rect 12633 7497 12667 7531
rect 15485 7497 15519 7531
rect 17785 7497 17819 7531
rect 21189 7497 21223 7531
rect 11069 7429 11103 7463
rect 16129 7429 16163 7463
rect 16865 7429 16899 7463
rect 17693 7429 17727 7463
rect 20545 7429 20579 7463
rect 21097 7429 21131 7463
rect 25145 7429 25179 7463
rect 22293 7361 22327 7395
rect 23949 7361 23983 7395
rect 9045 7293 9079 7327
rect 9321 7293 9355 7327
rect 12725 7293 12759 7327
rect 12817 7293 12851 7327
rect 13737 7293 13771 7327
rect 14013 7293 14047 7327
rect 17877 7293 17911 7327
rect 18521 7293 18555 7327
rect 18797 7293 18831 7327
rect 21281 7293 21315 7327
rect 23305 7293 23339 7327
rect 10793 7225 10827 7259
rect 16313 7225 16347 7259
rect 12265 7157 12299 7191
rect 16681 7157 16715 7191
rect 17325 7157 17359 7191
rect 20269 7157 20303 7191
rect 20729 7157 20763 7191
rect 12541 6953 12575 6987
rect 20453 6953 20487 6987
rect 10793 6817 10827 6851
rect 14197 6817 14231 6851
rect 17417 6817 17451 6851
rect 18889 6817 18923 6851
rect 19901 6817 19935 6851
rect 20085 6817 20119 6851
rect 25053 6817 25087 6851
rect 25145 6817 25179 6851
rect 13737 6749 13771 6783
rect 15485 6749 15519 6783
rect 17141 6749 17175 6783
rect 20913 6749 20947 6783
rect 22661 6749 22695 6783
rect 11069 6681 11103 6715
rect 14657 6681 14691 6715
rect 16497 6681 16531 6715
rect 21833 6681 21867 6715
rect 23857 6681 23891 6715
rect 12817 6613 12851 6647
rect 13553 6613 13587 6647
rect 14749 6613 14783 6647
rect 19441 6613 19475 6647
rect 19809 6613 19843 6647
rect 24593 6613 24627 6647
rect 24961 6613 24995 6647
rect 10425 6409 10459 6443
rect 12173 6409 12207 6443
rect 12817 6409 12851 6443
rect 13369 6409 13403 6443
rect 17325 6409 17359 6443
rect 17969 6409 18003 6443
rect 24593 6409 24627 6443
rect 10885 6341 10919 6375
rect 10793 6273 10827 6307
rect 12081 6273 12115 6307
rect 13737 6273 13771 6307
rect 13829 6273 13863 6307
rect 14381 6273 14415 6307
rect 15117 6273 15151 6307
rect 17233 6273 17267 6307
rect 18245 6273 18279 6307
rect 20269 6273 20303 6307
rect 22017 6273 22051 6307
rect 24777 6273 24811 6307
rect 10977 6205 11011 6239
rect 12265 6205 12299 6239
rect 13921 6205 13955 6239
rect 16129 6205 16163 6239
rect 17417 6205 17451 6239
rect 19441 6205 19475 6239
rect 21281 6205 21315 6239
rect 22293 6205 22327 6239
rect 11713 6137 11747 6171
rect 16865 6137 16899 6171
rect 13001 6069 13035 6103
rect 23765 6069 23799 6103
rect 24041 6069 24075 6103
rect 24225 6069 24259 6103
rect 11805 5865 11839 5899
rect 13553 5865 13587 5899
rect 14197 5865 14231 5899
rect 14749 5865 14783 5899
rect 17693 5865 17727 5899
rect 23857 5865 23891 5899
rect 25237 5865 25271 5899
rect 18153 5797 18187 5831
rect 24869 5797 24903 5831
rect 10333 5729 10367 5763
rect 12265 5729 12299 5763
rect 14473 5729 14507 5763
rect 15209 5729 15243 5763
rect 15393 5729 15427 5763
rect 18613 5729 18647 5763
rect 18705 5729 18739 5763
rect 19901 5729 19935 5763
rect 21741 5729 21775 5763
rect 10057 5661 10091 5695
rect 12541 5661 12575 5695
rect 13737 5661 13771 5695
rect 15945 5661 15979 5695
rect 18521 5661 18555 5695
rect 19625 5661 19659 5695
rect 21465 5661 21499 5695
rect 23213 5661 23247 5695
rect 24041 5661 24075 5695
rect 24685 5661 24719 5695
rect 16221 5593 16255 5627
rect 23397 5593 23431 5627
rect 15117 5525 15151 5559
rect 25329 5525 25363 5559
rect 10977 5321 11011 5355
rect 14933 5321 14967 5355
rect 20545 5321 20579 5355
rect 11529 5253 11563 5287
rect 13461 5253 13495 5287
rect 17877 5253 17911 5287
rect 21557 5253 21591 5287
rect 10701 5185 10735 5219
rect 11161 5185 11195 5219
rect 13185 5185 13219 5219
rect 17141 5185 17175 5219
rect 18797 5185 18831 5219
rect 21097 5185 21131 5219
rect 22109 5185 22143 5219
rect 23857 5185 23891 5219
rect 11805 5117 11839 5151
rect 11897 5117 11931 5151
rect 12173 5117 12207 5151
rect 15485 5117 15519 5151
rect 15761 5117 15795 5151
rect 19073 5117 19107 5151
rect 22477 5117 22511 5151
rect 24317 5117 24351 5151
rect 21189 4981 21223 5015
rect 10149 4777 10183 4811
rect 21281 4777 21315 4811
rect 24777 4777 24811 4811
rect 10425 4709 10459 4743
rect 16865 4709 16899 4743
rect 25329 4709 25363 4743
rect 2053 4641 2087 4675
rect 5089 4641 5123 4675
rect 11345 4641 11379 4675
rect 15117 4641 15151 4675
rect 19533 4641 19567 4675
rect 1777 4573 1811 4607
rect 3985 4573 4019 4607
rect 7113 4573 7147 4607
rect 9873 4573 9907 4607
rect 10609 4573 10643 4607
rect 11069 4573 11103 4607
rect 12541 4573 12575 4607
rect 14473 4573 14507 4607
rect 17601 4573 17635 4607
rect 21833 4573 21867 4607
rect 23673 4573 23707 4607
rect 24133 4573 24167 4607
rect 4629 4505 4663 4539
rect 5365 4505 5399 4539
rect 7389 4505 7423 4539
rect 9781 4505 9815 4539
rect 13553 4505 13587 4539
rect 15393 4505 15427 4539
rect 18337 4505 18371 4539
rect 19809 4505 19843 4539
rect 22661 4505 22695 4539
rect 24685 4505 24719 4539
rect 25145 4505 25179 4539
rect 1593 4437 1627 4471
rect 14289 4437 14323 4471
rect 14749 4437 14783 4471
rect 23765 4437 23799 4471
rect 2237 4233 2271 4267
rect 15669 4233 15703 4267
rect 16129 4233 16163 4267
rect 21557 4233 21591 4267
rect 22017 4233 22051 4267
rect 24685 4233 24719 4267
rect 14197 4165 14231 4199
rect 22477 4165 22511 4199
rect 1593 4097 1627 4131
rect 2881 4097 2915 4131
rect 3157 4097 3191 4131
rect 4353 4097 4387 4131
rect 9505 4097 9539 4131
rect 10609 4097 10643 4131
rect 12265 4097 12299 4131
rect 13921 4097 13955 4131
rect 17049 4097 17083 4131
rect 18705 4097 18739 4131
rect 20913 4097 20947 4131
rect 21005 4097 21039 4131
rect 21833 4097 21867 4131
rect 25145 4097 25179 4131
rect 10333 4029 10367 4063
rect 11621 4029 11655 4063
rect 13277 4029 13311 4063
rect 17325 4029 17359 4063
rect 19165 4029 19199 4063
rect 21189 4029 21223 4063
rect 24133 4029 24167 4063
rect 2697 3961 2731 3995
rect 4169 3961 4203 3995
rect 9321 3961 9355 3995
rect 9873 3961 9907 3995
rect 3893 3893 3927 3927
rect 4813 3893 4847 3927
rect 6101 3893 6135 3927
rect 7021 3893 7055 3927
rect 9045 3893 9079 3927
rect 10057 3893 10091 3927
rect 11805 3893 11839 3927
rect 20545 3893 20579 3927
rect 25329 3893 25363 3927
rect 2881 3689 2915 3723
rect 4261 3689 4295 3723
rect 8401 3689 8435 3723
rect 10425 3689 10459 3723
rect 23857 3689 23891 3723
rect 6377 3621 6411 3655
rect 7113 3621 7147 3655
rect 9689 3621 9723 3655
rect 1869 3553 1903 3587
rect 5181 3553 5215 3587
rect 11069 3553 11103 3587
rect 12817 3553 12851 3587
rect 14749 3553 14783 3587
rect 16589 3553 16623 3587
rect 18061 3553 18095 3587
rect 19901 3553 19935 3587
rect 21741 3553 21775 3587
rect 23213 3553 23247 3587
rect 1593 3485 1627 3519
rect 3065 3485 3099 3519
rect 3525 3485 3559 3519
rect 4445 3485 4479 3519
rect 4905 3485 4939 3519
rect 6561 3485 6595 3519
rect 7297 3485 7331 3519
rect 8585 3485 8619 3519
rect 8953 3485 8987 3519
rect 9873 3485 9907 3519
rect 10609 3485 10643 3519
rect 11345 3485 11379 3519
rect 12449 3485 12483 3519
rect 14473 3485 14507 3519
rect 16313 3485 16347 3519
rect 18337 3485 18371 3519
rect 19441 3485 19475 3519
rect 21373 3485 21407 3519
rect 24041 3485 24075 3519
rect 24593 3485 24627 3519
rect 7849 3417 7883 3451
rect 3341 3349 3375 3383
rect 3801 3349 3835 3383
rect 6101 3349 6135 3383
rect 7757 3349 7791 3383
rect 9229 3349 9263 3383
rect 9413 3349 9447 3383
rect 25237 3349 25271 3383
rect 7205 3145 7239 3179
rect 9689 3145 9723 3179
rect 10333 3145 10367 3179
rect 10977 3145 11011 3179
rect 21281 3145 21315 3179
rect 22201 3145 22235 3179
rect 22937 3145 22971 3179
rect 23673 3145 23707 3179
rect 24225 3145 24259 3179
rect 9413 3077 9447 3111
rect 20637 3077 20671 3111
rect 20821 3077 20855 3111
rect 22109 3077 22143 3111
rect 22845 3077 22879 3111
rect 23581 3077 23615 3111
rect 25421 3077 25455 3111
rect 2421 3009 2455 3043
rect 3709 3009 3743 3043
rect 5457 3009 5491 3043
rect 6745 3009 6779 3043
rect 7389 3009 7423 3043
rect 9045 3009 9079 3043
rect 9873 3009 9907 3043
rect 10517 3009 10551 3043
rect 11161 3009 11195 3043
rect 11989 3009 12023 3043
rect 13185 3009 13219 3043
rect 14841 3009 14875 3043
rect 17049 3009 17083 3043
rect 18889 3009 18923 3043
rect 24409 3009 24443 3043
rect 25145 3009 25179 3043
rect 2145 2941 2179 2975
rect 3433 2941 3467 2975
rect 5181 2941 5215 2975
rect 7849 2941 7883 2975
rect 9229 2941 9263 2975
rect 11713 2941 11747 2975
rect 13645 2941 13679 2975
rect 15301 2941 15335 2975
rect 17325 2941 17359 2975
rect 19165 2941 19199 2975
rect 6561 2873 6595 2907
rect 24961 2873 24995 2907
rect 4537 2805 4571 2839
rect 4905 2805 4939 2839
rect 8079 2805 8113 2839
rect 8401 2601 8435 2635
rect 16129 2601 16163 2635
rect 18705 2601 18739 2635
rect 21281 2533 21315 2567
rect 2881 2465 2915 2499
rect 5457 2465 5491 2499
rect 6837 2465 6871 2499
rect 10977 2465 11011 2499
rect 14933 2465 14967 2499
rect 16405 2465 16439 2499
rect 17325 2465 17359 2499
rect 19901 2465 19935 2499
rect 22477 2465 22511 2499
rect 23857 2465 23891 2499
rect 2605 2397 2639 2431
rect 3985 2397 4019 2431
rect 4721 2397 4755 2431
rect 5181 2397 5215 2431
rect 6653 2397 6687 2431
rect 7297 2397 7331 2431
rect 7941 2397 7975 2431
rect 8585 2397 8619 2431
rect 9321 2397 9355 2431
rect 9873 2397 9907 2431
rect 11897 2397 11931 2431
rect 12449 2397 12483 2431
rect 14105 2397 14139 2431
rect 14473 2397 14507 2431
rect 16865 2397 16899 2431
rect 18889 2397 18923 2431
rect 19441 2397 19475 2431
rect 21465 2397 21499 2431
rect 22201 2397 22235 2431
rect 24593 2397 24627 2431
rect 4261 2329 4295 2363
rect 13277 2329 13311 2363
rect 3801 2261 3835 2295
rect 4537 2261 4571 2295
rect 6469 2261 6503 2295
rect 7113 2261 7147 2295
rect 7757 2261 7791 2295
rect 9137 2261 9171 2295
rect 11713 2261 11747 2295
rect 25237 2261 25271 2295
<< metal1 >>
rect 1104 54426 25852 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 25852 54426
rect 1104 54352 25852 54374
rect 13814 54272 13820 54324
rect 13872 54272 13878 54324
rect 16546 54284 18276 54312
rect 2225 54179 2283 54185
rect 2225 54145 2237 54179
rect 2271 54176 2283 54179
rect 4062 54176 4068 54188
rect 2271 54148 4068 54176
rect 2271 54145 2283 54148
rect 2225 54139 2283 54145
rect 4062 54136 4068 54148
rect 4120 54136 4126 54188
rect 4798 54136 4804 54188
rect 4856 54136 4862 54188
rect 7374 54136 7380 54188
rect 7432 54136 7438 54188
rect 9582 54136 9588 54188
rect 9640 54136 9646 54188
rect 11698 54136 11704 54188
rect 11756 54176 11762 54188
rect 12161 54179 12219 54185
rect 12161 54176 12173 54179
rect 11756 54148 12173 54176
rect 11756 54136 11762 54148
rect 12161 54145 12173 54148
rect 12207 54145 12219 54179
rect 13832 54176 13860 54272
rect 16546 54244 16574 54284
rect 14568 54216 16574 54244
rect 14461 54179 14519 54185
rect 14461 54176 14473 54179
rect 13832 54148 14473 54176
rect 12161 54139 12219 54145
rect 14461 54145 14473 54148
rect 14507 54145 14519 54179
rect 14461 54139 14519 54145
rect 2406 54068 2412 54120
rect 2464 54108 2470 54120
rect 2501 54111 2559 54117
rect 2501 54108 2513 54111
rect 2464 54080 2513 54108
rect 2464 54068 2470 54080
rect 2501 54077 2513 54080
rect 2547 54077 2559 54111
rect 2501 54071 2559 54077
rect 5166 54068 5172 54120
rect 5224 54068 5230 54120
rect 7834 54068 7840 54120
rect 7892 54068 7898 54120
rect 9306 54068 9312 54120
rect 9364 54108 9370 54120
rect 9861 54111 9919 54117
rect 9861 54108 9873 54111
rect 9364 54080 9873 54108
rect 9364 54068 9370 54080
rect 9861 54077 9873 54080
rect 9907 54077 9919 54111
rect 9861 54071 9919 54077
rect 12342 54068 12348 54120
rect 12400 54108 12406 54120
rect 12621 54111 12679 54117
rect 12621 54108 12633 54111
rect 12400 54080 12633 54108
rect 12400 54068 12406 54080
rect 12621 54077 12633 54080
rect 12667 54077 12679 54111
rect 14568 54108 14596 54216
rect 14826 54136 14832 54188
rect 14884 54176 14890 54188
rect 15105 54179 15163 54185
rect 15105 54176 15117 54179
rect 14884 54148 15117 54176
rect 14884 54136 14890 54148
rect 15105 54145 15117 54148
rect 15151 54176 15163 54179
rect 15381 54179 15439 54185
rect 15381 54176 15393 54179
rect 15151 54148 15393 54176
rect 15151 54145 15163 54148
rect 15105 54139 15163 54145
rect 15381 54145 15393 54148
rect 15427 54145 15439 54179
rect 15381 54139 15439 54145
rect 16574 54136 16580 54188
rect 16632 54176 16638 54188
rect 17037 54179 17095 54185
rect 17037 54176 17049 54179
rect 16632 54148 17049 54176
rect 16632 54136 16638 54148
rect 17037 54145 17049 54148
rect 17083 54176 17095 54179
rect 17313 54179 17371 54185
rect 17313 54176 17325 54179
rect 17083 54148 17325 54176
rect 17083 54145 17095 54148
rect 17037 54139 17095 54145
rect 17313 54145 17325 54148
rect 17359 54145 17371 54179
rect 17313 54139 17371 54145
rect 17586 54136 17592 54188
rect 17644 54176 17650 54188
rect 17865 54179 17923 54185
rect 17865 54176 17877 54179
rect 17644 54148 17877 54176
rect 17644 54136 17650 54148
rect 17865 54145 17877 54148
rect 17911 54176 17923 54179
rect 18141 54179 18199 54185
rect 18141 54176 18153 54179
rect 17911 54148 18153 54176
rect 17911 54145 17923 54148
rect 17865 54139 17923 54145
rect 18141 54145 18153 54148
rect 18187 54145 18199 54179
rect 18141 54139 18199 54145
rect 12621 54071 12679 54077
rect 12728 54080 14596 54108
rect 18248 54108 18276 54284
rect 18966 54272 18972 54324
rect 19024 54272 19030 54324
rect 18984 54176 19012 54272
rect 19429 54179 19487 54185
rect 19429 54176 19441 54179
rect 18984 54148 19441 54176
rect 19429 54145 19441 54148
rect 19475 54145 19487 54179
rect 19429 54139 19487 54145
rect 20714 54136 20720 54188
rect 20772 54176 20778 54188
rect 21269 54179 21327 54185
rect 21269 54176 21281 54179
rect 20772 54148 21281 54176
rect 20772 54136 20778 54148
rect 21269 54145 21281 54148
rect 21315 54145 21327 54179
rect 21269 54139 21327 54145
rect 21726 54136 21732 54188
rect 21784 54176 21790 54188
rect 22005 54179 22063 54185
rect 22005 54176 22017 54179
rect 21784 54148 22017 54176
rect 21784 54136 21790 54148
rect 22005 54145 22017 54148
rect 22051 54176 22063 54179
rect 22557 54179 22615 54185
rect 22557 54176 22569 54179
rect 22051 54148 22569 54176
rect 22051 54145 22063 54148
rect 22005 54139 22063 54145
rect 22557 54145 22569 54148
rect 22603 54145 22615 54179
rect 22557 54139 22615 54145
rect 23106 54136 23112 54188
rect 23164 54176 23170 54188
rect 23201 54179 23259 54185
rect 23201 54176 23213 54179
rect 23164 54148 23213 54176
rect 23164 54136 23170 54148
rect 23201 54145 23213 54148
rect 23247 54176 23259 54179
rect 23753 54179 23811 54185
rect 23753 54176 23765 54179
rect 23247 54148 23765 54176
rect 23247 54145 23259 54148
rect 23201 54139 23259 54145
rect 23753 54145 23765 54148
rect 23799 54145 23811 54179
rect 23753 54139 23811 54145
rect 24029 54179 24087 54185
rect 24029 54145 24041 54179
rect 24075 54176 24087 54179
rect 24673 54179 24731 54185
rect 24673 54176 24685 54179
rect 24075 54148 24685 54176
rect 24075 54145 24087 54148
rect 24029 54139 24087 54145
rect 24673 54145 24685 54148
rect 24719 54176 24731 54179
rect 25866 54176 25872 54188
rect 24719 54148 25872 54176
rect 24719 54145 24731 54148
rect 24673 54139 24731 54145
rect 25866 54136 25872 54148
rect 25924 54136 25930 54188
rect 19705 54111 19763 54117
rect 19705 54108 19717 54111
rect 18248 54080 19717 54108
rect 8570 54000 8576 54052
rect 8628 54040 8634 54052
rect 12728 54040 12756 54080
rect 19705 54077 19717 54080
rect 19751 54077 19763 54111
rect 19705 54071 19763 54077
rect 8628 54012 12756 54040
rect 8628 54000 8634 54012
rect 13906 54000 13912 54052
rect 13964 54040 13970 54052
rect 14921 54043 14979 54049
rect 14921 54040 14933 54043
rect 13964 54012 14933 54040
rect 13964 54000 13970 54012
rect 14921 54009 14933 54012
rect 14967 54009 14979 54043
rect 14921 54003 14979 54009
rect 15654 54000 15660 54052
rect 15712 54040 15718 54052
rect 17681 54043 17739 54049
rect 17681 54040 17693 54043
rect 15712 54012 17693 54040
rect 15712 54000 15718 54012
rect 17681 54009 17693 54012
rect 17727 54009 17739 54043
rect 17681 54003 17739 54009
rect 20162 54000 20168 54052
rect 20220 54040 20226 54052
rect 22189 54043 22247 54049
rect 22189 54040 22201 54043
rect 20220 54012 22201 54040
rect 20220 54000 20226 54012
rect 22189 54009 22201 54012
rect 22235 54009 22247 54043
rect 22189 54003 22247 54009
rect 12710 53932 12716 53984
rect 12768 53972 12774 53984
rect 14277 53975 14335 53981
rect 14277 53972 14289 53975
rect 12768 53944 14289 53972
rect 12768 53932 12774 53944
rect 14277 53941 14289 53944
rect 14323 53941 14335 53975
rect 14277 53935 14335 53941
rect 15562 53932 15568 53984
rect 15620 53972 15626 53984
rect 16853 53975 16911 53981
rect 16853 53972 16865 53975
rect 15620 53944 16865 53972
rect 15620 53932 15626 53944
rect 16853 53941 16865 53944
rect 16899 53941 16911 53975
rect 16853 53935 16911 53941
rect 16942 53932 16948 53984
rect 17000 53972 17006 53984
rect 20901 53975 20959 53981
rect 20901 53972 20913 53975
rect 17000 53944 20913 53972
rect 17000 53932 17006 53944
rect 20901 53941 20913 53944
rect 20947 53941 20959 53975
rect 20901 53935 20959 53941
rect 22094 53932 22100 53984
rect 22152 53972 22158 53984
rect 23385 53975 23443 53981
rect 23385 53972 23397 53975
rect 22152 53944 23397 53972
rect 22152 53932 22158 53944
rect 23385 53941 23397 53944
rect 23431 53941 23443 53975
rect 23385 53935 23443 53941
rect 24213 53975 24271 53981
rect 24213 53941 24225 53975
rect 24259 53972 24271 53975
rect 25038 53972 25044 53984
rect 24259 53944 25044 53972
rect 24259 53941 24271 53944
rect 24213 53935 24271 53941
rect 25038 53932 25044 53944
rect 25096 53932 25102 53984
rect 25314 53932 25320 53984
rect 25372 53932 25378 53984
rect 1104 53882 25852 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 25852 53882
rect 1104 53808 25852 53830
rect 24486 53728 24492 53780
rect 24544 53728 24550 53780
rect 24762 53728 24768 53780
rect 24820 53728 24826 53780
rect 10686 53660 10692 53712
rect 10744 53660 10750 53712
rect 1026 53592 1032 53644
rect 1084 53632 1090 53644
rect 2041 53635 2099 53641
rect 2041 53632 2053 53635
rect 1084 53604 2053 53632
rect 1084 53592 1090 53604
rect 2041 53601 2053 53604
rect 2087 53601 2099 53635
rect 2041 53595 2099 53601
rect 3786 53592 3792 53644
rect 3844 53632 3850 53644
rect 4433 53635 4491 53641
rect 4433 53632 4445 53635
rect 3844 53604 4445 53632
rect 3844 53592 3850 53604
rect 4433 53601 4445 53604
rect 4479 53601 4491 53635
rect 4433 53595 4491 53601
rect 6546 53592 6552 53644
rect 6604 53632 6610 53644
rect 7101 53635 7159 53641
rect 7101 53632 7113 53635
rect 6604 53604 7113 53632
rect 6604 53592 6610 53604
rect 7101 53601 7113 53604
rect 7147 53601 7159 53635
rect 10704 53632 10732 53660
rect 11241 53635 11299 53641
rect 11241 53632 11253 53635
rect 10704 53604 11253 53632
rect 7101 53595 7159 53601
rect 11241 53601 11253 53604
rect 11287 53601 11299 53635
rect 11241 53595 11299 53601
rect 1765 53567 1823 53573
rect 1765 53533 1777 53567
rect 1811 53533 1823 53567
rect 1765 53527 1823 53533
rect 1780 53496 1808 53527
rect 4154 53524 4160 53576
rect 4212 53524 4218 53576
rect 6825 53567 6883 53573
rect 6825 53533 6837 53567
rect 6871 53564 6883 53567
rect 7834 53564 7840 53576
rect 6871 53536 7840 53564
rect 6871 53533 6883 53536
rect 6825 53527 6883 53533
rect 7834 53524 7840 53536
rect 7892 53524 7898 53576
rect 10686 53524 10692 53576
rect 10744 53564 10750 53576
rect 10781 53567 10839 53573
rect 10781 53564 10793 53567
rect 10744 53536 10793 53564
rect 10744 53524 10750 53536
rect 10781 53533 10793 53536
rect 10827 53533 10839 53567
rect 10781 53527 10839 53533
rect 22741 53567 22799 53573
rect 22741 53533 22753 53567
rect 22787 53564 22799 53567
rect 23109 53567 23167 53573
rect 23109 53564 23121 53567
rect 22787 53536 23121 53564
rect 22787 53533 22799 53536
rect 22741 53527 22799 53533
rect 23109 53533 23121 53536
rect 23155 53564 23167 53567
rect 23382 53564 23388 53576
rect 23155 53536 23388 53564
rect 23155 53533 23167 53536
rect 23109 53527 23167 53533
rect 23382 53524 23388 53536
rect 23440 53524 23446 53576
rect 23753 53567 23811 53573
rect 23753 53533 23765 53567
rect 23799 53564 23811 53567
rect 24486 53564 24492 53576
rect 23799 53536 24492 53564
rect 23799 53533 23811 53536
rect 23753 53527 23811 53533
rect 24486 53524 24492 53536
rect 24544 53524 24550 53576
rect 25038 53524 25044 53576
rect 25096 53524 25102 53576
rect 5534 53496 5540 53508
rect 1780 53468 5540 53496
rect 5534 53456 5540 53468
rect 5592 53456 5598 53508
rect 22830 53388 22836 53440
rect 22888 53428 22894 53440
rect 23201 53431 23259 53437
rect 23201 53428 23213 53431
rect 22888 53400 23213 53428
rect 22888 53388 22894 53400
rect 23201 53397 23213 53400
rect 23247 53397 23259 53431
rect 23201 53391 23259 53397
rect 23934 53388 23940 53440
rect 23992 53388 23998 53440
rect 25225 53431 25283 53437
rect 25225 53397 25237 53431
rect 25271 53428 25283 53431
rect 25866 53428 25872 53440
rect 25271 53400 25872 53428
rect 25271 53397 25283 53400
rect 25225 53391 25283 53397
rect 25866 53388 25872 53400
rect 25924 53388 25930 53440
rect 1104 53338 25852 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 25852 53338
rect 1104 53264 25852 53286
rect 4062 53184 4068 53236
rect 4120 53224 4126 53236
rect 5169 53227 5227 53233
rect 5169 53224 5181 53227
rect 4120 53196 5181 53224
rect 4120 53184 4126 53196
rect 5169 53193 5181 53196
rect 5215 53193 5227 53227
rect 5169 53187 5227 53193
rect 5353 53091 5411 53097
rect 5353 53057 5365 53091
rect 5399 53088 5411 53091
rect 7742 53088 7748 53100
rect 5399 53060 7748 53088
rect 5399 53057 5411 53060
rect 5353 53051 5411 53057
rect 7742 53048 7748 53060
rect 7800 53048 7806 53100
rect 23569 53091 23627 53097
rect 23569 53057 23581 53091
rect 23615 53057 23627 53091
rect 23569 53051 23627 53057
rect 24305 53091 24363 53097
rect 24305 53057 24317 53091
rect 24351 53088 24363 53091
rect 24762 53088 24768 53100
rect 24351 53060 24768 53088
rect 24351 53057 24363 53060
rect 24305 53051 24363 53057
rect 23584 53020 23612 53051
rect 24762 53048 24768 53060
rect 24820 53048 24826 53100
rect 25038 53048 25044 53100
rect 25096 53048 25102 53100
rect 24394 53020 24400 53032
rect 23584 52992 24400 53020
rect 24394 52980 24400 52992
rect 24452 52980 24458 53032
rect 18690 52912 18696 52964
rect 18748 52952 18754 52964
rect 25225 52955 25283 52961
rect 25225 52952 25237 52955
rect 18748 52924 25237 52952
rect 18748 52912 18754 52924
rect 25225 52921 25237 52924
rect 25271 52921 25283 52955
rect 25225 52915 25283 52921
rect 23750 52844 23756 52896
rect 23808 52844 23814 52896
rect 24486 52844 24492 52896
rect 24544 52844 24550 52896
rect 1104 52794 25852 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 25852 52794
rect 1104 52720 25852 52742
rect 4154 52640 4160 52692
rect 4212 52680 4218 52692
rect 6549 52683 6607 52689
rect 6549 52680 6561 52683
rect 4212 52652 6561 52680
rect 4212 52640 4218 52652
rect 6549 52649 6561 52652
rect 6595 52649 6607 52683
rect 6549 52643 6607 52649
rect 24029 52683 24087 52689
rect 24029 52649 24041 52683
rect 24075 52680 24087 52683
rect 24394 52680 24400 52692
rect 24075 52652 24400 52680
rect 24075 52649 24087 52652
rect 24029 52643 24087 52649
rect 24394 52640 24400 52652
rect 24452 52640 24458 52692
rect 6733 52479 6791 52485
rect 6733 52445 6745 52479
rect 6779 52476 6791 52479
rect 9490 52476 9496 52488
rect 6779 52448 9496 52476
rect 6779 52445 6791 52448
rect 6733 52439 6791 52445
rect 9490 52436 9496 52448
rect 9548 52436 9554 52488
rect 24581 52479 24639 52485
rect 24581 52445 24593 52479
rect 24627 52476 24639 52479
rect 25317 52479 25375 52485
rect 24627 52448 24992 52476
rect 24627 52445 24639 52448
rect 24581 52439 24639 52445
rect 24964 52420 24992 52448
rect 25317 52445 25329 52479
rect 25363 52476 25375 52479
rect 26510 52476 26516 52488
rect 25363 52448 26516 52476
rect 25363 52445 25375 52448
rect 25317 52439 25375 52445
rect 26510 52436 26516 52448
rect 26568 52436 26574 52488
rect 24946 52368 24952 52420
rect 25004 52368 25010 52420
rect 1104 52250 25852 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 25852 52250
rect 1104 52176 25852 52198
rect 24857 52139 24915 52145
rect 24857 52105 24869 52139
rect 24903 52136 24915 52139
rect 25038 52136 25044 52148
rect 24903 52108 25044 52136
rect 24903 52105 24915 52108
rect 24857 52099 24915 52105
rect 25038 52096 25044 52108
rect 25096 52096 25102 52148
rect 25314 51960 25320 52012
rect 25372 51960 25378 52012
rect 23382 51756 23388 51808
rect 23440 51796 23446 51808
rect 25133 51799 25191 51805
rect 25133 51796 25145 51799
rect 23440 51768 25145 51796
rect 23440 51756 23446 51768
rect 25133 51765 25145 51768
rect 25179 51765 25191 51799
rect 25133 51759 25191 51765
rect 1104 51706 25852 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 25852 51706
rect 1104 51632 25852 51654
rect 7374 51552 7380 51604
rect 7432 51592 7438 51604
rect 8297 51595 8355 51601
rect 8297 51592 8309 51595
rect 7432 51564 8309 51592
rect 7432 51552 7438 51564
rect 8297 51561 8309 51564
rect 8343 51561 8355 51595
rect 8297 51555 8355 51561
rect 7834 51484 7840 51536
rect 7892 51524 7898 51536
rect 9217 51527 9275 51533
rect 9217 51524 9229 51527
rect 7892 51496 9229 51524
rect 7892 51484 7898 51496
rect 9217 51493 9229 51496
rect 9263 51493 9275 51527
rect 9217 51487 9275 51493
rect 4798 51348 4804 51400
rect 4856 51388 4862 51400
rect 7837 51391 7895 51397
rect 7837 51388 7849 51391
rect 4856 51360 7849 51388
rect 4856 51348 4862 51360
rect 7837 51357 7849 51360
rect 7883 51357 7895 51391
rect 7837 51351 7895 51357
rect 8478 51348 8484 51400
rect 8536 51348 8542 51400
rect 9401 51391 9459 51397
rect 9401 51357 9413 51391
rect 9447 51388 9459 51391
rect 10502 51388 10508 51400
rect 9447 51360 10508 51388
rect 9447 51357 9459 51360
rect 9401 51351 9459 51357
rect 10502 51348 10508 51360
rect 10560 51348 10566 51400
rect 7653 51323 7711 51329
rect 7653 51289 7665 51323
rect 7699 51320 7711 51323
rect 10778 51320 10784 51332
rect 7699 51292 10784 51320
rect 7699 51289 7711 51292
rect 7653 51283 7711 51289
rect 10778 51280 10784 51292
rect 10836 51280 10842 51332
rect 24581 51323 24639 51329
rect 24581 51289 24593 51323
rect 24627 51320 24639 51323
rect 24946 51320 24952 51332
rect 24627 51292 24952 51320
rect 24627 51289 24639 51292
rect 24581 51283 24639 51289
rect 24946 51280 24952 51292
rect 25004 51280 25010 51332
rect 25317 51323 25375 51329
rect 25317 51289 25329 51323
rect 25363 51320 25375 51323
rect 26602 51320 26608 51332
rect 25363 51292 26608 51320
rect 25363 51289 25375 51292
rect 25317 51283 25375 51289
rect 26602 51280 26608 51292
rect 26660 51280 26666 51332
rect 1104 51162 25852 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 25852 51162
rect 1104 51088 25852 51110
rect 24581 50915 24639 50921
rect 24581 50881 24593 50915
rect 24627 50912 24639 50915
rect 24946 50912 24952 50924
rect 24627 50884 24952 50912
rect 24627 50881 24639 50884
rect 24581 50875 24639 50881
rect 24946 50872 24952 50884
rect 25004 50872 25010 50924
rect 18598 50668 18604 50720
rect 18656 50708 18662 50720
rect 25041 50711 25099 50717
rect 25041 50708 25053 50711
rect 18656 50680 25053 50708
rect 18656 50668 18662 50680
rect 25041 50677 25053 50680
rect 25087 50677 25099 50711
rect 25041 50671 25099 50677
rect 1104 50618 25852 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 25852 50618
rect 1104 50544 25852 50566
rect 5534 50464 5540 50516
rect 5592 50504 5598 50516
rect 7837 50507 7895 50513
rect 7837 50504 7849 50507
rect 5592 50476 7849 50504
rect 5592 50464 5598 50476
rect 7837 50473 7849 50476
rect 7883 50504 7895 50507
rect 8386 50504 8392 50516
rect 7883 50476 8392 50504
rect 7883 50473 7895 50476
rect 7837 50467 7895 50473
rect 8386 50464 8392 50476
rect 8444 50464 8450 50516
rect 9582 50464 9588 50516
rect 9640 50464 9646 50516
rect 7742 50396 7748 50448
rect 7800 50436 7806 50448
rect 8021 50439 8079 50445
rect 8021 50436 8033 50439
rect 7800 50408 8033 50436
rect 7800 50396 7806 50408
rect 8021 50405 8033 50408
rect 8067 50405 8079 50439
rect 8021 50399 8079 50405
rect 8389 50371 8447 50377
rect 8389 50368 8401 50371
rect 7576 50340 8401 50368
rect 7576 50309 7604 50340
rect 8389 50337 8401 50340
rect 8435 50368 8447 50371
rect 8570 50368 8576 50380
rect 8435 50340 8576 50368
rect 8435 50337 8447 50340
rect 8389 50331 8447 50337
rect 8570 50328 8576 50340
rect 8628 50328 8634 50380
rect 7561 50303 7619 50309
rect 7561 50269 7573 50303
rect 7607 50269 7619 50303
rect 7561 50263 7619 50269
rect 9493 50235 9551 50241
rect 9493 50201 9505 50235
rect 9539 50232 9551 50235
rect 9582 50232 9588 50244
rect 9539 50204 9588 50232
rect 9539 50201 9551 50204
rect 9493 50195 9551 50201
rect 9582 50192 9588 50204
rect 9640 50192 9646 50244
rect 25498 50124 25504 50176
rect 25556 50124 25562 50176
rect 1104 50074 25852 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 25852 50074
rect 1104 50000 25852 50022
rect 24489 49827 24547 49833
rect 24489 49793 24501 49827
rect 24535 49824 24547 49827
rect 25498 49824 25504 49836
rect 24535 49796 25504 49824
rect 24535 49793 24547 49796
rect 24489 49787 24547 49793
rect 25498 49784 25504 49796
rect 25556 49784 25562 49836
rect 24670 49716 24676 49768
rect 24728 49756 24734 49768
rect 24765 49759 24823 49765
rect 24765 49756 24777 49759
rect 24728 49728 24777 49756
rect 24728 49716 24734 49728
rect 24765 49725 24777 49728
rect 24811 49725 24823 49759
rect 24765 49719 24823 49725
rect 1104 49530 25852 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 25852 49530
rect 1104 49456 25852 49478
rect 10686 49308 10692 49360
rect 10744 49308 10750 49360
rect 11698 49308 11704 49360
rect 11756 49308 11762 49360
rect 10226 49104 10232 49156
rect 10284 49144 10290 49156
rect 10505 49147 10563 49153
rect 10505 49144 10517 49147
rect 10284 49116 10517 49144
rect 10284 49104 10290 49116
rect 10505 49113 10517 49116
rect 10551 49113 10563 49147
rect 10505 49107 10563 49113
rect 10870 49104 10876 49156
rect 10928 49144 10934 49156
rect 11517 49147 11575 49153
rect 11517 49144 11529 49147
rect 10928 49116 11529 49144
rect 10928 49104 10934 49116
rect 11517 49113 11529 49116
rect 11563 49113 11575 49147
rect 11517 49107 11575 49113
rect 24765 49147 24823 49153
rect 24765 49113 24777 49147
rect 24811 49144 24823 49147
rect 25130 49144 25136 49156
rect 24811 49116 25136 49144
rect 24811 49113 24823 49116
rect 24765 49107 24823 49113
rect 25130 49104 25136 49116
rect 25188 49104 25194 49156
rect 20070 49036 20076 49088
rect 20128 49076 20134 49088
rect 25225 49079 25283 49085
rect 25225 49076 25237 49079
rect 20128 49048 25237 49076
rect 20128 49036 20134 49048
rect 25225 49045 25237 49048
rect 25271 49045 25283 49079
rect 25225 49039 25283 49045
rect 1104 48986 25852 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 25852 48986
rect 1104 48912 25852 48934
rect 9122 48872 9128 48884
rect 6656 48844 9128 48872
rect 6656 48745 6684 48844
rect 9122 48832 9128 48844
rect 9180 48832 9186 48884
rect 6641 48739 6699 48745
rect 6641 48705 6653 48739
rect 6687 48705 6699 48739
rect 8050 48708 8800 48736
rect 6641 48699 6699 48705
rect 6917 48671 6975 48677
rect 6917 48637 6929 48671
rect 6963 48668 6975 48671
rect 8294 48668 8300 48680
rect 6963 48640 8300 48668
rect 6963 48637 6975 48640
rect 6917 48631 6975 48637
rect 8294 48628 8300 48640
rect 8352 48628 8358 48680
rect 8386 48628 8392 48680
rect 8444 48628 8450 48680
rect 8772 48609 8800 48708
rect 8757 48603 8815 48609
rect 8757 48569 8769 48603
rect 8803 48600 8815 48603
rect 9950 48600 9956 48612
rect 8803 48572 9956 48600
rect 8803 48569 8815 48572
rect 8757 48563 8815 48569
rect 9950 48560 9956 48572
rect 10008 48560 10014 48612
rect 8941 48535 8999 48541
rect 8941 48501 8953 48535
rect 8987 48532 8999 48535
rect 9122 48532 9128 48544
rect 8987 48504 9128 48532
rect 8987 48501 8999 48504
rect 8941 48495 8999 48501
rect 9122 48492 9128 48504
rect 9180 48492 9186 48544
rect 25130 48492 25136 48544
rect 25188 48532 25194 48544
rect 25409 48535 25467 48541
rect 25409 48532 25421 48535
rect 25188 48504 25421 48532
rect 25188 48492 25194 48504
rect 25409 48501 25421 48504
rect 25455 48501 25467 48535
rect 25409 48495 25467 48501
rect 1104 48442 25852 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 25852 48442
rect 1104 48368 25852 48390
rect 7742 48084 7748 48136
rect 7800 48124 7806 48136
rect 10356 48127 10414 48133
rect 10356 48124 10368 48127
rect 7800 48096 10368 48124
rect 7800 48084 7806 48096
rect 10356 48093 10368 48096
rect 10402 48093 10414 48127
rect 10356 48087 10414 48093
rect 23382 48084 23388 48136
rect 23440 48084 23446 48136
rect 25130 48084 25136 48136
rect 25188 48084 25194 48136
rect 17586 48016 17592 48068
rect 17644 48056 17650 48068
rect 25317 48059 25375 48065
rect 25317 48056 25329 48059
rect 17644 48028 25329 48056
rect 17644 48016 17650 48028
rect 25317 48025 25329 48028
rect 25363 48025 25375 48059
rect 25317 48019 25375 48025
rect 10459 47991 10517 47997
rect 10459 47957 10471 47991
rect 10505 47988 10517 47991
rect 12618 47988 12624 48000
rect 10505 47960 12624 47988
rect 10505 47957 10517 47960
rect 10459 47951 10517 47957
rect 12618 47948 12624 47960
rect 12676 47948 12682 48000
rect 24026 47948 24032 48000
rect 24084 47948 24090 48000
rect 1104 47898 25852 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 25852 47898
rect 1104 47824 25852 47846
rect 9214 47744 9220 47796
rect 9272 47784 9278 47796
rect 9490 47784 9496 47796
rect 9272 47756 9496 47784
rect 9272 47744 9278 47756
rect 9490 47744 9496 47756
rect 9548 47784 9554 47796
rect 9861 47787 9919 47793
rect 9861 47784 9873 47787
rect 9548 47756 9873 47784
rect 9548 47744 9554 47756
rect 9861 47753 9873 47756
rect 9907 47753 9919 47787
rect 9861 47747 9919 47753
rect 8570 47676 8576 47728
rect 8628 47716 8634 47728
rect 10137 47719 10195 47725
rect 10137 47716 10149 47719
rect 8628 47688 10149 47716
rect 8628 47676 8634 47688
rect 9416 47657 9444 47688
rect 10137 47685 10149 47688
rect 10183 47716 10195 47719
rect 10962 47716 10968 47728
rect 10183 47688 10968 47716
rect 10183 47685 10195 47688
rect 10137 47679 10195 47685
rect 10962 47676 10968 47688
rect 11020 47676 11026 47728
rect 9401 47651 9459 47657
rect 9401 47617 9413 47651
rect 9447 47648 9459 47651
rect 24857 47651 24915 47657
rect 9447 47620 9481 47648
rect 9447 47617 9459 47620
rect 9401 47611 9459 47617
rect 24857 47617 24869 47651
rect 24903 47648 24915 47651
rect 25314 47648 25320 47660
rect 24903 47620 25320 47648
rect 24903 47617 24915 47620
rect 24857 47611 24915 47617
rect 25314 47608 25320 47620
rect 25372 47608 25378 47660
rect 8294 47404 8300 47456
rect 8352 47444 8358 47456
rect 9490 47444 9496 47456
rect 8352 47416 9496 47444
rect 8352 47404 8358 47416
rect 9490 47404 9496 47416
rect 9548 47404 9554 47456
rect 24946 47404 24952 47456
rect 25004 47444 25010 47456
rect 25133 47447 25191 47453
rect 25133 47444 25145 47447
rect 25004 47416 25145 47444
rect 25004 47404 25010 47416
rect 25133 47413 25145 47416
rect 25179 47413 25191 47447
rect 25133 47407 25191 47413
rect 1104 47354 25852 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 25852 47354
rect 1104 47280 25852 47302
rect 9214 46996 9220 47048
rect 9272 47036 9278 47048
rect 11644 47039 11702 47045
rect 11644 47036 11656 47039
rect 9272 47008 11656 47036
rect 9272 46996 9278 47008
rect 11644 47005 11656 47008
rect 11690 47005 11702 47039
rect 11644 46999 11702 47005
rect 11747 46971 11805 46977
rect 11747 46937 11759 46971
rect 11793 46968 11805 46971
rect 13722 46968 13728 46980
rect 11793 46940 13728 46968
rect 11793 46937 11805 46940
rect 11747 46931 11805 46937
rect 13722 46928 13728 46940
rect 13780 46928 13786 46980
rect 25314 46860 25320 46912
rect 25372 46900 25378 46912
rect 25409 46903 25467 46909
rect 25409 46900 25421 46903
rect 25372 46872 25421 46900
rect 25372 46860 25378 46872
rect 25409 46869 25421 46872
rect 25455 46869 25467 46903
rect 25409 46863 25467 46869
rect 1104 46810 25852 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 25852 46810
rect 1104 46736 25852 46758
rect 10778 46656 10784 46708
rect 10836 46656 10842 46708
rect 10962 46656 10968 46708
rect 11020 46696 11026 46708
rect 11057 46699 11115 46705
rect 11057 46696 11069 46699
rect 11020 46668 11069 46696
rect 11020 46656 11026 46668
rect 11057 46665 11069 46668
rect 11103 46665 11115 46699
rect 11057 46659 11115 46665
rect 10980 46628 11008 46656
rect 10336 46600 11008 46628
rect 10336 46569 10364 46600
rect 10321 46563 10379 46569
rect 10321 46529 10333 46563
rect 10367 46529 10379 46563
rect 10321 46523 10379 46529
rect 10704 46424 10732 46600
rect 13722 46588 13728 46640
rect 13780 46628 13786 46640
rect 14093 46631 14151 46637
rect 14093 46628 14105 46631
rect 13780 46600 14105 46628
rect 13780 46588 13786 46600
rect 14093 46597 14105 46600
rect 14139 46597 14151 46631
rect 14093 46591 14151 46597
rect 10778 46520 10784 46572
rect 10836 46560 10842 46572
rect 12564 46563 12622 46569
rect 12564 46560 12576 46563
rect 10836 46532 12576 46560
rect 10836 46520 10842 46532
rect 12564 46529 12576 46532
rect 12610 46529 12622 46563
rect 12564 46523 12622 46529
rect 13906 46520 13912 46572
rect 13964 46520 13970 46572
rect 25314 46520 25320 46572
rect 25372 46520 25378 46572
rect 15746 46452 15752 46504
rect 15804 46452 15810 46504
rect 10778 46424 10784 46436
rect 10704 46396 10784 46424
rect 10778 46384 10784 46396
rect 10836 46384 10842 46436
rect 10410 46316 10416 46368
rect 10468 46316 10474 46368
rect 12667 46359 12725 46365
rect 12667 46325 12679 46359
rect 12713 46356 12725 46359
rect 15010 46356 15016 46368
rect 12713 46328 15016 46356
rect 12713 46325 12725 46328
rect 12667 46319 12725 46325
rect 15010 46316 15016 46328
rect 15068 46316 15074 46368
rect 25133 46359 25191 46365
rect 25133 46325 25145 46359
rect 25179 46356 25191 46359
rect 25682 46356 25688 46368
rect 25179 46328 25688 46356
rect 25179 46325 25191 46328
rect 25133 46319 25191 46325
rect 25682 46316 25688 46328
rect 25740 46316 25746 46368
rect 1104 46266 25852 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 25852 46266
rect 1104 46192 25852 46214
rect 8478 46112 8484 46164
rect 8536 46112 8542 46164
rect 15562 46084 15568 46096
rect 14844 46056 15568 46084
rect 7742 45976 7748 46028
rect 7800 46016 7806 46028
rect 14844 46025 14872 46056
rect 15562 46044 15568 46056
rect 15620 46044 15626 46096
rect 8113 46019 8171 46025
rect 8113 46016 8125 46019
rect 7800 45988 8125 46016
rect 7800 45976 7806 45988
rect 8113 45985 8125 45988
rect 8159 45985 8171 46019
rect 8113 45979 8171 45985
rect 14829 46019 14887 46025
rect 14829 45985 14841 46019
rect 14875 45985 14887 46019
rect 14829 45979 14887 45985
rect 15010 45976 15016 46028
rect 15068 45976 15074 46028
rect 16482 45976 16488 46028
rect 16540 45976 16546 46028
rect 7834 45908 7840 45960
rect 7892 45948 7898 45960
rect 7929 45951 7987 45957
rect 7929 45948 7941 45951
rect 7892 45920 7941 45948
rect 7892 45908 7898 45920
rect 7929 45917 7941 45920
rect 7975 45917 7987 45951
rect 7929 45911 7987 45917
rect 12526 45908 12532 45960
rect 12584 45948 12590 45960
rect 13300 45951 13358 45957
rect 13300 45948 13312 45951
rect 12584 45920 13312 45948
rect 12584 45908 12590 45920
rect 13300 45917 13312 45920
rect 13346 45917 13358 45951
rect 13300 45911 13358 45917
rect 24857 45951 24915 45957
rect 24857 45917 24869 45951
rect 24903 45948 24915 45951
rect 25314 45948 25320 45960
rect 24903 45920 25320 45948
rect 24903 45917 24915 45920
rect 24857 45911 24915 45917
rect 25314 45908 25320 45920
rect 25372 45908 25378 45960
rect 13403 45815 13461 45821
rect 13403 45781 13415 45815
rect 13449 45812 13461 45815
rect 15102 45812 15108 45824
rect 13449 45784 15108 45812
rect 13449 45781 13461 45784
rect 13403 45775 13461 45781
rect 15102 45772 15108 45784
rect 15160 45772 15166 45824
rect 25133 45815 25191 45821
rect 25133 45781 25145 45815
rect 25179 45812 25191 45815
rect 26050 45812 26056 45824
rect 25179 45784 26056 45812
rect 25179 45781 25191 45784
rect 25133 45775 25191 45781
rect 26050 45772 26056 45784
rect 26108 45772 26114 45824
rect 1104 45722 25852 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 25852 45722
rect 1104 45648 25852 45670
rect 10502 45500 10508 45552
rect 10560 45540 10566 45552
rect 12526 45540 12532 45552
rect 10560 45512 12532 45540
rect 10560 45500 10566 45512
rect 12526 45500 12532 45512
rect 12584 45500 12590 45552
rect 12618 45500 12624 45552
rect 12676 45540 12682 45552
rect 12897 45543 12955 45549
rect 12897 45540 12909 45543
rect 12676 45512 12909 45540
rect 12676 45500 12682 45512
rect 12897 45509 12909 45512
rect 12943 45509 12955 45543
rect 12897 45503 12955 45509
rect 12710 45432 12716 45484
rect 12768 45432 12774 45484
rect 14550 45364 14556 45416
rect 14608 45364 14614 45416
rect 25314 45228 25320 45280
rect 25372 45268 25378 45280
rect 25409 45271 25467 45277
rect 25409 45268 25421 45271
rect 25372 45240 25421 45268
rect 25372 45228 25378 45240
rect 25409 45237 25421 45240
rect 25455 45237 25467 45271
rect 25409 45231 25467 45237
rect 1104 45178 25852 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 25852 45178
rect 1104 45104 25852 45126
rect 9490 45024 9496 45076
rect 9548 45064 9554 45076
rect 10873 45067 10931 45073
rect 10873 45064 10885 45067
rect 9548 45036 10885 45064
rect 9548 45024 9554 45036
rect 10873 45033 10885 45036
rect 10919 45033 10931 45067
rect 10873 45027 10931 45033
rect 9950 44888 9956 44940
rect 10008 44928 10014 44940
rect 10008 44900 10640 44928
rect 10008 44888 10014 44900
rect 9122 44820 9128 44872
rect 9180 44820 9186 44872
rect 9401 44795 9459 44801
rect 9401 44761 9413 44795
rect 9447 44792 9459 44795
rect 9674 44792 9680 44804
rect 9447 44764 9680 44792
rect 9447 44761 9459 44764
rect 9401 44755 9459 44761
rect 9674 44752 9680 44764
rect 9732 44752 9738 44804
rect 10612 44792 10640 44900
rect 15654 44888 15660 44940
rect 15712 44888 15718 44940
rect 25314 44820 25320 44872
rect 25372 44820 25378 44872
rect 11241 44795 11299 44801
rect 11241 44792 11253 44795
rect 10612 44778 11253 44792
rect 10626 44764 11253 44778
rect 11241 44761 11253 44764
rect 11287 44792 11299 44795
rect 11514 44792 11520 44804
rect 11287 44764 11520 44792
rect 11287 44761 11299 44764
rect 11241 44755 11299 44761
rect 11514 44752 11520 44764
rect 11572 44752 11578 44804
rect 15102 44752 15108 44804
rect 15160 44792 15166 44804
rect 15841 44795 15899 44801
rect 15841 44792 15853 44795
rect 15160 44764 15853 44792
rect 15160 44752 15166 44764
rect 15841 44761 15853 44764
rect 15887 44761 15899 44795
rect 15841 44755 15899 44761
rect 17497 44795 17555 44801
rect 17497 44761 17509 44795
rect 17543 44792 17555 44795
rect 19978 44792 19984 44804
rect 17543 44764 19984 44792
rect 17543 44761 17555 44764
rect 17497 44755 17555 44761
rect 19978 44752 19984 44764
rect 20036 44752 20042 44804
rect 9692 44724 9720 44752
rect 10410 44724 10416 44736
rect 9692 44696 10416 44724
rect 10410 44684 10416 44696
rect 10468 44684 10474 44736
rect 11425 44727 11483 44733
rect 11425 44693 11437 44727
rect 11471 44724 11483 44727
rect 11698 44724 11704 44736
rect 11471 44696 11704 44724
rect 11471 44693 11483 44696
rect 11425 44687 11483 44693
rect 11698 44684 11704 44696
rect 11756 44684 11762 44736
rect 25133 44727 25191 44733
rect 25133 44693 25145 44727
rect 25179 44724 25191 44727
rect 25222 44724 25228 44736
rect 25179 44696 25228 44724
rect 25179 44693 25191 44696
rect 25133 44687 25191 44693
rect 25222 44684 25228 44696
rect 25280 44684 25286 44736
rect 1104 44634 25852 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 25852 44634
rect 1104 44560 25852 44582
rect 9582 44480 9588 44532
rect 9640 44480 9646 44532
rect 9125 44387 9183 44393
rect 9125 44353 9137 44387
rect 9171 44384 9183 44387
rect 9214 44384 9220 44396
rect 9171 44356 9220 44384
rect 9171 44353 9183 44356
rect 9125 44347 9183 44353
rect 9214 44344 9220 44356
rect 9272 44344 9278 44396
rect 10597 44387 10655 44393
rect 10597 44353 10609 44387
rect 10643 44384 10655 44387
rect 10778 44384 10784 44396
rect 10643 44356 10784 44384
rect 10643 44353 10655 44356
rect 10597 44347 10655 44353
rect 10778 44344 10784 44356
rect 10836 44384 10842 44396
rect 11517 44387 11575 44393
rect 11517 44384 11529 44387
rect 10836 44356 11529 44384
rect 10836 44344 10842 44356
rect 11517 44353 11529 44356
rect 11563 44353 11575 44387
rect 11517 44347 11575 44353
rect 24762 44344 24768 44396
rect 24820 44384 24826 44396
rect 25133 44387 25191 44393
rect 25133 44384 25145 44387
rect 24820 44356 25145 44384
rect 24820 44344 24826 44356
rect 25133 44353 25145 44356
rect 25179 44353 25191 44387
rect 25133 44347 25191 44353
rect 8941 44319 8999 44325
rect 8941 44285 8953 44319
rect 8987 44316 8999 44319
rect 9030 44316 9036 44328
rect 8987 44288 9036 44316
rect 8987 44285 8999 44288
rect 8941 44279 8999 44285
rect 9030 44276 9036 44288
rect 9088 44276 9094 44328
rect 10502 44208 10508 44260
rect 10560 44248 10566 44260
rect 10560 44220 11008 44248
rect 10560 44208 10566 44220
rect 10980 44192 11008 44220
rect 10686 44140 10692 44192
rect 10744 44140 10750 44192
rect 10962 44140 10968 44192
rect 11020 44180 11026 44192
rect 11057 44183 11115 44189
rect 11057 44180 11069 44183
rect 11020 44152 11069 44180
rect 11020 44140 11026 44152
rect 11057 44149 11069 44152
rect 11103 44149 11115 44183
rect 11057 44143 11115 44149
rect 16850 44140 16856 44192
rect 16908 44180 16914 44192
rect 22830 44180 22836 44192
rect 16908 44152 22836 44180
rect 16908 44140 16914 44152
rect 22830 44140 22836 44152
rect 22888 44140 22894 44192
rect 24854 44140 24860 44192
rect 24912 44180 24918 44192
rect 25225 44183 25283 44189
rect 25225 44180 25237 44183
rect 24912 44152 25237 44180
rect 24912 44140 24918 44152
rect 25225 44149 25237 44152
rect 25271 44149 25283 44183
rect 25225 44143 25283 44149
rect 1104 44090 25852 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 25852 44090
rect 1104 44016 25852 44038
rect 16574 43936 16580 43988
rect 16632 43976 16638 43988
rect 22097 43979 22155 43985
rect 22097 43976 22109 43979
rect 16632 43948 22109 43976
rect 16632 43936 16638 43948
rect 22097 43945 22109 43948
rect 22143 43945 22155 43979
rect 22097 43939 22155 43945
rect 20625 43843 20683 43849
rect 20625 43809 20637 43843
rect 20671 43840 20683 43843
rect 24026 43840 24032 43852
rect 20671 43812 24032 43840
rect 20671 43809 20683 43812
rect 20625 43803 20683 43809
rect 24026 43800 24032 43812
rect 24084 43800 24090 43852
rect 19518 43732 19524 43784
rect 19576 43772 19582 43784
rect 20349 43775 20407 43781
rect 20349 43772 20361 43775
rect 19576 43744 20361 43772
rect 19576 43732 19582 43744
rect 20349 43741 20361 43744
rect 20395 43741 20407 43775
rect 20349 43735 20407 43741
rect 21082 43704 21088 43716
rect 21008 43676 21088 43704
rect 21008 43636 21036 43676
rect 21082 43664 21088 43676
rect 21140 43664 21146 43716
rect 22373 43707 22431 43713
rect 22373 43704 22385 43707
rect 21928 43676 22385 43704
rect 21928 43636 21956 43676
rect 22373 43673 22385 43676
rect 22419 43673 22431 43707
rect 22373 43667 22431 43673
rect 21008 43608 21956 43636
rect 25498 43596 25504 43648
rect 25556 43596 25562 43648
rect 1104 43546 25852 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 25852 43546
rect 1104 43472 25852 43494
rect 25133 43367 25191 43373
rect 25133 43333 25145 43367
rect 25179 43364 25191 43367
rect 25498 43364 25504 43376
rect 25179 43336 25504 43364
rect 25179 43333 25191 43336
rect 25133 43327 25191 43333
rect 25498 43324 25504 43336
rect 25556 43324 25562 43376
rect 24210 43052 24216 43104
rect 24268 43092 24274 43104
rect 25225 43095 25283 43101
rect 25225 43092 25237 43095
rect 24268 43064 25237 43092
rect 24268 43052 24274 43064
rect 25225 43061 25237 43064
rect 25271 43061 25283 43095
rect 25225 43055 25283 43061
rect 1104 43002 25852 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 25852 43002
rect 1104 42928 25852 42950
rect 10226 42712 10232 42764
rect 10284 42712 10290 42764
rect 8938 42644 8944 42696
rect 8996 42684 9002 42696
rect 9585 42687 9643 42693
rect 9585 42684 9597 42687
rect 8996 42656 9597 42684
rect 8996 42644 9002 42656
rect 9585 42653 9597 42656
rect 9631 42653 9643 42687
rect 9585 42647 9643 42653
rect 9769 42687 9827 42693
rect 9769 42653 9781 42687
rect 9815 42684 9827 42687
rect 10594 42684 10600 42696
rect 9815 42656 10600 42684
rect 9815 42653 9827 42656
rect 9769 42647 9827 42653
rect 10594 42644 10600 42656
rect 10652 42644 10658 42696
rect 24765 42619 24823 42625
rect 24765 42585 24777 42619
rect 24811 42616 24823 42619
rect 25130 42616 25136 42628
rect 24811 42588 25136 42616
rect 24811 42585 24823 42588
rect 24765 42579 24823 42585
rect 25130 42576 25136 42588
rect 25188 42576 25194 42628
rect 24302 42508 24308 42560
rect 24360 42548 24366 42560
rect 25225 42551 25283 42557
rect 25225 42548 25237 42551
rect 24360 42520 25237 42548
rect 24360 42508 24366 42520
rect 25225 42517 25237 42520
rect 25271 42517 25283 42551
rect 25225 42511 25283 42517
rect 1104 42458 25852 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 25852 42458
rect 1104 42384 25852 42406
rect 9674 42304 9680 42356
rect 9732 42344 9738 42356
rect 11149 42347 11207 42353
rect 11149 42344 11161 42347
rect 9732 42316 11161 42344
rect 9732 42304 9738 42316
rect 11149 42313 11161 42316
rect 11195 42313 11207 42347
rect 11149 42307 11207 42313
rect 11514 42276 11520 42288
rect 10902 42248 11520 42276
rect 11514 42236 11520 42248
rect 11572 42236 11578 42288
rect 9122 42100 9128 42152
rect 9180 42140 9186 42152
rect 9401 42143 9459 42149
rect 9401 42140 9413 42143
rect 9180 42112 9413 42140
rect 9180 42100 9186 42112
rect 9401 42109 9413 42112
rect 9447 42109 9459 42143
rect 9401 42103 9459 42109
rect 9677 42143 9735 42149
rect 9677 42109 9689 42143
rect 9723 42140 9735 42143
rect 9766 42140 9772 42152
rect 9723 42112 9772 42140
rect 9723 42109 9735 42112
rect 9677 42103 9735 42109
rect 9416 42004 9444 42103
rect 9766 42100 9772 42112
rect 9824 42140 9830 42152
rect 10686 42140 10692 42152
rect 9824 42112 10692 42140
rect 9824 42100 9830 42112
rect 10686 42100 10692 42112
rect 10744 42100 10750 42152
rect 10704 42044 11744 42072
rect 10704 42004 10732 42044
rect 11716 42016 11744 42044
rect 15562 42032 15568 42084
rect 15620 42072 15626 42084
rect 24486 42072 24492 42084
rect 15620 42044 24492 42072
rect 15620 42032 15626 42044
rect 24486 42032 24492 42044
rect 24544 42032 24550 42084
rect 9416 41976 10732 42004
rect 11514 41964 11520 42016
rect 11572 41964 11578 42016
rect 11698 41964 11704 42016
rect 11756 41964 11762 42016
rect 25130 41964 25136 42016
rect 25188 42004 25194 42016
rect 25409 42007 25467 42013
rect 25409 42004 25421 42007
rect 25188 41976 25421 42004
rect 25188 41964 25194 41976
rect 25409 41973 25421 41976
rect 25455 41973 25467 42007
rect 25409 41967 25467 41973
rect 1104 41914 25852 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 25852 41914
rect 1104 41840 25852 41862
rect 10870 41760 10876 41812
rect 10928 41760 10934 41812
rect 16206 41692 16212 41744
rect 16264 41732 16270 41744
rect 18690 41732 18696 41744
rect 16264 41704 18696 41732
rect 16264 41692 16270 41704
rect 18690 41692 18696 41704
rect 18748 41692 18754 41744
rect 10413 41667 10471 41673
rect 10413 41633 10425 41667
rect 10459 41664 10471 41667
rect 10962 41664 10968 41676
rect 10459 41636 10968 41664
rect 10459 41633 10471 41636
rect 10413 41627 10471 41633
rect 10962 41624 10968 41636
rect 11020 41624 11026 41676
rect 10226 41556 10232 41608
rect 10284 41556 10290 41608
rect 25130 41556 25136 41608
rect 25188 41556 25194 41608
rect 21358 41488 21364 41540
rect 21416 41528 21422 41540
rect 25317 41531 25375 41537
rect 25317 41528 25329 41531
rect 21416 41500 25329 41528
rect 21416 41488 21422 41500
rect 25317 41497 25329 41500
rect 25363 41497 25375 41531
rect 25317 41491 25375 41497
rect 20254 41420 20260 41472
rect 20312 41460 20318 41472
rect 24670 41460 24676 41472
rect 20312 41432 24676 41460
rect 20312 41420 20318 41432
rect 24670 41420 24676 41432
rect 24728 41420 24734 41472
rect 1104 41370 25852 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 25852 41370
rect 1104 41296 25852 41318
rect 24857 41123 24915 41129
rect 24857 41089 24869 41123
rect 24903 41120 24915 41123
rect 25314 41120 25320 41132
rect 24903 41092 25320 41120
rect 24903 41089 24915 41092
rect 24857 41083 24915 41089
rect 25314 41080 25320 41092
rect 25372 41080 25378 41132
rect 25038 40876 25044 40928
rect 25096 40916 25102 40928
rect 25133 40919 25191 40925
rect 25133 40916 25145 40919
rect 25096 40888 25145 40916
rect 25096 40876 25102 40888
rect 25133 40885 25145 40888
rect 25179 40885 25191 40919
rect 25133 40879 25191 40885
rect 1104 40826 25852 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 25852 40826
rect 1104 40752 25852 40774
rect 25498 40332 25504 40384
rect 25556 40332 25562 40384
rect 1104 40282 25852 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 25852 40282
rect 1104 40208 25852 40230
rect 23290 40128 23296 40180
rect 23348 40168 23354 40180
rect 25133 40171 25191 40177
rect 25133 40168 25145 40171
rect 23348 40140 25145 40168
rect 23348 40128 23354 40140
rect 25133 40137 25145 40140
rect 25179 40137 25191 40171
rect 25133 40131 25191 40137
rect 25498 40100 25504 40112
rect 25332 40072 25504 40100
rect 25332 40041 25360 40072
rect 25498 40060 25504 40072
rect 25556 40060 25562 40112
rect 25317 40035 25375 40041
rect 25317 40001 25329 40035
rect 25363 40001 25375 40035
rect 25317 39995 25375 40001
rect 1104 39738 25852 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 25852 39738
rect 1104 39664 25852 39686
rect 24857 39423 24915 39429
rect 24857 39389 24869 39423
rect 24903 39420 24915 39423
rect 25314 39420 25320 39432
rect 24903 39392 25320 39420
rect 24903 39389 24915 39392
rect 24857 39383 24915 39389
rect 25314 39380 25320 39392
rect 25372 39380 25378 39432
rect 21910 39244 21916 39296
rect 21968 39284 21974 39296
rect 25133 39287 25191 39293
rect 25133 39284 25145 39287
rect 21968 39256 25145 39284
rect 21968 39244 21974 39256
rect 25133 39253 25145 39256
rect 25179 39253 25191 39287
rect 25133 39247 25191 39253
rect 1104 39194 25852 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 25852 39194
rect 1104 39120 25852 39142
rect 25314 38700 25320 38752
rect 25372 38740 25378 38752
rect 25409 38743 25467 38749
rect 25409 38740 25421 38743
rect 25372 38712 25421 38740
rect 25372 38700 25378 38712
rect 25409 38709 25421 38712
rect 25455 38709 25467 38743
rect 25409 38703 25467 38709
rect 1104 38650 25852 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 25852 38650
rect 1104 38576 25852 38598
rect 25314 38292 25320 38344
rect 25372 38292 25378 38344
rect 25133 38199 25191 38205
rect 25133 38165 25145 38199
rect 25179 38196 25191 38199
rect 25406 38196 25412 38208
rect 25179 38168 25412 38196
rect 25179 38165 25191 38168
rect 25133 38159 25191 38165
rect 25406 38156 25412 38168
rect 25464 38156 25470 38208
rect 1104 38106 25852 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 25852 38106
rect 1104 38032 25852 38054
rect 7834 37952 7840 38004
rect 7892 37992 7898 38004
rect 8665 37995 8723 38001
rect 8665 37992 8677 37995
rect 7892 37964 8677 37992
rect 7892 37952 7898 37964
rect 8665 37961 8677 37964
rect 8711 37961 8723 37995
rect 8665 37955 8723 37961
rect 8846 37816 8852 37868
rect 8904 37816 8910 37868
rect 24765 37859 24823 37865
rect 24765 37825 24777 37859
rect 24811 37856 24823 37859
rect 25130 37856 25136 37868
rect 24811 37828 25136 37856
rect 24811 37825 24823 37828
rect 24765 37819 24823 37825
rect 25130 37816 25136 37828
rect 25188 37816 25194 37868
rect 25317 37723 25375 37729
rect 25317 37689 25329 37723
rect 25363 37720 25375 37723
rect 25774 37720 25780 37732
rect 25363 37692 25780 37720
rect 25363 37689 25375 37692
rect 25317 37683 25375 37689
rect 25774 37680 25780 37692
rect 25832 37680 25838 37732
rect 1104 37562 25852 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 25852 37562
rect 1104 37488 25852 37510
rect 16298 37272 16304 37324
rect 16356 37312 16362 37324
rect 18598 37312 18604 37324
rect 16356 37284 18604 37312
rect 16356 37272 16362 37284
rect 18598 37272 18604 37284
rect 18656 37272 18662 37324
rect 25498 37068 25504 37120
rect 25556 37068 25562 37120
rect 1104 37018 25852 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 25852 37018
rect 1104 36944 25852 36966
rect 25133 36839 25191 36845
rect 25133 36805 25145 36839
rect 25179 36836 25191 36839
rect 25498 36836 25504 36848
rect 25179 36808 25504 36836
rect 25179 36805 25191 36808
rect 25133 36799 25191 36805
rect 25498 36796 25504 36808
rect 25556 36796 25562 36848
rect 25317 36635 25375 36641
rect 25317 36601 25329 36635
rect 25363 36632 25375 36635
rect 25590 36632 25596 36644
rect 25363 36604 25596 36632
rect 25363 36601 25375 36604
rect 25317 36595 25375 36601
rect 25590 36592 25596 36604
rect 25648 36592 25654 36644
rect 1104 36474 25852 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 25852 36474
rect 1104 36400 25852 36422
rect 24857 36159 24915 36165
rect 24857 36125 24869 36159
rect 24903 36156 24915 36159
rect 25314 36156 25320 36168
rect 24903 36128 25320 36156
rect 24903 36125 24915 36128
rect 24857 36119 24915 36125
rect 25314 36116 25320 36128
rect 25372 36116 25378 36168
rect 25130 35980 25136 36032
rect 25188 35980 25194 36032
rect 1104 35930 25852 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 25852 35930
rect 1104 35856 25852 35878
rect 11698 35816 11704 35828
rect 9416 35788 11704 35816
rect 9416 35689 9444 35788
rect 11698 35776 11704 35788
rect 11756 35776 11762 35828
rect 22465 35819 22523 35825
rect 22465 35785 22477 35819
rect 22511 35816 22523 35819
rect 26050 35816 26056 35828
rect 22511 35788 26056 35816
rect 22511 35785 22523 35788
rect 22465 35779 22523 35785
rect 26050 35776 26056 35788
rect 26108 35776 26114 35828
rect 11514 35748 11520 35760
rect 10902 35720 11520 35748
rect 11514 35708 11520 35720
rect 11572 35748 11578 35760
rect 12158 35748 12164 35760
rect 11572 35720 12164 35748
rect 11572 35708 11578 35720
rect 12158 35708 12164 35720
rect 12216 35708 12222 35760
rect 21177 35751 21235 35757
rect 21177 35717 21189 35751
rect 21223 35748 21235 35751
rect 25682 35748 25688 35760
rect 21223 35720 25688 35748
rect 21223 35717 21235 35720
rect 21177 35711 21235 35717
rect 25682 35708 25688 35720
rect 25740 35708 25746 35760
rect 9401 35683 9459 35689
rect 9401 35649 9413 35683
rect 9447 35649 9459 35683
rect 21085 35683 21143 35689
rect 21085 35680 21097 35683
rect 9401 35643 9459 35649
rect 20364 35652 21097 35680
rect 9674 35572 9680 35624
rect 9732 35572 9738 35624
rect 9766 35572 9772 35624
rect 9824 35612 9830 35624
rect 11149 35615 11207 35621
rect 11149 35612 11161 35615
rect 9824 35584 11161 35612
rect 9824 35572 9830 35584
rect 11149 35581 11161 35584
rect 11195 35581 11207 35615
rect 11149 35575 11207 35581
rect 11790 35436 11796 35488
rect 11848 35436 11854 35488
rect 15746 35436 15752 35488
rect 15804 35476 15810 35488
rect 20364 35485 20392 35652
rect 21085 35649 21097 35652
rect 21131 35680 21143 35683
rect 21131 35652 21772 35680
rect 21131 35649 21143 35652
rect 21085 35643 21143 35649
rect 21269 35615 21327 35621
rect 21269 35581 21281 35615
rect 21315 35581 21327 35615
rect 21744 35612 21772 35652
rect 21818 35640 21824 35692
rect 21876 35680 21882 35692
rect 22373 35683 22431 35689
rect 22373 35680 22385 35683
rect 21876 35652 22385 35680
rect 21876 35640 21882 35652
rect 22373 35649 22385 35652
rect 22419 35649 22431 35683
rect 22373 35643 22431 35649
rect 22186 35612 22192 35624
rect 21744 35584 22192 35612
rect 21269 35575 21327 35581
rect 21284 35544 21312 35575
rect 22186 35572 22192 35584
rect 22244 35572 22250 35624
rect 22554 35572 22560 35624
rect 22612 35572 22618 35624
rect 21192 35516 21312 35544
rect 21192 35488 21220 35516
rect 20349 35479 20407 35485
rect 20349 35476 20361 35479
rect 15804 35448 20361 35476
rect 15804 35436 15810 35448
rect 20349 35445 20361 35448
rect 20395 35445 20407 35479
rect 20349 35439 20407 35445
rect 20622 35436 20628 35488
rect 20680 35476 20686 35488
rect 20717 35479 20775 35485
rect 20717 35476 20729 35479
rect 20680 35448 20729 35476
rect 20680 35436 20686 35448
rect 20717 35445 20729 35448
rect 20763 35445 20775 35479
rect 20717 35439 20775 35445
rect 21174 35436 21180 35488
rect 21232 35436 21238 35488
rect 22002 35436 22008 35488
rect 22060 35436 22066 35488
rect 25314 35436 25320 35488
rect 25372 35476 25378 35488
rect 25409 35479 25467 35485
rect 25409 35476 25421 35479
rect 25372 35448 25421 35476
rect 25372 35436 25378 35448
rect 25409 35445 25421 35448
rect 25455 35445 25467 35479
rect 25409 35439 25467 35445
rect 1104 35386 25852 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 25852 35386
rect 1104 35312 25852 35334
rect 22738 35096 22744 35148
rect 22796 35136 22802 35148
rect 23293 35139 23351 35145
rect 23293 35136 23305 35139
rect 22796 35108 23305 35136
rect 22796 35096 22802 35108
rect 23293 35105 23305 35108
rect 23339 35105 23351 35139
rect 23293 35099 23351 35105
rect 23201 35071 23259 35077
rect 23201 35037 23213 35071
rect 23247 35068 23259 35071
rect 25222 35068 25228 35080
rect 23247 35040 25228 35068
rect 23247 35037 23259 35040
rect 23201 35031 23259 35037
rect 25222 35028 25228 35040
rect 25280 35028 25286 35080
rect 25314 35028 25320 35080
rect 25372 35028 25378 35080
rect 19978 34960 19984 35012
rect 20036 35000 20042 35012
rect 20438 35000 20444 35012
rect 20036 34972 20444 35000
rect 20036 34960 20042 34972
rect 20438 34960 20444 34972
rect 20496 35000 20502 35012
rect 22373 35003 22431 35009
rect 22373 35000 22385 35003
rect 20496 34972 22385 35000
rect 20496 34960 20502 34972
rect 22373 34969 22385 34972
rect 22419 35000 22431 35003
rect 23109 35003 23167 35009
rect 23109 35000 23121 35003
rect 22419 34972 23121 35000
rect 22419 34969 22431 34972
rect 22373 34963 22431 34969
rect 23109 34969 23121 34972
rect 23155 34969 23167 35003
rect 23109 34963 23167 34969
rect 16482 34892 16488 34944
rect 16540 34932 16546 34944
rect 21818 34932 21824 34944
rect 16540 34904 21824 34932
rect 16540 34892 16546 34904
rect 21818 34892 21824 34904
rect 21876 34892 21882 34944
rect 22462 34892 22468 34944
rect 22520 34932 22526 34944
rect 22741 34935 22799 34941
rect 22741 34932 22753 34935
rect 22520 34904 22753 34932
rect 22520 34892 22526 34904
rect 22741 34901 22753 34904
rect 22787 34901 22799 34935
rect 22741 34895 22799 34901
rect 25133 34935 25191 34941
rect 25133 34901 25145 34935
rect 25179 34932 25191 34935
rect 25682 34932 25688 34944
rect 25179 34904 25688 34932
rect 25179 34901 25191 34904
rect 25133 34895 25191 34901
rect 25682 34892 25688 34904
rect 25740 34892 25746 34944
rect 1104 34842 25852 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 25852 34842
rect 1104 34768 25852 34790
rect 20806 34688 20812 34740
rect 20864 34728 20870 34740
rect 25133 34731 25191 34737
rect 25133 34728 25145 34731
rect 20864 34700 25145 34728
rect 20864 34688 20870 34700
rect 25133 34697 25145 34700
rect 25179 34697 25191 34731
rect 25133 34691 25191 34697
rect 24857 34595 24915 34601
rect 24857 34561 24869 34595
rect 24903 34592 24915 34595
rect 25314 34592 25320 34604
rect 24903 34564 25320 34592
rect 24903 34561 24915 34564
rect 24857 34555 24915 34561
rect 25314 34552 25320 34564
rect 25372 34552 25378 34604
rect 21082 34348 21088 34400
rect 21140 34388 21146 34400
rect 21358 34388 21364 34400
rect 21140 34360 21364 34388
rect 21140 34348 21146 34360
rect 21358 34348 21364 34360
rect 21416 34348 21422 34400
rect 1104 34298 25852 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 25852 34298
rect 1104 34224 25852 34246
rect 9030 34144 9036 34196
rect 9088 34184 9094 34196
rect 9125 34187 9183 34193
rect 9125 34184 9137 34187
rect 9088 34156 9137 34184
rect 9088 34144 9094 34156
rect 9125 34153 9137 34156
rect 9171 34153 9183 34187
rect 9125 34147 9183 34153
rect 11790 34008 11796 34060
rect 11848 34048 11854 34060
rect 15381 34051 15439 34057
rect 15381 34048 15393 34051
rect 11848 34020 15393 34048
rect 11848 34008 11854 34020
rect 15381 34017 15393 34020
rect 15427 34017 15439 34051
rect 15381 34011 15439 34017
rect 19702 34008 19708 34060
rect 19760 34048 19766 34060
rect 21637 34051 21695 34057
rect 21637 34048 21649 34051
rect 19760 34020 21649 34048
rect 19760 34008 19766 34020
rect 21637 34017 21649 34020
rect 21683 34048 21695 34051
rect 22278 34048 22284 34060
rect 21683 34020 22284 34048
rect 21683 34017 21695 34020
rect 21637 34011 21695 34017
rect 22278 34008 22284 34020
rect 22336 34008 22342 34060
rect 9214 33940 9220 33992
rect 9272 33980 9278 33992
rect 9309 33983 9367 33989
rect 9309 33980 9321 33983
rect 9272 33952 9321 33980
rect 9272 33940 9278 33952
rect 9309 33949 9321 33952
rect 9355 33949 9367 33983
rect 9309 33943 9367 33949
rect 19426 33940 19432 33992
rect 19484 33940 19490 33992
rect 24857 33983 24915 33989
rect 24857 33949 24869 33983
rect 24903 33980 24915 33983
rect 25314 33980 25320 33992
rect 24903 33952 25320 33980
rect 24903 33949 24915 33952
rect 24857 33943 24915 33949
rect 25314 33940 25320 33952
rect 25372 33940 25378 33992
rect 14645 33915 14703 33921
rect 14645 33881 14657 33915
rect 14691 33912 14703 33915
rect 15378 33912 15384 33924
rect 14691 33884 15384 33912
rect 14691 33881 14703 33884
rect 14645 33875 14703 33881
rect 15378 33872 15384 33884
rect 15436 33912 15442 33924
rect 15841 33915 15899 33921
rect 15841 33912 15853 33915
rect 15436 33884 15853 33912
rect 15436 33872 15442 33884
rect 15841 33881 15853 33884
rect 15887 33881 15899 33915
rect 15841 33875 15899 33881
rect 19705 33915 19763 33921
rect 19705 33881 19717 33915
rect 19751 33912 19763 33915
rect 19794 33912 19800 33924
rect 19751 33884 19800 33912
rect 19751 33881 19763 33884
rect 19705 33875 19763 33881
rect 19794 33872 19800 33884
rect 19852 33872 19858 33924
rect 21358 33912 21364 33924
rect 20930 33884 21364 33912
rect 21358 33872 21364 33884
rect 21416 33872 21422 33924
rect 21913 33915 21971 33921
rect 21913 33881 21925 33915
rect 21959 33881 21971 33915
rect 23138 33884 23704 33912
rect 21913 33875 21971 33881
rect 21174 33804 21180 33856
rect 21232 33804 21238 33856
rect 21928 33844 21956 33875
rect 23676 33856 23704 33884
rect 22922 33844 22928 33856
rect 21928 33816 22928 33844
rect 22922 33804 22928 33816
rect 22980 33804 22986 33856
rect 23198 33804 23204 33856
rect 23256 33844 23262 33856
rect 23385 33847 23443 33853
rect 23385 33844 23397 33847
rect 23256 33816 23397 33844
rect 23256 33804 23262 33816
rect 23385 33813 23397 33816
rect 23431 33813 23443 33847
rect 23385 33807 23443 33813
rect 23658 33804 23664 33856
rect 23716 33804 23722 33856
rect 25133 33847 25191 33853
rect 25133 33813 25145 33847
rect 25179 33844 25191 33847
rect 26234 33844 26240 33856
rect 25179 33816 26240 33844
rect 25179 33813 25191 33816
rect 25133 33807 25191 33813
rect 26234 33804 26240 33816
rect 26292 33804 26298 33856
rect 1104 33754 25852 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 25852 33754
rect 1104 33680 25852 33702
rect 22554 33640 22560 33652
rect 19812 33612 22560 33640
rect 19812 33581 19840 33612
rect 22554 33600 22560 33612
rect 22612 33640 22618 33652
rect 23198 33640 23204 33652
rect 22612 33612 23204 33640
rect 22612 33600 22618 33612
rect 23198 33600 23204 33612
rect 23256 33600 23262 33652
rect 19797 33575 19855 33581
rect 19797 33541 19809 33575
rect 19843 33541 19855 33575
rect 21358 33572 21364 33584
rect 21022 33544 21364 33572
rect 19797 33535 19855 33541
rect 21358 33532 21364 33544
rect 21416 33532 21422 33584
rect 22278 33572 22284 33584
rect 22020 33544 22284 33572
rect 19518 33464 19524 33516
rect 19576 33464 19582 33516
rect 22020 33513 22048 33544
rect 22278 33532 22284 33544
rect 22336 33532 22342 33584
rect 23658 33572 23664 33584
rect 23506 33544 23664 33572
rect 23658 33532 23664 33544
rect 23716 33532 23722 33584
rect 22005 33507 22063 33513
rect 22005 33473 22017 33507
rect 22051 33473 22063 33507
rect 25317 33507 25375 33513
rect 25317 33504 25329 33507
rect 22005 33467 22063 33473
rect 24872 33476 25329 33504
rect 19794 33396 19800 33448
rect 19852 33436 19858 33448
rect 20530 33436 20536 33448
rect 19852 33408 20536 33436
rect 19852 33396 19858 33408
rect 20530 33396 20536 33408
rect 20588 33436 20594 33448
rect 21269 33439 21327 33445
rect 21269 33436 21281 33439
rect 20588 33408 21281 33436
rect 20588 33396 20594 33408
rect 21269 33405 21281 33408
rect 21315 33405 21327 33439
rect 21269 33399 21327 33405
rect 22281 33439 22339 33445
rect 22281 33405 22293 33439
rect 22327 33436 22339 33439
rect 22370 33436 22376 33448
rect 22327 33408 22376 33436
rect 22327 33405 22339 33408
rect 22281 33399 22339 33405
rect 22370 33396 22376 33408
rect 22428 33396 22434 33448
rect 22922 33396 22928 33448
rect 22980 33436 22986 33448
rect 23753 33439 23811 33445
rect 23753 33436 23765 33439
rect 22980 33408 23765 33436
rect 22980 33396 22986 33408
rect 23753 33405 23765 33408
rect 23799 33405 23811 33439
rect 23753 33399 23811 33405
rect 21358 33260 21364 33312
rect 21416 33300 21422 33312
rect 21545 33303 21603 33309
rect 21545 33300 21557 33303
rect 21416 33272 21557 33300
rect 21416 33260 21422 33272
rect 21545 33269 21557 33272
rect 21591 33269 21603 33303
rect 21545 33263 21603 33269
rect 23658 33260 23664 33312
rect 23716 33300 23722 33312
rect 24121 33303 24179 33309
rect 24121 33300 24133 33303
rect 23716 33272 24133 33300
rect 23716 33260 23722 33272
rect 24121 33269 24133 33272
rect 24167 33300 24179 33303
rect 24305 33303 24363 33309
rect 24305 33300 24317 33303
rect 24167 33272 24317 33300
rect 24167 33269 24179 33272
rect 24121 33263 24179 33269
rect 24305 33269 24317 33272
rect 24351 33269 24363 33303
rect 24305 33263 24363 33269
rect 24581 33303 24639 33309
rect 24581 33269 24593 33303
rect 24627 33300 24639 33303
rect 24670 33300 24676 33312
rect 24627 33272 24676 33300
rect 24627 33269 24639 33272
rect 24581 33263 24639 33269
rect 24670 33260 24676 33272
rect 24728 33260 24734 33312
rect 24762 33260 24768 33312
rect 24820 33300 24826 33312
rect 24872 33309 24900 33476
rect 25317 33473 25329 33476
rect 25363 33473 25375 33507
rect 25317 33467 25375 33473
rect 24857 33303 24915 33309
rect 24857 33300 24869 33303
rect 24820 33272 24869 33300
rect 24820 33260 24826 33272
rect 24857 33269 24869 33272
rect 24903 33269 24915 33303
rect 24857 33263 24915 33269
rect 25133 33303 25191 33309
rect 25133 33269 25145 33303
rect 25179 33300 25191 33303
rect 25958 33300 25964 33312
rect 25179 33272 25964 33300
rect 25179 33269 25191 33272
rect 25133 33263 25191 33269
rect 25958 33260 25964 33272
rect 26016 33260 26022 33312
rect 1104 33210 25852 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 25852 33210
rect 1104 33136 25852 33158
rect 16758 33056 16764 33108
rect 16816 33056 16822 33108
rect 22370 33056 22376 33108
rect 22428 33096 22434 33108
rect 22738 33096 22744 33108
rect 22428 33068 22744 33096
rect 22428 33056 22434 33068
rect 22738 33056 22744 33068
rect 22796 33096 22802 33108
rect 24029 33099 24087 33105
rect 24029 33096 24041 33099
rect 22796 33068 24041 33096
rect 22796 33056 22802 33068
rect 24029 33065 24041 33068
rect 24075 33065 24087 33099
rect 24029 33059 24087 33065
rect 25314 33028 25320 33040
rect 24688 33000 25320 33028
rect 16114 32920 16120 32972
rect 16172 32960 16178 32972
rect 16574 32960 16580 32972
rect 16172 32932 16580 32960
rect 16172 32920 16178 32932
rect 16574 32920 16580 32932
rect 16632 32960 16638 32972
rect 17037 32963 17095 32969
rect 16632 32932 16677 32960
rect 16632 32920 16638 32932
rect 17037 32929 17049 32963
rect 17083 32960 17095 32963
rect 17862 32960 17868 32972
rect 17083 32932 17868 32960
rect 17083 32929 17095 32932
rect 17037 32923 17095 32929
rect 16025 32895 16083 32901
rect 16025 32861 16037 32895
rect 16071 32892 16083 32895
rect 16758 32892 16764 32904
rect 16071 32864 16764 32892
rect 16071 32861 16083 32864
rect 16025 32855 16083 32861
rect 16758 32852 16764 32864
rect 16816 32892 16822 32904
rect 17126 32892 17132 32904
rect 16816 32864 17132 32892
rect 16816 32852 16822 32864
rect 17126 32852 17132 32864
rect 17184 32852 17190 32904
rect 15933 32827 15991 32833
rect 15933 32793 15945 32827
rect 15979 32824 15991 32827
rect 17236 32824 17264 32932
rect 17862 32920 17868 32932
rect 17920 32960 17926 32972
rect 17920 32932 21956 32960
rect 17920 32920 17926 32932
rect 19426 32852 19432 32904
rect 19484 32892 19490 32904
rect 20625 32895 20683 32901
rect 20625 32892 20637 32895
rect 19484 32864 20637 32892
rect 19484 32852 19490 32864
rect 20625 32861 20637 32864
rect 20671 32861 20683 32895
rect 20625 32855 20683 32861
rect 15979 32796 17264 32824
rect 19889 32827 19947 32833
rect 15979 32793 15991 32796
rect 15933 32787 15991 32793
rect 19889 32793 19901 32827
rect 19935 32824 19947 32827
rect 19935 32796 19969 32824
rect 19935 32793 19947 32796
rect 19889 32787 19947 32793
rect 12618 32716 12624 32768
rect 12676 32756 12682 32768
rect 15565 32759 15623 32765
rect 15565 32756 15577 32759
rect 12676 32728 15577 32756
rect 12676 32716 12682 32728
rect 15565 32725 15577 32728
rect 15611 32725 15623 32759
rect 15565 32719 15623 32725
rect 17034 32716 17040 32768
rect 17092 32756 17098 32768
rect 19613 32759 19671 32765
rect 19613 32756 19625 32759
rect 17092 32728 19625 32756
rect 17092 32716 17098 32728
rect 19613 32725 19625 32728
rect 19659 32756 19671 32759
rect 19904 32756 19932 32787
rect 21818 32756 21824 32768
rect 19659 32728 21824 32756
rect 19659 32725 19671 32728
rect 19613 32719 19671 32725
rect 21818 32716 21824 32728
rect 21876 32716 21882 32768
rect 21928 32756 21956 32932
rect 22278 32920 22284 32972
rect 22336 32920 22342 32972
rect 22557 32963 22615 32969
rect 22557 32929 22569 32963
rect 22603 32960 22615 32963
rect 24688 32960 24716 33000
rect 25314 32988 25320 33000
rect 25372 32988 25378 33040
rect 22603 32932 24716 32960
rect 22603 32929 22615 32932
rect 22557 32923 22615 32929
rect 25038 32920 25044 32972
rect 25096 32920 25102 32972
rect 25222 32920 25228 32972
rect 25280 32920 25286 32972
rect 23658 32852 23664 32904
rect 23716 32852 23722 32904
rect 24946 32852 24952 32904
rect 25004 32892 25010 32904
rect 25406 32892 25412 32904
rect 25004 32864 25412 32892
rect 25004 32852 25010 32864
rect 25406 32852 25412 32864
rect 25464 32852 25470 32904
rect 24670 32784 24676 32836
rect 24728 32824 24734 32836
rect 24728 32796 24992 32824
rect 24728 32784 24734 32796
rect 23842 32756 23848 32768
rect 21928 32728 23848 32756
rect 23842 32716 23848 32728
rect 23900 32716 23906 32768
rect 24581 32759 24639 32765
rect 24581 32725 24593 32759
rect 24627 32756 24639 32759
rect 24854 32756 24860 32768
rect 24627 32728 24860 32756
rect 24627 32725 24639 32728
rect 24581 32719 24639 32725
rect 24854 32716 24860 32728
rect 24912 32716 24918 32768
rect 24964 32765 24992 32796
rect 24949 32759 25007 32765
rect 24949 32725 24961 32759
rect 24995 32725 25007 32759
rect 24949 32719 25007 32725
rect 1104 32666 25852 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 25852 32666
rect 1104 32592 25852 32614
rect 17034 32552 17040 32564
rect 16546 32524 17040 32552
rect 15378 32444 15384 32496
rect 15436 32484 15442 32496
rect 16546 32484 16574 32524
rect 17034 32512 17040 32524
rect 17092 32512 17098 32564
rect 23934 32552 23940 32564
rect 18616 32524 23940 32552
rect 15436 32456 16574 32484
rect 15436 32444 15442 32456
rect 16666 32444 16672 32496
rect 16724 32484 16730 32496
rect 16853 32487 16911 32493
rect 16853 32484 16865 32487
rect 16724 32456 16865 32484
rect 16724 32444 16730 32456
rect 16853 32453 16865 32456
rect 16899 32484 16911 32487
rect 18616 32484 18644 32524
rect 23934 32512 23940 32524
rect 23992 32512 23998 32564
rect 25225 32555 25283 32561
rect 25225 32521 25237 32555
rect 25271 32552 25283 32555
rect 25314 32552 25320 32564
rect 25271 32524 25320 32552
rect 25271 32521 25283 32524
rect 25225 32515 25283 32521
rect 25314 32512 25320 32524
rect 25372 32552 25378 32564
rect 26050 32552 26056 32564
rect 25372 32524 26056 32552
rect 25372 32512 25378 32524
rect 26050 32512 26056 32524
rect 26108 32512 26114 32564
rect 16899 32456 18644 32484
rect 16899 32453 16911 32456
rect 16853 32447 16911 32453
rect 22278 32444 22284 32496
rect 22336 32484 22342 32496
rect 22833 32487 22891 32493
rect 22833 32484 22845 32487
rect 22336 32456 22845 32484
rect 22336 32444 22342 32456
rect 22833 32453 22845 32456
rect 22879 32484 22891 32487
rect 22879 32456 23520 32484
rect 22879 32453 22891 32456
rect 22833 32447 22891 32453
rect 20470 32388 21312 32416
rect 13354 32308 13360 32360
rect 13412 32348 13418 32360
rect 16117 32351 16175 32357
rect 16117 32348 16129 32351
rect 13412 32320 16129 32348
rect 13412 32308 13418 32320
rect 16117 32317 16129 32320
rect 16163 32348 16175 32351
rect 16758 32348 16764 32360
rect 16163 32320 16764 32348
rect 16163 32317 16175 32320
rect 16117 32311 16175 32317
rect 16758 32308 16764 32320
rect 16816 32308 16822 32360
rect 19061 32351 19119 32357
rect 19061 32317 19073 32351
rect 19107 32317 19119 32351
rect 19061 32311 19119 32317
rect 19337 32351 19395 32357
rect 19337 32317 19349 32351
rect 19383 32348 19395 32351
rect 21174 32348 21180 32360
rect 19383 32320 21180 32348
rect 19383 32317 19395 32320
rect 19337 32311 19395 32317
rect 16574 32172 16580 32224
rect 16632 32212 16638 32224
rect 18966 32212 18972 32224
rect 16632 32184 18972 32212
rect 16632 32172 16638 32184
rect 18966 32172 18972 32184
rect 19024 32172 19030 32224
rect 19076 32212 19104 32311
rect 21174 32308 21180 32320
rect 21232 32308 21238 32360
rect 19426 32212 19432 32224
rect 19076 32184 19432 32212
rect 19426 32172 19432 32184
rect 19484 32172 19490 32224
rect 20809 32215 20867 32221
rect 20809 32181 20821 32215
rect 20855 32212 20867 32215
rect 20898 32212 20904 32224
rect 20855 32184 20904 32212
rect 20855 32181 20867 32184
rect 20809 32175 20867 32181
rect 20898 32172 20904 32184
rect 20956 32172 20962 32224
rect 21177 32215 21235 32221
rect 21177 32181 21189 32215
rect 21223 32212 21235 32215
rect 21284 32212 21312 32388
rect 21818 32376 21824 32428
rect 21876 32416 21882 32428
rect 23492 32425 23520 32456
rect 24762 32444 24768 32496
rect 24820 32444 24826 32496
rect 22097 32419 22155 32425
rect 22097 32416 22109 32419
rect 21876 32388 22109 32416
rect 21876 32376 21882 32388
rect 22097 32385 22109 32388
rect 22143 32385 22155 32419
rect 22097 32379 22155 32385
rect 23477 32419 23535 32425
rect 23477 32385 23489 32419
rect 23523 32385 23535 32419
rect 23477 32379 23535 32385
rect 23753 32351 23811 32357
rect 23753 32317 23765 32351
rect 23799 32348 23811 32351
rect 25222 32348 25228 32360
rect 23799 32320 25228 32348
rect 23799 32317 23811 32320
rect 23753 32311 23811 32317
rect 25222 32308 25228 32320
rect 25280 32308 25286 32360
rect 21450 32240 21456 32292
rect 21508 32280 21514 32292
rect 21508 32252 21956 32280
rect 21508 32240 21514 32252
rect 21358 32212 21364 32224
rect 21223 32184 21364 32212
rect 21223 32181 21235 32184
rect 21177 32175 21235 32181
rect 21358 32172 21364 32184
rect 21416 32172 21422 32224
rect 21637 32215 21695 32221
rect 21637 32181 21649 32215
rect 21683 32212 21695 32215
rect 21818 32212 21824 32224
rect 21683 32184 21824 32212
rect 21683 32181 21695 32184
rect 21637 32175 21695 32181
rect 21818 32172 21824 32184
rect 21876 32172 21882 32224
rect 21928 32212 21956 32252
rect 26510 32212 26516 32224
rect 21928 32184 26516 32212
rect 26510 32172 26516 32184
rect 26568 32172 26574 32224
rect 1104 32122 25852 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 25852 32122
rect 1104 32048 25852 32070
rect 17024 32011 17082 32017
rect 17024 31977 17036 32011
rect 17070 32008 17082 32011
rect 18506 32008 18512 32020
rect 17070 31980 18512 32008
rect 17070 31977 17082 31980
rect 17024 31971 17082 31977
rect 18506 31968 18512 31980
rect 18564 31968 18570 32020
rect 18966 31968 18972 32020
rect 19024 32008 19030 32020
rect 21450 32008 21456 32020
rect 19024 31980 21456 32008
rect 19024 31968 19030 31980
rect 21450 31968 21456 31980
rect 21508 31968 21514 32020
rect 22186 31968 22192 32020
rect 22244 32008 22250 32020
rect 22649 32011 22707 32017
rect 22649 32008 22661 32011
rect 22244 31980 22661 32008
rect 22244 31968 22250 31980
rect 22649 31977 22661 31980
rect 22695 31977 22707 32011
rect 22649 31971 22707 31977
rect 12526 31900 12532 31952
rect 12584 31940 12590 31952
rect 15565 31943 15623 31949
rect 15565 31940 15577 31943
rect 12584 31912 15577 31940
rect 12584 31900 12590 31912
rect 15565 31909 15577 31912
rect 15611 31909 15623 31943
rect 15565 31903 15623 31909
rect 20732 31912 22232 31940
rect 16114 31832 16120 31884
rect 16172 31832 16178 31884
rect 17678 31832 17684 31884
rect 17736 31872 17742 31884
rect 18509 31875 18567 31881
rect 18509 31872 18521 31875
rect 17736 31844 18521 31872
rect 17736 31832 17742 31844
rect 18509 31841 18521 31844
rect 18555 31841 18567 31875
rect 18509 31835 18567 31841
rect 19702 31832 19708 31884
rect 19760 31872 19766 31884
rect 20732 31872 20760 31912
rect 19760 31844 20760 31872
rect 19760 31832 19766 31844
rect 21910 31832 21916 31884
rect 21968 31872 21974 31884
rect 22204 31881 22232 31912
rect 22097 31875 22155 31881
rect 22097 31872 22109 31875
rect 21968 31844 22109 31872
rect 21968 31832 21974 31844
rect 22097 31841 22109 31844
rect 22143 31841 22155 31875
rect 22097 31835 22155 31841
rect 22189 31875 22247 31881
rect 22189 31841 22201 31875
rect 22235 31841 22247 31875
rect 22189 31835 22247 31841
rect 16025 31807 16083 31813
rect 16025 31773 16037 31807
rect 16071 31804 16083 31807
rect 16574 31804 16580 31816
rect 16071 31776 16580 31804
rect 16071 31773 16083 31776
rect 16025 31767 16083 31773
rect 16574 31764 16580 31776
rect 16632 31764 16638 31816
rect 16758 31764 16764 31816
rect 16816 31764 16822 31816
rect 19426 31764 19432 31816
rect 19484 31764 19490 31816
rect 21358 31736 21364 31748
rect 18262 31708 18920 31736
rect 20930 31708 21364 31736
rect 15933 31671 15991 31677
rect 15933 31637 15945 31671
rect 15979 31668 15991 31671
rect 16666 31668 16672 31680
rect 15979 31640 16672 31668
rect 15979 31637 15991 31640
rect 15933 31631 15991 31637
rect 16666 31628 16672 31640
rect 16724 31628 16730 31680
rect 18892 31677 18920 31708
rect 21358 31696 21364 31708
rect 21416 31696 21422 31748
rect 22554 31736 22560 31748
rect 22066 31708 22560 31736
rect 22066 31680 22094 31708
rect 22554 31696 22560 31708
rect 22612 31696 22618 31748
rect 22664 31736 22692 31971
rect 22738 31900 22744 31952
rect 22796 31940 22802 31952
rect 23017 31943 23075 31949
rect 23017 31940 23029 31943
rect 22796 31912 23029 31940
rect 22796 31900 22802 31912
rect 23017 31909 23029 31912
rect 23063 31909 23075 31943
rect 23017 31903 23075 31909
rect 25038 31900 25044 31952
rect 25096 31940 25102 31952
rect 25133 31943 25191 31949
rect 25133 31940 25145 31943
rect 25096 31912 25145 31940
rect 25096 31900 25102 31912
rect 25133 31909 25145 31912
rect 25179 31909 25191 31943
rect 25133 31903 25191 31909
rect 23290 31832 23296 31884
rect 23348 31872 23354 31884
rect 23477 31875 23535 31881
rect 23477 31872 23489 31875
rect 23348 31844 23489 31872
rect 23348 31832 23354 31844
rect 23477 31841 23489 31844
rect 23523 31841 23535 31875
rect 23477 31835 23535 31841
rect 23569 31875 23627 31881
rect 23569 31841 23581 31875
rect 23615 31841 23627 31875
rect 23569 31835 23627 31841
rect 23014 31764 23020 31816
rect 23072 31804 23078 31816
rect 23584 31804 23612 31835
rect 23072 31776 23612 31804
rect 24857 31807 24915 31813
rect 23072 31764 23078 31776
rect 24857 31773 24869 31807
rect 24903 31804 24915 31807
rect 25314 31804 25320 31816
rect 24903 31776 25320 31804
rect 24903 31773 24915 31776
rect 24857 31767 24915 31773
rect 25314 31764 25320 31776
rect 25372 31764 25378 31816
rect 23385 31739 23443 31745
rect 23385 31736 23397 31739
rect 22664 31708 23397 31736
rect 23385 31705 23397 31708
rect 23431 31705 23443 31739
rect 23385 31699 23443 31705
rect 18877 31671 18935 31677
rect 18877 31637 18889 31671
rect 18923 31668 18935 31671
rect 18966 31668 18972 31680
rect 18923 31640 18972 31668
rect 18923 31637 18935 31640
rect 18877 31631 18935 31637
rect 18966 31628 18972 31640
rect 19024 31628 19030 31680
rect 20990 31628 20996 31680
rect 21048 31668 21054 31680
rect 21177 31671 21235 31677
rect 21177 31668 21189 31671
rect 21048 31640 21189 31668
rect 21048 31628 21054 31640
rect 21177 31637 21189 31640
rect 21223 31637 21235 31671
rect 21177 31631 21235 31637
rect 21634 31628 21640 31680
rect 21692 31628 21698 31680
rect 22002 31628 22008 31680
rect 22060 31640 22094 31680
rect 24673 31671 24731 31677
rect 22060 31628 22066 31640
rect 24673 31637 24685 31671
rect 24719 31668 24731 31671
rect 24762 31668 24768 31680
rect 24719 31640 24768 31668
rect 24719 31637 24731 31640
rect 24673 31631 24731 31637
rect 24762 31628 24768 31640
rect 24820 31628 24826 31680
rect 1104 31578 25852 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 25852 31578
rect 1104 31504 25852 31526
rect 15749 31467 15807 31473
rect 15749 31464 15761 31467
rect 14936 31436 15761 31464
rect 14936 31408 14964 31436
rect 15749 31433 15761 31436
rect 15795 31464 15807 31467
rect 19153 31467 19211 31473
rect 15795 31436 19012 31464
rect 15795 31433 15807 31436
rect 15749 31427 15807 31433
rect 18984 31408 19012 31436
rect 19153 31433 19165 31467
rect 19199 31464 19211 31467
rect 19702 31464 19708 31476
rect 19199 31436 19708 31464
rect 19199 31433 19211 31436
rect 19153 31427 19211 31433
rect 19702 31424 19708 31436
rect 19760 31424 19766 31476
rect 21358 31424 21364 31476
rect 21416 31424 21422 31476
rect 21545 31467 21603 31473
rect 21545 31433 21557 31467
rect 21591 31464 21603 31467
rect 21726 31464 21732 31476
rect 21591 31436 21732 31464
rect 21591 31433 21603 31436
rect 21545 31427 21603 31433
rect 21726 31424 21732 31436
rect 21784 31464 21790 31476
rect 22002 31464 22008 31476
rect 21784 31436 22008 31464
rect 21784 31424 21790 31436
rect 22002 31424 22008 31436
rect 22060 31424 22066 31476
rect 23566 31424 23572 31476
rect 23624 31464 23630 31476
rect 24213 31467 24271 31473
rect 24213 31464 24225 31467
rect 23624 31436 24225 31464
rect 23624 31424 23630 31436
rect 24213 31433 24225 31436
rect 24259 31433 24271 31467
rect 24213 31427 24271 31433
rect 25498 31424 25504 31476
rect 25556 31424 25562 31476
rect 14918 31396 14924 31408
rect 14858 31368 14924 31396
rect 14918 31356 14924 31368
rect 14976 31356 14982 31408
rect 18966 31396 18972 31408
rect 18906 31368 18972 31396
rect 18966 31356 18972 31368
rect 19024 31396 19030 31408
rect 19521 31399 19579 31405
rect 19521 31396 19533 31399
rect 19024 31368 19533 31396
rect 19024 31356 19030 31368
rect 19521 31365 19533 31368
rect 19567 31396 19579 31399
rect 21376 31396 21404 31424
rect 19567 31368 21404 31396
rect 19567 31365 19579 31368
rect 19521 31359 19579 31365
rect 22646 31356 22652 31408
rect 22704 31396 22710 31408
rect 22741 31399 22799 31405
rect 22741 31396 22753 31399
rect 22704 31368 22753 31396
rect 22704 31356 22710 31368
rect 22741 31365 22753 31368
rect 22787 31396 22799 31399
rect 23014 31396 23020 31408
rect 22787 31368 23020 31396
rect 22787 31365 22799 31368
rect 22741 31359 22799 31365
rect 23014 31356 23020 31368
rect 23072 31356 23078 31408
rect 25516 31396 25544 31424
rect 24044 31368 25544 31396
rect 16758 31288 16764 31340
rect 16816 31328 16822 31340
rect 17405 31331 17463 31337
rect 17405 31328 17417 31331
rect 16816 31300 17417 31328
rect 16816 31288 16822 31300
rect 17405 31297 17417 31300
rect 17451 31297 17463 31331
rect 17405 31291 17463 31297
rect 20438 31288 20444 31340
rect 20496 31288 20502 31340
rect 20533 31331 20591 31337
rect 20533 31297 20545 31331
rect 20579 31328 20591 31331
rect 20579 31300 22232 31328
rect 20579 31297 20591 31300
rect 20533 31291 20591 31297
rect 13354 31220 13360 31272
rect 13412 31220 13418 31272
rect 13633 31263 13691 31269
rect 13633 31229 13645 31263
rect 13679 31260 13691 31263
rect 15473 31263 15531 31269
rect 15473 31260 15485 31263
rect 13679 31232 15485 31260
rect 13679 31229 13691 31232
rect 13633 31223 13691 31229
rect 15473 31229 15485 31232
rect 15519 31260 15531 31263
rect 16114 31260 16120 31272
rect 15519 31232 16120 31260
rect 15519 31229 15531 31232
rect 15473 31223 15531 31229
rect 16114 31220 16120 31232
rect 16172 31260 16178 31272
rect 16393 31263 16451 31269
rect 16393 31260 16405 31263
rect 16172 31232 16405 31260
rect 16172 31220 16178 31232
rect 16393 31229 16405 31232
rect 16439 31229 16451 31263
rect 16393 31223 16451 31229
rect 17678 31220 17684 31272
rect 17736 31220 17742 31272
rect 18690 31220 18696 31272
rect 18748 31260 18754 31272
rect 20625 31263 20683 31269
rect 20625 31260 20637 31263
rect 18748 31232 20637 31260
rect 18748 31220 18754 31232
rect 20625 31229 20637 31232
rect 20671 31229 20683 31263
rect 22204 31260 22232 31300
rect 22278 31288 22284 31340
rect 22336 31328 22342 31340
rect 22465 31331 22523 31337
rect 22465 31328 22477 31331
rect 22336 31300 22477 31328
rect 22336 31288 22342 31300
rect 22465 31297 22477 31300
rect 22511 31297 22523 31331
rect 22465 31291 22523 31297
rect 23842 31288 23848 31340
rect 23900 31288 23906 31340
rect 24044 31260 24072 31368
rect 25317 31331 25375 31337
rect 25317 31297 25329 31331
rect 25363 31328 25375 31331
rect 25498 31328 25504 31340
rect 25363 31300 25504 31328
rect 25363 31297 25375 31300
rect 25317 31291 25375 31297
rect 25498 31288 25504 31300
rect 25556 31288 25562 31340
rect 22204 31232 24072 31260
rect 20625 31223 20683 31229
rect 25130 31220 25136 31272
rect 25188 31260 25194 31272
rect 25866 31260 25872 31272
rect 25188 31232 25872 31260
rect 25188 31220 25194 31232
rect 25866 31220 25872 31232
rect 25924 31220 25930 31272
rect 20073 31195 20131 31201
rect 20073 31192 20085 31195
rect 18708 31164 20085 31192
rect 13814 31084 13820 31136
rect 13872 31124 13878 31136
rect 15105 31127 15163 31133
rect 15105 31124 15117 31127
rect 13872 31096 15117 31124
rect 13872 31084 13878 31096
rect 15105 31093 15117 31096
rect 15151 31093 15163 31127
rect 15105 31087 15163 31093
rect 16574 31084 16580 31136
rect 16632 31124 16638 31136
rect 16758 31124 16764 31136
rect 16632 31096 16764 31124
rect 16632 31084 16638 31096
rect 16758 31084 16764 31096
rect 16816 31084 16822 31136
rect 17494 31084 17500 31136
rect 17552 31124 17558 31136
rect 18708 31124 18736 31164
rect 20073 31161 20085 31164
rect 20119 31161 20131 31195
rect 20073 31155 20131 31161
rect 17552 31096 18736 31124
rect 19797 31127 19855 31133
rect 17552 31084 17558 31096
rect 19797 31093 19809 31127
rect 19843 31124 19855 31127
rect 20438 31124 20444 31136
rect 19843 31096 20444 31124
rect 19843 31093 19855 31096
rect 19797 31087 19855 31093
rect 20438 31084 20444 31096
rect 20496 31124 20502 31136
rect 21174 31124 21180 31136
rect 20496 31096 21180 31124
rect 20496 31084 20502 31096
rect 21174 31084 21180 31096
rect 21232 31084 21238 31136
rect 23842 31084 23848 31136
rect 23900 31124 23906 31136
rect 24581 31127 24639 31133
rect 24581 31124 24593 31127
rect 23900 31096 24593 31124
rect 23900 31084 23906 31096
rect 24581 31093 24593 31096
rect 24627 31124 24639 31127
rect 24762 31124 24768 31136
rect 24627 31096 24768 31124
rect 24627 31093 24639 31096
rect 24581 31087 24639 31093
rect 24762 31084 24768 31096
rect 24820 31084 24826 31136
rect 25130 31084 25136 31136
rect 25188 31084 25194 31136
rect 1104 31034 25852 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 25852 31034
rect 1104 30960 25852 30982
rect 9125 30923 9183 30929
rect 9125 30889 9137 30923
rect 9171 30920 9183 30923
rect 10226 30920 10232 30932
rect 9171 30892 10232 30920
rect 9171 30889 9183 30892
rect 9125 30883 9183 30889
rect 10226 30880 10232 30892
rect 10284 30880 10290 30932
rect 15378 30880 15384 30932
rect 15436 30920 15442 30932
rect 15565 30923 15623 30929
rect 15565 30920 15577 30923
rect 15436 30892 15577 30920
rect 15436 30880 15442 30892
rect 15565 30889 15577 30892
rect 15611 30920 15623 30923
rect 15749 30923 15807 30929
rect 15749 30920 15761 30923
rect 15611 30892 15761 30920
rect 15611 30889 15623 30892
rect 15565 30883 15623 30889
rect 15749 30889 15761 30892
rect 15795 30889 15807 30923
rect 15749 30883 15807 30889
rect 18509 30923 18567 30929
rect 18509 30889 18521 30923
rect 18555 30920 18567 30923
rect 18690 30920 18696 30932
rect 18555 30892 18696 30920
rect 18555 30889 18567 30892
rect 18509 30883 18567 30889
rect 18690 30880 18696 30892
rect 18748 30880 18754 30932
rect 18877 30923 18935 30929
rect 18877 30889 18889 30923
rect 18923 30920 18935 30923
rect 18966 30920 18972 30932
rect 18923 30892 18972 30920
rect 18923 30889 18935 30892
rect 18877 30883 18935 30889
rect 18966 30880 18972 30892
rect 19024 30880 19030 30932
rect 22465 30923 22523 30929
rect 22465 30889 22477 30923
rect 22511 30920 22523 30923
rect 22646 30920 22652 30932
rect 22511 30892 22652 30920
rect 22511 30889 22523 30892
rect 22465 30883 22523 30889
rect 22646 30880 22652 30892
rect 22704 30880 22710 30932
rect 22833 30923 22891 30929
rect 22833 30889 22845 30923
rect 22879 30920 22891 30923
rect 23842 30920 23848 30932
rect 22879 30892 23848 30920
rect 22879 30889 22891 30892
rect 22833 30883 22891 30889
rect 16761 30787 16819 30793
rect 16761 30753 16773 30787
rect 16807 30784 16819 30787
rect 19426 30784 19432 30796
rect 16807 30756 19432 30784
rect 16807 30753 16819 30756
rect 16761 30747 16819 30753
rect 19426 30744 19432 30756
rect 19484 30784 19490 30796
rect 20717 30787 20775 30793
rect 20717 30784 20729 30787
rect 19484 30756 20729 30784
rect 19484 30744 19490 30756
rect 20717 30753 20729 30756
rect 20763 30753 20775 30787
rect 20717 30747 20775 30753
rect 21358 30744 21364 30796
rect 21416 30784 21422 30796
rect 21416 30756 22140 30784
rect 21416 30744 21422 30756
rect 8754 30676 8760 30728
rect 8812 30716 8818 30728
rect 9309 30719 9367 30725
rect 9309 30716 9321 30719
rect 8812 30688 9321 30716
rect 8812 30676 8818 30688
rect 9309 30685 9321 30688
rect 9355 30685 9367 30719
rect 9309 30679 9367 30685
rect 14090 30676 14096 30728
rect 14148 30716 14154 30728
rect 14369 30719 14427 30725
rect 14369 30716 14381 30719
rect 14148 30688 14381 30716
rect 14148 30676 14154 30688
rect 14369 30685 14381 30688
rect 14415 30716 14427 30719
rect 15378 30716 15384 30728
rect 14415 30688 15384 30716
rect 14415 30685 14427 30688
rect 14369 30679 14427 30685
rect 15378 30676 15384 30688
rect 15436 30676 15442 30728
rect 22112 30716 22140 30756
rect 22848 30716 22876 30883
rect 23842 30880 23848 30892
rect 23900 30880 23906 30932
rect 25498 30880 25504 30932
rect 25556 30880 25562 30932
rect 22112 30702 22876 30716
rect 22126 30688 22876 30702
rect 15102 30608 15108 30660
rect 15160 30608 15166 30660
rect 17037 30651 17095 30657
rect 17037 30617 17049 30651
rect 17083 30617 17095 30651
rect 18966 30648 18972 30660
rect 18262 30620 18972 30648
rect 17037 30611 17095 30617
rect 17052 30580 17080 30611
rect 18966 30608 18972 30620
rect 19024 30608 19030 30660
rect 20990 30608 20996 30660
rect 21048 30608 21054 30660
rect 22646 30608 22652 30660
rect 22704 30648 22710 30660
rect 24581 30651 24639 30657
rect 24581 30648 24593 30651
rect 22704 30620 24593 30648
rect 22704 30608 22710 30620
rect 24581 30617 24593 30620
rect 24627 30617 24639 30651
rect 24581 30611 24639 30617
rect 18782 30580 18788 30592
rect 17052 30552 18788 30580
rect 18782 30540 18788 30552
rect 18840 30540 18846 30592
rect 20070 30540 20076 30592
rect 20128 30540 20134 30592
rect 1104 30490 25852 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 25852 30490
rect 1104 30416 25852 30438
rect 13354 30376 13360 30388
rect 12406 30348 13360 30376
rect 12406 30308 12434 30348
rect 13354 30336 13360 30348
rect 13412 30336 13418 30388
rect 15933 30379 15991 30385
rect 15933 30345 15945 30379
rect 15979 30376 15991 30379
rect 16574 30376 16580 30388
rect 15979 30348 16580 30376
rect 15979 30345 15991 30348
rect 15933 30339 15991 30345
rect 16574 30336 16580 30348
rect 16632 30376 16638 30388
rect 16761 30379 16819 30385
rect 16761 30376 16773 30379
rect 16632 30348 16773 30376
rect 16632 30336 16638 30348
rect 16761 30345 16773 30348
rect 16807 30376 16819 30379
rect 16807 30348 18184 30376
rect 16807 30345 16819 30348
rect 16761 30339 16819 30345
rect 11808 30280 12434 30308
rect 7650 30200 7656 30252
rect 7708 30240 7714 30252
rect 11808 30249 11836 30280
rect 12710 30268 12716 30320
rect 12768 30268 12774 30320
rect 14090 30268 14096 30320
rect 14148 30268 14154 30320
rect 14550 30268 14556 30320
rect 14608 30308 14614 30320
rect 14608 30280 18092 30308
rect 14608 30268 14614 30280
rect 9125 30243 9183 30249
rect 9125 30240 9137 30243
rect 7708 30212 9137 30240
rect 7708 30200 7714 30212
rect 9125 30209 9137 30212
rect 9171 30209 9183 30243
rect 9125 30203 9183 30209
rect 11793 30243 11851 30249
rect 11793 30209 11805 30243
rect 11839 30209 11851 30243
rect 11793 30203 11851 30209
rect 15841 30243 15899 30249
rect 15841 30209 15853 30243
rect 15887 30240 15899 30243
rect 16850 30240 16856 30252
rect 15887 30212 16856 30240
rect 15887 30209 15899 30212
rect 15841 30203 15899 30209
rect 16850 30200 16856 30212
rect 16908 30200 16914 30252
rect 12066 30132 12072 30184
rect 12124 30132 12130 30184
rect 12158 30132 12164 30184
rect 12216 30172 12222 30184
rect 12710 30172 12716 30184
rect 12216 30144 12716 30172
rect 12216 30132 12222 30144
rect 12710 30132 12716 30144
rect 12768 30132 12774 30184
rect 13354 30132 13360 30184
rect 13412 30172 13418 30184
rect 14829 30175 14887 30181
rect 14829 30172 14841 30175
rect 13412 30144 14841 30172
rect 13412 30132 13418 30144
rect 14829 30141 14841 30144
rect 14875 30141 14887 30175
rect 14829 30135 14887 30141
rect 16022 30132 16028 30184
rect 16080 30132 16086 30184
rect 18064 30172 18092 30280
rect 18156 30240 18184 30348
rect 18966 30336 18972 30388
rect 19024 30336 19030 30388
rect 20070 30336 20076 30388
rect 20128 30376 20134 30388
rect 20257 30379 20315 30385
rect 20257 30376 20269 30379
rect 20128 30348 20269 30376
rect 20128 30336 20134 30348
rect 20257 30345 20269 30348
rect 20303 30345 20315 30379
rect 20257 30339 20315 30345
rect 18322 30268 18328 30320
rect 18380 30308 18386 30320
rect 18984 30308 19012 30336
rect 18380 30280 19012 30308
rect 20349 30311 20407 30317
rect 18380 30268 18386 30280
rect 20349 30277 20361 30311
rect 20395 30308 20407 30311
rect 21910 30308 21916 30320
rect 20395 30280 21916 30308
rect 20395 30277 20407 30280
rect 20349 30271 20407 30277
rect 21910 30268 21916 30280
rect 21968 30268 21974 30320
rect 22462 30268 22468 30320
rect 22520 30268 22526 30320
rect 22830 30268 22836 30320
rect 22888 30268 22894 30320
rect 24854 30308 24860 30320
rect 24794 30280 24860 30308
rect 24854 30268 24860 30280
rect 24912 30268 24918 30320
rect 21269 30243 21327 30249
rect 18156 30212 20668 30240
rect 19978 30172 19984 30184
rect 18064 30144 19984 30172
rect 19978 30132 19984 30144
rect 20036 30132 20042 30184
rect 20530 30132 20536 30184
rect 20588 30132 20594 30184
rect 20640 30172 20668 30212
rect 21269 30209 21281 30243
rect 21315 30240 21327 30243
rect 22373 30243 22431 30249
rect 22373 30240 22385 30243
rect 21315 30212 22385 30240
rect 21315 30209 21327 30212
rect 21269 30203 21327 30209
rect 22373 30209 22385 30212
rect 22419 30209 22431 30243
rect 22848 30240 22876 30268
rect 22373 30203 22431 30209
rect 22664 30212 22876 30240
rect 22664 30181 22692 30212
rect 22649 30175 22707 30181
rect 20640 30144 22232 30172
rect 8938 30064 8944 30116
rect 8996 30064 9002 30116
rect 16482 30064 16488 30116
rect 16540 30104 16546 30116
rect 22094 30104 22100 30116
rect 16540 30076 22100 30104
rect 16540 30064 16546 30076
rect 22094 30064 22100 30076
rect 22152 30064 22158 30116
rect 11514 29996 11520 30048
rect 11572 30036 11578 30048
rect 13541 30039 13599 30045
rect 13541 30036 13553 30039
rect 11572 30008 13553 30036
rect 11572 29996 11578 30008
rect 13541 30005 13553 30008
rect 13587 30036 13599 30039
rect 13630 30036 13636 30048
rect 13587 30008 13636 30036
rect 13587 30005 13599 30008
rect 13541 29999 13599 30005
rect 13630 29996 13636 30008
rect 13688 29996 13694 30048
rect 15473 30039 15531 30045
rect 15473 30005 15485 30039
rect 15519 30036 15531 30039
rect 15930 30036 15936 30048
rect 15519 30008 15936 30036
rect 15519 30005 15531 30008
rect 15473 29999 15531 30005
rect 15930 29996 15936 30008
rect 15988 29996 15994 30048
rect 19794 29996 19800 30048
rect 19852 30036 19858 30048
rect 19889 30039 19947 30045
rect 19889 30036 19901 30039
rect 19852 30008 19901 30036
rect 19852 29996 19858 30008
rect 19889 30005 19901 30008
rect 19935 30005 19947 30039
rect 19889 29999 19947 30005
rect 21910 29996 21916 30048
rect 21968 30036 21974 30048
rect 22005 30039 22063 30045
rect 22005 30036 22017 30039
rect 21968 30008 22017 30036
rect 21968 29996 21974 30008
rect 22005 30005 22017 30008
rect 22051 30005 22063 30039
rect 22204 30036 22232 30144
rect 22649 30141 22661 30175
rect 22695 30141 22707 30175
rect 22649 30135 22707 30141
rect 22830 30132 22836 30184
rect 22888 30172 22894 30184
rect 23293 30175 23351 30181
rect 23293 30172 23305 30175
rect 22888 30144 23305 30172
rect 22888 30132 22894 30144
rect 23293 30141 23305 30144
rect 23339 30141 23351 30175
rect 23293 30135 23351 30141
rect 23566 30132 23572 30184
rect 23624 30132 23630 30184
rect 25041 30175 25099 30181
rect 25041 30141 25053 30175
rect 25087 30172 25099 30175
rect 25222 30172 25228 30184
rect 25087 30144 25228 30172
rect 25087 30141 25099 30144
rect 25041 30135 25099 30141
rect 25222 30132 25228 30144
rect 25280 30132 25286 30184
rect 26142 30104 26148 30116
rect 24596 30076 26148 30104
rect 24596 30036 24624 30076
rect 26142 30064 26148 30076
rect 26200 30064 26206 30116
rect 22204 30008 24624 30036
rect 22005 29999 22063 30005
rect 24854 29996 24860 30048
rect 24912 30036 24918 30048
rect 25222 30036 25228 30048
rect 24912 30008 25228 30036
rect 24912 29996 24918 30008
rect 25222 29996 25228 30008
rect 25280 30036 25286 30048
rect 25317 30039 25375 30045
rect 25317 30036 25329 30039
rect 25280 30008 25329 30036
rect 25280 29996 25286 30008
rect 25317 30005 25329 30008
rect 25363 30005 25375 30039
rect 25317 29999 25375 30005
rect 1104 29946 25852 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 25852 29946
rect 1104 29872 25852 29894
rect 12066 29792 12072 29844
rect 12124 29832 12130 29844
rect 13449 29835 13507 29841
rect 12124 29804 12940 29832
rect 12124 29792 12130 29804
rect 12912 29773 12940 29804
rect 13449 29801 13461 29835
rect 13495 29832 13507 29835
rect 13814 29832 13820 29844
rect 13495 29804 13820 29832
rect 13495 29801 13507 29804
rect 13449 29795 13507 29801
rect 13814 29792 13820 29804
rect 13872 29792 13878 29844
rect 16301 29835 16359 29841
rect 16301 29801 16313 29835
rect 16347 29832 16359 29835
rect 23845 29835 23903 29841
rect 16347 29804 22094 29832
rect 16347 29801 16359 29804
rect 16301 29795 16359 29801
rect 12897 29767 12955 29773
rect 12897 29733 12909 29767
rect 12943 29764 12955 29767
rect 12943 29736 15884 29764
rect 12943 29733 12955 29736
rect 12897 29727 12955 29733
rect 11149 29699 11207 29705
rect 11149 29665 11161 29699
rect 11195 29696 11207 29699
rect 11422 29696 11428 29708
rect 11195 29668 11428 29696
rect 11195 29665 11207 29668
rect 11149 29659 11207 29665
rect 11422 29656 11428 29668
rect 11480 29696 11486 29708
rect 13354 29696 13360 29708
rect 11480 29668 13360 29696
rect 11480 29656 11486 29668
rect 13354 29656 13360 29668
rect 13412 29656 13418 29708
rect 15856 29705 15884 29736
rect 15841 29699 15899 29705
rect 15841 29665 15853 29699
rect 15887 29696 15899 29699
rect 16022 29696 16028 29708
rect 15887 29668 16028 29696
rect 15887 29665 15899 29668
rect 15841 29659 15899 29665
rect 16022 29656 16028 29668
rect 16080 29656 16086 29708
rect 15565 29631 15623 29637
rect 15565 29597 15577 29631
rect 15611 29628 15623 29631
rect 15654 29628 15660 29640
rect 15611 29600 15660 29628
rect 15611 29597 15623 29600
rect 15565 29591 15623 29597
rect 15654 29588 15660 29600
rect 15712 29628 15718 29640
rect 16316 29628 16344 29795
rect 16482 29724 16488 29776
rect 16540 29724 16546 29776
rect 18414 29724 18420 29776
rect 18472 29764 18478 29776
rect 20165 29767 20223 29773
rect 20165 29764 20177 29767
rect 18472 29736 20177 29764
rect 18472 29724 18478 29736
rect 20165 29733 20177 29736
rect 20211 29733 20223 29767
rect 20165 29727 20223 29733
rect 17037 29699 17095 29705
rect 17037 29665 17049 29699
rect 17083 29696 17095 29699
rect 19334 29696 19340 29708
rect 17083 29668 19340 29696
rect 17083 29665 17095 29668
rect 17037 29659 17095 29665
rect 19334 29656 19340 29668
rect 19392 29656 19398 29708
rect 20717 29699 20775 29705
rect 20717 29696 20729 29699
rect 19444 29668 20729 29696
rect 18874 29628 18880 29640
rect 15712 29600 16344 29628
rect 18616 29600 18880 29628
rect 15712 29588 15718 29600
rect 11330 29520 11336 29572
rect 11388 29560 11394 29572
rect 11425 29563 11483 29569
rect 11425 29560 11437 29563
rect 11388 29532 11437 29560
rect 11388 29520 11394 29532
rect 11425 29529 11437 29532
rect 11471 29529 11483 29563
rect 12710 29560 12716 29572
rect 12650 29532 12716 29560
rect 11425 29523 11483 29529
rect 12710 29520 12716 29532
rect 12768 29520 12774 29572
rect 17313 29563 17371 29569
rect 17313 29529 17325 29563
rect 17359 29529 17371 29563
rect 17313 29523 17371 29529
rect 12728 29492 12756 29520
rect 13265 29495 13323 29501
rect 13265 29492 13277 29495
rect 12728 29464 13277 29492
rect 13265 29461 13277 29464
rect 13311 29492 13323 29495
rect 13725 29495 13783 29501
rect 13725 29492 13737 29495
rect 13311 29464 13737 29492
rect 13311 29461 13323 29464
rect 13265 29455 13323 29461
rect 13725 29461 13737 29464
rect 13771 29492 13783 29495
rect 14918 29492 14924 29504
rect 13771 29464 14924 29492
rect 13771 29461 13783 29464
rect 13725 29455 13783 29461
rect 14918 29452 14924 29464
rect 14976 29452 14982 29504
rect 15194 29452 15200 29504
rect 15252 29452 15258 29504
rect 15657 29495 15715 29501
rect 15657 29461 15669 29495
rect 15703 29492 15715 29495
rect 16114 29492 16120 29504
rect 15703 29464 16120 29492
rect 15703 29461 15715 29464
rect 15657 29455 15715 29461
rect 16114 29452 16120 29464
rect 16172 29492 16178 29504
rect 16482 29492 16488 29504
rect 16172 29464 16488 29492
rect 16172 29452 16178 29464
rect 16482 29452 16488 29464
rect 16540 29452 16546 29504
rect 17328 29492 17356 29523
rect 18322 29520 18328 29572
rect 18380 29520 18386 29572
rect 18616 29492 18644 29600
rect 18874 29588 18880 29600
rect 18932 29628 18938 29640
rect 19444 29628 19472 29668
rect 20717 29665 20729 29668
rect 20763 29665 20775 29699
rect 22066 29696 22094 29804
rect 23845 29801 23857 29835
rect 23891 29832 23903 29835
rect 26142 29832 26148 29844
rect 23891 29804 26148 29832
rect 23891 29801 23903 29804
rect 23845 29795 23903 29801
rect 26142 29792 26148 29804
rect 26200 29792 26206 29844
rect 23382 29724 23388 29776
rect 23440 29764 23446 29776
rect 25133 29767 25191 29773
rect 25133 29764 25145 29767
rect 23440 29736 25145 29764
rect 23440 29724 23446 29736
rect 25133 29733 25145 29736
rect 25179 29733 25191 29767
rect 25133 29727 25191 29733
rect 26602 29696 26608 29708
rect 22066 29668 26608 29696
rect 20717 29659 20775 29665
rect 26602 29656 26608 29668
rect 26660 29656 26666 29708
rect 18932 29600 19472 29628
rect 20625 29631 20683 29637
rect 18932 29588 18938 29600
rect 20625 29597 20637 29631
rect 20671 29628 20683 29631
rect 20806 29628 20812 29640
rect 20671 29600 20812 29628
rect 20671 29597 20683 29600
rect 20625 29591 20683 29597
rect 20806 29588 20812 29600
rect 20864 29588 20870 29640
rect 23385 29631 23443 29637
rect 23385 29597 23397 29631
rect 23431 29597 23443 29631
rect 23385 29591 23443 29597
rect 24029 29631 24087 29637
rect 24029 29597 24041 29631
rect 24075 29628 24087 29631
rect 24486 29628 24492 29640
rect 24075 29600 24492 29628
rect 24075 29597 24087 29600
rect 24029 29591 24087 29597
rect 22925 29563 22983 29569
rect 22925 29529 22937 29563
rect 22971 29560 22983 29563
rect 23400 29560 23428 29591
rect 24486 29588 24492 29600
rect 24544 29588 24550 29640
rect 25314 29588 25320 29640
rect 25372 29588 25378 29640
rect 24854 29560 24860 29572
rect 22971 29532 24860 29560
rect 22971 29529 22983 29532
rect 22925 29523 22983 29529
rect 24854 29520 24860 29532
rect 24912 29520 24918 29572
rect 17328 29464 18644 29492
rect 18782 29452 18788 29504
rect 18840 29452 18846 29504
rect 19150 29452 19156 29504
rect 19208 29492 19214 29504
rect 19429 29495 19487 29501
rect 19429 29492 19441 29495
rect 19208 29464 19441 29492
rect 19208 29452 19214 29464
rect 19429 29461 19441 29464
rect 19475 29461 19487 29495
rect 19429 29455 19487 29461
rect 19978 29452 19984 29504
rect 20036 29492 20042 29504
rect 20533 29495 20591 29501
rect 20533 29492 20545 29495
rect 20036 29464 20545 29492
rect 20036 29452 20042 29464
rect 20533 29461 20545 29464
rect 20579 29461 20591 29495
rect 20533 29455 20591 29461
rect 22462 29452 22468 29504
rect 22520 29492 22526 29504
rect 23201 29495 23259 29501
rect 23201 29492 23213 29495
rect 22520 29464 23213 29492
rect 22520 29452 22526 29464
rect 23201 29461 23213 29464
rect 23247 29461 23259 29495
rect 23201 29455 23259 29461
rect 24486 29452 24492 29504
rect 24544 29452 24550 29504
rect 24765 29495 24823 29501
rect 24765 29461 24777 29495
rect 24811 29492 24823 29495
rect 25222 29492 25228 29504
rect 24811 29464 25228 29492
rect 24811 29461 24823 29464
rect 24765 29455 24823 29461
rect 25222 29452 25228 29464
rect 25280 29452 25286 29504
rect 1104 29402 25852 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 25852 29402
rect 1104 29328 25852 29350
rect 8846 29248 8852 29300
rect 8904 29288 8910 29300
rect 9493 29291 9551 29297
rect 9493 29288 9505 29291
rect 8904 29260 9505 29288
rect 8904 29248 8910 29260
rect 9493 29257 9505 29260
rect 9539 29257 9551 29291
rect 9493 29251 9551 29257
rect 9861 29291 9919 29297
rect 9861 29257 9873 29291
rect 9907 29288 9919 29291
rect 10410 29288 10416 29300
rect 9907 29260 10416 29288
rect 9907 29257 9919 29260
rect 9861 29251 9919 29257
rect 10410 29248 10416 29260
rect 10468 29248 10474 29300
rect 12434 29248 12440 29300
rect 12492 29288 12498 29300
rect 12529 29291 12587 29297
rect 12529 29288 12541 29291
rect 12492 29260 12541 29288
rect 12492 29248 12498 29260
rect 12529 29257 12541 29260
rect 12575 29257 12587 29291
rect 12529 29251 12587 29257
rect 12618 29248 12624 29300
rect 12676 29248 12682 29300
rect 13814 29248 13820 29300
rect 13872 29248 13878 29300
rect 13906 29248 13912 29300
rect 13964 29288 13970 29300
rect 15105 29291 15163 29297
rect 15105 29288 15117 29291
rect 13964 29260 15117 29288
rect 13964 29248 13970 29260
rect 15105 29257 15117 29260
rect 15151 29257 15163 29291
rect 15105 29251 15163 29257
rect 9674 29180 9680 29232
rect 9732 29220 9738 29232
rect 13832 29220 13860 29248
rect 14918 29220 14924 29232
rect 9732 29192 10088 29220
rect 9732 29180 9738 29192
rect 10060 29093 10088 29192
rect 13280 29192 13860 29220
rect 14858 29192 14924 29220
rect 9953 29087 10011 29093
rect 9953 29053 9965 29087
rect 9999 29053 10011 29087
rect 9953 29047 10011 29053
rect 10045 29087 10103 29093
rect 10045 29053 10057 29087
rect 10091 29084 10103 29087
rect 10870 29084 10876 29096
rect 10091 29056 10876 29084
rect 10091 29053 10103 29056
rect 10045 29047 10103 29053
rect 9968 29016 9996 29047
rect 10870 29044 10876 29056
rect 10928 29044 10934 29096
rect 11790 29044 11796 29096
rect 11848 29084 11854 29096
rect 12805 29087 12863 29093
rect 12805 29084 12817 29087
rect 11848 29056 12817 29084
rect 11848 29044 11854 29056
rect 12805 29053 12817 29056
rect 12851 29084 12863 29087
rect 13280 29084 13308 29192
rect 14918 29180 14924 29192
rect 14976 29180 14982 29232
rect 13354 29112 13360 29164
rect 13412 29112 13418 29164
rect 15120 29152 15148 29251
rect 15194 29248 15200 29300
rect 15252 29288 15258 29300
rect 16025 29291 16083 29297
rect 16025 29288 16037 29291
rect 15252 29260 16037 29288
rect 15252 29248 15258 29260
rect 16025 29257 16037 29260
rect 16071 29257 16083 29291
rect 16025 29251 16083 29257
rect 17221 29291 17279 29297
rect 17221 29257 17233 29291
rect 17267 29288 17279 29291
rect 17494 29288 17500 29300
rect 17267 29260 17500 29288
rect 17267 29257 17279 29260
rect 17221 29251 17279 29257
rect 17494 29248 17500 29260
rect 17552 29288 17558 29300
rect 17862 29288 17868 29300
rect 17552 29260 17868 29288
rect 17552 29248 17558 29260
rect 17862 29248 17868 29260
rect 17920 29288 17926 29300
rect 18049 29291 18107 29297
rect 18049 29288 18061 29291
rect 17920 29260 18061 29288
rect 17920 29248 17926 29260
rect 18049 29257 18061 29260
rect 18095 29257 18107 29291
rect 18049 29251 18107 29257
rect 19150 29248 19156 29300
rect 19208 29248 19214 29300
rect 19245 29291 19303 29297
rect 19245 29257 19257 29291
rect 19291 29288 19303 29291
rect 20622 29288 20628 29300
rect 19291 29260 20628 29288
rect 19291 29257 19303 29260
rect 19245 29251 19303 29257
rect 20622 29248 20628 29260
rect 20680 29248 20686 29300
rect 23937 29291 23995 29297
rect 23937 29257 23949 29291
rect 23983 29288 23995 29291
rect 24118 29288 24124 29300
rect 23983 29260 24124 29288
rect 23983 29257 23995 29260
rect 23937 29251 23995 29257
rect 15930 29180 15936 29232
rect 15988 29180 15994 29232
rect 17034 29180 17040 29232
rect 17092 29220 17098 29232
rect 17313 29223 17371 29229
rect 17313 29220 17325 29223
rect 17092 29192 17325 29220
rect 17092 29180 17098 29192
rect 17313 29189 17325 29192
rect 17359 29220 17371 29223
rect 17957 29223 18015 29229
rect 17957 29220 17969 29223
rect 17359 29192 17969 29220
rect 17359 29189 17371 29192
rect 17313 29183 17371 29189
rect 17880 29164 17908 29192
rect 17957 29189 17969 29192
rect 18003 29189 18015 29223
rect 17957 29183 18015 29189
rect 19978 29180 19984 29232
rect 20036 29220 20042 29232
rect 20346 29220 20352 29232
rect 20036 29192 20352 29220
rect 20036 29180 20042 29192
rect 20346 29180 20352 29192
rect 20404 29220 20410 29232
rect 23952 29220 23980 29251
rect 24118 29248 24124 29260
rect 24176 29288 24182 29300
rect 24578 29288 24584 29300
rect 24176 29260 24584 29288
rect 24176 29248 24182 29260
rect 24578 29248 24584 29260
rect 24636 29248 24642 29300
rect 25314 29248 25320 29300
rect 25372 29288 25378 29300
rect 25409 29291 25467 29297
rect 25409 29288 25421 29291
rect 25372 29260 25421 29288
rect 25372 29248 25378 29260
rect 25409 29257 25421 29260
rect 25455 29257 25467 29291
rect 25409 29251 25467 29257
rect 20404 29192 23980 29220
rect 20404 29180 20410 29192
rect 17402 29152 17408 29164
rect 15120 29124 17408 29152
rect 17402 29112 17408 29124
rect 17460 29152 17466 29164
rect 17460 29124 17540 29152
rect 17460 29112 17466 29124
rect 12851 29056 13308 29084
rect 12851 29053 12863 29056
rect 12805 29047 12863 29053
rect 13630 29044 13636 29096
rect 13688 29084 13694 29096
rect 17512 29093 17540 29124
rect 17862 29112 17868 29164
rect 17920 29112 17926 29164
rect 22189 29155 22247 29161
rect 22189 29152 22201 29155
rect 22066 29124 22201 29152
rect 16117 29087 16175 29093
rect 16117 29084 16129 29087
rect 13688 29056 16129 29084
rect 13688 29044 13694 29056
rect 16117 29053 16129 29056
rect 16163 29053 16175 29087
rect 16117 29047 16175 29053
rect 17497 29087 17555 29093
rect 17497 29053 17509 29087
rect 17543 29053 17555 29087
rect 17497 29047 17555 29053
rect 19429 29087 19487 29093
rect 19429 29053 19441 29087
rect 19475 29084 19487 29087
rect 20898 29084 20904 29096
rect 19475 29056 20904 29084
rect 19475 29053 19487 29056
rect 19429 29047 19487 29053
rect 20898 29044 20904 29056
rect 20956 29044 20962 29096
rect 10226 29016 10232 29028
rect 9968 28988 10232 29016
rect 10226 28976 10232 28988
rect 10284 28976 10290 29028
rect 12158 28976 12164 29028
rect 12216 28976 12222 29028
rect 14642 28976 14648 29028
rect 14700 29016 14706 29028
rect 15565 29019 15623 29025
rect 15565 29016 15577 29019
rect 14700 28988 15577 29016
rect 14700 28976 14706 28988
rect 15565 28985 15577 28988
rect 15611 28985 15623 29019
rect 15565 28979 15623 28985
rect 15746 28976 15752 29028
rect 15804 29016 15810 29028
rect 16853 29019 16911 29025
rect 16853 29016 16865 29019
rect 15804 28988 16865 29016
rect 15804 28976 15810 28988
rect 16853 28985 16865 28988
rect 16899 28985 16911 29019
rect 18785 29019 18843 29025
rect 18785 29016 18797 29019
rect 16853 28979 16911 28985
rect 16960 28988 18797 29016
rect 13620 28951 13678 28957
rect 13620 28917 13632 28951
rect 13666 28948 13678 28951
rect 14090 28948 14096 28960
rect 13666 28920 14096 28948
rect 13666 28917 13678 28920
rect 13620 28911 13678 28917
rect 14090 28908 14096 28920
rect 14148 28908 14154 28960
rect 15286 28908 15292 28960
rect 15344 28948 15350 28960
rect 16960 28948 16988 28988
rect 18785 28985 18797 28988
rect 18831 28985 18843 29019
rect 18785 28979 18843 28985
rect 21818 28976 21824 29028
rect 21876 29016 21882 29028
rect 22066 29016 22094 29124
rect 22189 29121 22201 29124
rect 22235 29121 22247 29155
rect 22189 29115 22247 29121
rect 24029 29155 24087 29161
rect 24029 29121 24041 29155
rect 24075 29152 24087 29155
rect 25317 29155 25375 29161
rect 25317 29152 25329 29155
rect 24075 29124 25329 29152
rect 24075 29121 24087 29124
rect 24029 29115 24087 29121
rect 25317 29121 25329 29124
rect 25363 29152 25375 29155
rect 25406 29152 25412 29164
rect 25363 29124 25412 29152
rect 25363 29121 25375 29124
rect 25317 29115 25375 29121
rect 25406 29112 25412 29124
rect 25464 29112 25470 29164
rect 22830 29044 22836 29096
rect 22888 29084 22894 29096
rect 22925 29087 22983 29093
rect 22925 29084 22937 29087
rect 22888 29056 22937 29084
rect 22888 29044 22894 29056
rect 22925 29053 22937 29056
rect 22971 29053 22983 29087
rect 22925 29047 22983 29053
rect 23750 29044 23756 29096
rect 23808 29084 23814 29096
rect 24121 29087 24179 29093
rect 24121 29084 24133 29087
rect 23808 29056 24133 29084
rect 23808 29044 23814 29056
rect 24121 29053 24133 29056
rect 24167 29053 24179 29087
rect 24121 29047 24179 29053
rect 24765 29087 24823 29093
rect 24765 29053 24777 29087
rect 24811 29084 24823 29087
rect 24946 29084 24952 29096
rect 24811 29056 24952 29084
rect 24811 29053 24823 29056
rect 24765 29047 24823 29053
rect 24946 29044 24952 29056
rect 25004 29044 25010 29096
rect 21876 28988 22094 29016
rect 23569 29019 23627 29025
rect 21876 28976 21882 28988
rect 23569 28985 23581 29019
rect 23615 29016 23627 29019
rect 24670 29016 24676 29028
rect 23615 28988 24676 29016
rect 23615 28985 23627 28988
rect 23569 28979 23627 28985
rect 24670 28976 24676 28988
rect 24728 28976 24734 29028
rect 15344 28920 16988 28948
rect 15344 28908 15350 28920
rect 1104 28858 25852 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 25852 28858
rect 1104 28784 25852 28806
rect 10870 28704 10876 28756
rect 10928 28704 10934 28756
rect 13541 28747 13599 28753
rect 13541 28744 13553 28747
rect 12820 28716 13553 28744
rect 9125 28611 9183 28617
rect 9125 28577 9137 28611
rect 9171 28608 9183 28611
rect 11422 28608 11428 28620
rect 9171 28580 11428 28608
rect 9171 28577 9183 28580
rect 9125 28571 9183 28577
rect 11422 28568 11428 28580
rect 11480 28568 11486 28620
rect 11698 28568 11704 28620
rect 11756 28608 11762 28620
rect 12710 28608 12716 28620
rect 11756 28580 12716 28608
rect 11756 28568 11762 28580
rect 12710 28568 12716 28580
rect 12768 28608 12774 28620
rect 12820 28608 12848 28716
rect 13541 28713 13553 28716
rect 13587 28744 13599 28747
rect 13722 28744 13728 28756
rect 13587 28716 13728 28744
rect 13587 28713 13599 28716
rect 13541 28707 13599 28713
rect 13722 28704 13728 28716
rect 13780 28744 13786 28756
rect 14918 28744 14924 28756
rect 13780 28716 14924 28744
rect 13780 28704 13786 28716
rect 14918 28704 14924 28716
rect 14976 28744 14982 28756
rect 15841 28747 15899 28753
rect 15841 28744 15853 28747
rect 14976 28716 15853 28744
rect 14976 28704 14982 28716
rect 15841 28713 15853 28716
rect 15887 28713 15899 28747
rect 15841 28707 15899 28713
rect 18874 28704 18880 28756
rect 18932 28704 18938 28756
rect 22373 28747 22431 28753
rect 22373 28713 22385 28747
rect 22419 28744 22431 28747
rect 23750 28744 23756 28756
rect 22419 28716 23756 28744
rect 22419 28713 22431 28716
rect 22373 28707 22431 28713
rect 23750 28704 23756 28716
rect 23808 28704 23814 28756
rect 16482 28676 16488 28688
rect 15304 28648 16488 28676
rect 12768 28580 12848 28608
rect 12768 28568 12774 28580
rect 12820 28526 12848 28580
rect 13173 28611 13231 28617
rect 13173 28577 13185 28611
rect 13219 28608 13231 28611
rect 14090 28608 14096 28620
rect 13219 28580 14096 28608
rect 13219 28577 13231 28580
rect 13173 28571 13231 28577
rect 14090 28568 14096 28580
rect 14148 28568 14154 28620
rect 15304 28617 15332 28648
rect 16482 28636 16488 28648
rect 16540 28636 16546 28688
rect 22833 28679 22891 28685
rect 22833 28676 22845 28679
rect 22066 28648 22845 28676
rect 15289 28611 15347 28617
rect 15289 28577 15301 28611
rect 15335 28577 15347 28611
rect 15289 28571 15347 28577
rect 15378 28568 15384 28620
rect 15436 28568 15442 28620
rect 17405 28611 17463 28617
rect 17405 28577 17417 28611
rect 17451 28608 17463 28611
rect 18966 28608 18972 28620
rect 17451 28580 18972 28608
rect 17451 28577 17463 28580
rect 17405 28571 17463 28577
rect 18966 28568 18972 28580
rect 19024 28568 19030 28620
rect 20073 28611 20131 28617
rect 20073 28577 20085 28611
rect 20119 28608 20131 28611
rect 20990 28608 20996 28620
rect 20119 28580 20996 28608
rect 20119 28577 20131 28580
rect 20073 28571 20131 28577
rect 20990 28568 20996 28580
rect 21048 28568 21054 28620
rect 21358 28568 21364 28620
rect 21416 28608 21422 28620
rect 22066 28608 22094 28648
rect 22833 28645 22845 28648
rect 22879 28645 22891 28679
rect 24762 28676 24768 28688
rect 22833 28639 22891 28645
rect 23308 28648 24768 28676
rect 21416 28580 22094 28608
rect 21416 28568 21422 28580
rect 22186 28568 22192 28620
rect 22244 28608 22250 28620
rect 23308 28608 23336 28648
rect 24762 28636 24768 28648
rect 24820 28636 24826 28688
rect 22244 28580 23336 28608
rect 23385 28611 23443 28617
rect 22244 28568 22250 28580
rect 23385 28577 23397 28611
rect 23431 28608 23443 28611
rect 23658 28608 23664 28620
rect 23431 28580 23664 28608
rect 23431 28577 23443 28580
rect 23385 28571 23443 28577
rect 23658 28568 23664 28580
rect 23716 28568 23722 28620
rect 24854 28568 24860 28620
rect 24912 28608 24918 28620
rect 25041 28611 25099 28617
rect 25041 28608 25053 28611
rect 24912 28580 25053 28608
rect 24912 28568 24918 28580
rect 25041 28577 25053 28580
rect 25087 28577 25099 28611
rect 25041 28571 25099 28577
rect 25225 28611 25283 28617
rect 25225 28577 25237 28611
rect 25271 28608 25283 28611
rect 26050 28608 26056 28620
rect 25271 28580 26056 28608
rect 25271 28577 25283 28580
rect 25225 28571 25283 28577
rect 26050 28568 26056 28580
rect 26108 28568 26114 28620
rect 15102 28500 15108 28552
rect 15160 28540 15166 28552
rect 17129 28543 17187 28549
rect 17129 28540 17141 28543
rect 15160 28512 17141 28540
rect 15160 28500 15166 28512
rect 17129 28509 17141 28512
rect 17175 28509 17187 28543
rect 17129 28503 17187 28509
rect 19334 28500 19340 28552
rect 19392 28540 19398 28552
rect 20622 28540 20628 28552
rect 19392 28512 20628 28540
rect 19392 28500 19398 28512
rect 20622 28500 20628 28512
rect 20680 28500 20686 28552
rect 22278 28500 22284 28552
rect 22336 28540 22342 28552
rect 22554 28540 22560 28552
rect 22336 28512 22560 28540
rect 22336 28500 22342 28512
rect 22554 28500 22560 28512
rect 22612 28540 22618 28552
rect 23201 28543 23259 28549
rect 23201 28540 23213 28543
rect 22612 28512 23213 28540
rect 22612 28500 22618 28512
rect 23201 28509 23213 28512
rect 23247 28540 23259 28543
rect 24029 28543 24087 28549
rect 24029 28540 24041 28543
rect 23247 28512 24041 28540
rect 23247 28509 23259 28512
rect 23201 28503 23259 28509
rect 24029 28509 24041 28512
rect 24075 28509 24087 28543
rect 24029 28503 24087 28509
rect 24946 28500 24952 28552
rect 25004 28500 25010 28552
rect 9401 28475 9459 28481
rect 9401 28441 9413 28475
rect 9447 28472 9459 28475
rect 9674 28472 9680 28484
rect 9447 28444 9680 28472
rect 9447 28441 9459 28444
rect 9401 28435 9459 28441
rect 9674 28432 9680 28444
rect 9732 28432 9738 28484
rect 11606 28472 11612 28484
rect 10626 28444 11612 28472
rect 11606 28432 11612 28444
rect 11664 28432 11670 28484
rect 11701 28475 11759 28481
rect 11701 28441 11713 28475
rect 11747 28441 11759 28475
rect 11701 28435 11759 28441
rect 15197 28475 15255 28481
rect 15197 28441 15209 28475
rect 15243 28472 15255 28475
rect 16298 28472 16304 28484
rect 15243 28444 16304 28472
rect 15243 28441 15255 28444
rect 15197 28435 15255 28441
rect 11514 28364 11520 28416
rect 11572 28404 11578 28416
rect 11716 28404 11744 28435
rect 16040 28416 16068 28444
rect 16298 28432 16304 28444
rect 16356 28432 16362 28484
rect 18874 28472 18880 28484
rect 18630 28444 18880 28472
rect 18874 28432 18880 28444
rect 18932 28432 18938 28484
rect 20898 28432 20904 28484
rect 20956 28432 20962 28484
rect 23293 28475 23351 28481
rect 22126 28444 22692 28472
rect 11572 28376 11744 28404
rect 11572 28364 11578 28376
rect 14826 28364 14832 28416
rect 14884 28364 14890 28416
rect 16022 28364 16028 28416
rect 16080 28364 16086 28416
rect 16209 28407 16267 28413
rect 16209 28373 16221 28407
rect 16255 28404 16267 28407
rect 16482 28404 16488 28416
rect 16255 28376 16488 28404
rect 16255 28373 16267 28376
rect 16209 28367 16267 28373
rect 16482 28364 16488 28376
rect 16540 28364 16546 28416
rect 18690 28364 18696 28416
rect 18748 28404 18754 28416
rect 19429 28407 19487 28413
rect 19429 28404 19441 28407
rect 18748 28376 19441 28404
rect 18748 28364 18754 28376
rect 19429 28373 19441 28376
rect 19475 28373 19487 28407
rect 19429 28367 19487 28373
rect 19702 28364 19708 28416
rect 19760 28404 19766 28416
rect 19797 28407 19855 28413
rect 19797 28404 19809 28407
rect 19760 28376 19809 28404
rect 19760 28364 19766 28376
rect 19797 28373 19809 28376
rect 19843 28373 19855 28407
rect 19797 28367 19855 28373
rect 19889 28407 19947 28413
rect 19889 28373 19901 28407
rect 19935 28404 19947 28407
rect 21634 28404 21640 28416
rect 19935 28376 21640 28404
rect 19935 28373 19947 28376
rect 19889 28367 19947 28373
rect 21634 28364 21640 28376
rect 21692 28364 21698 28416
rect 21726 28364 21732 28416
rect 21784 28404 21790 28416
rect 22204 28404 22232 28444
rect 21784 28376 22232 28404
rect 22664 28404 22692 28444
rect 23293 28441 23305 28475
rect 23339 28472 23351 28475
rect 25958 28472 25964 28484
rect 23339 28444 25964 28472
rect 23339 28441 23351 28444
rect 23293 28435 23351 28441
rect 25958 28432 25964 28444
rect 26016 28432 26022 28484
rect 23934 28404 23940 28416
rect 22664 28376 23940 28404
rect 21784 28364 21790 28376
rect 23934 28364 23940 28376
rect 23992 28364 23998 28416
rect 24394 28364 24400 28416
rect 24452 28404 24458 28416
rect 24581 28407 24639 28413
rect 24581 28404 24593 28407
rect 24452 28376 24593 28404
rect 24452 28364 24458 28376
rect 24581 28373 24593 28376
rect 24627 28373 24639 28407
rect 24581 28367 24639 28373
rect 1104 28314 25852 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 25852 28314
rect 1104 28240 25852 28262
rect 11057 28203 11115 28209
rect 11057 28169 11069 28203
rect 11103 28200 11115 28203
rect 11606 28200 11612 28212
rect 11103 28172 11612 28200
rect 11103 28169 11115 28172
rect 11057 28163 11115 28169
rect 11606 28160 11612 28172
rect 11664 28160 11670 28212
rect 13722 28200 13728 28212
rect 13280 28172 13728 28200
rect 11977 28135 12035 28141
rect 11977 28132 11989 28135
rect 11072 28104 11989 28132
rect 11072 28076 11100 28104
rect 11977 28101 11989 28104
rect 12023 28101 12035 28135
rect 13280 28132 13308 28172
rect 13722 28160 13728 28172
rect 13780 28160 13786 28212
rect 15562 28160 15568 28212
rect 15620 28200 15626 28212
rect 16393 28203 16451 28209
rect 16393 28200 16405 28203
rect 15620 28172 16405 28200
rect 15620 28160 15626 28172
rect 16393 28169 16405 28172
rect 16439 28169 16451 28203
rect 16393 28163 16451 28169
rect 18874 28160 18880 28212
rect 18932 28200 18938 28212
rect 18969 28203 19027 28209
rect 18969 28200 18981 28203
rect 18932 28172 18981 28200
rect 18932 28160 18938 28172
rect 18969 28169 18981 28172
rect 19015 28169 19027 28203
rect 18969 28163 19027 28169
rect 19702 28160 19708 28212
rect 19760 28160 19766 28212
rect 21545 28203 21603 28209
rect 21545 28200 21557 28203
rect 19812 28172 21557 28200
rect 13202 28104 13308 28132
rect 11977 28095 12035 28101
rect 13446 28092 13452 28144
rect 13504 28132 13510 28144
rect 19812 28132 19840 28172
rect 21545 28169 21557 28172
rect 21591 28200 21603 28203
rect 22186 28200 22192 28212
rect 21591 28172 22192 28200
rect 21591 28169 21603 28172
rect 21545 28163 21603 28169
rect 22186 28160 22192 28172
rect 22244 28200 22250 28212
rect 22373 28203 22431 28209
rect 22373 28200 22385 28203
rect 22244 28172 22385 28200
rect 22244 28160 22250 28172
rect 22373 28169 22385 28172
rect 22419 28169 22431 28203
rect 22373 28163 22431 28169
rect 22465 28203 22523 28209
rect 22465 28169 22477 28203
rect 22511 28200 22523 28203
rect 26234 28200 26240 28212
rect 22511 28172 26240 28200
rect 22511 28169 22523 28172
rect 22465 28163 22523 28169
rect 26234 28160 26240 28172
rect 26292 28160 26298 28212
rect 13504 28104 19840 28132
rect 13504 28092 13510 28104
rect 20622 28092 20628 28144
rect 20680 28132 20686 28144
rect 21085 28135 21143 28141
rect 21085 28132 21097 28135
rect 20680 28104 21097 28132
rect 20680 28092 20686 28104
rect 21085 28101 21097 28104
rect 21131 28101 21143 28135
rect 21085 28095 21143 28101
rect 11054 28024 11060 28076
rect 11112 28024 11118 28076
rect 15657 28067 15715 28073
rect 15657 28033 15669 28067
rect 15703 28064 15715 28067
rect 16298 28064 16304 28076
rect 15703 28036 16304 28064
rect 15703 28033 15715 28036
rect 15657 28027 15715 28033
rect 16298 28024 16304 28036
rect 16356 28024 16362 28076
rect 16666 28024 16672 28076
rect 16724 28064 16730 28076
rect 17221 28067 17279 28073
rect 17221 28064 17233 28067
rect 16724 28036 17233 28064
rect 16724 28024 16730 28036
rect 17221 28033 17233 28036
rect 17267 28064 17279 28067
rect 18782 28064 18788 28076
rect 17267 28036 18788 28064
rect 17267 28033 17279 28036
rect 17221 28027 17279 28033
rect 18782 28024 18788 28036
rect 18840 28024 18846 28076
rect 20349 28067 20407 28073
rect 20349 28033 20361 28067
rect 20395 28064 20407 28067
rect 21818 28064 21824 28076
rect 20395 28036 21824 28064
rect 20395 28033 20407 28036
rect 20349 28027 20407 28033
rect 11698 27956 11704 28008
rect 11756 27956 11762 28008
rect 15749 27999 15807 28005
rect 15749 27965 15761 27999
rect 15795 27965 15807 27999
rect 15749 27959 15807 27965
rect 10778 27888 10784 27940
rect 10836 27928 10842 27940
rect 15378 27928 15384 27940
rect 10836 27900 11652 27928
rect 10836 27888 10842 27900
rect 11624 27860 11652 27900
rect 13464 27900 15384 27928
rect 13464 27869 13492 27900
rect 15378 27888 15384 27900
rect 15436 27928 15442 27940
rect 15764 27928 15792 27959
rect 16758 27956 16764 28008
rect 16816 27996 16822 28008
rect 17313 27999 17371 28005
rect 17313 27996 17325 27999
rect 16816 27968 17325 27996
rect 16816 27956 16822 27968
rect 17313 27965 17325 27968
rect 17359 27965 17371 27999
rect 17313 27959 17371 27965
rect 15436 27900 15792 27928
rect 15436 27888 15442 27900
rect 13449 27863 13507 27869
rect 13449 27860 13461 27863
rect 11624 27832 13461 27860
rect 13449 27829 13461 27832
rect 13495 27829 13507 27863
rect 13449 27823 13507 27829
rect 13814 27820 13820 27872
rect 13872 27860 13878 27872
rect 15197 27863 15255 27869
rect 15197 27860 15209 27863
rect 13872 27832 15209 27860
rect 13872 27820 13878 27832
rect 15197 27829 15209 27832
rect 15243 27829 15255 27863
rect 15197 27823 15255 27829
rect 16298 27820 16304 27872
rect 16356 27820 16362 27872
rect 16850 27820 16856 27872
rect 16908 27820 16914 27872
rect 17328 27860 17356 27959
rect 17402 27956 17408 28008
rect 17460 27956 17466 28008
rect 17954 27956 17960 28008
rect 18012 27996 18018 28008
rect 18049 27999 18107 28005
rect 18049 27996 18061 27999
rect 18012 27968 18061 27996
rect 18012 27956 18018 27968
rect 18049 27965 18061 27968
rect 18095 27965 18107 27999
rect 18049 27959 18107 27965
rect 17678 27888 17684 27940
rect 17736 27928 17742 27940
rect 19337 27931 19395 27937
rect 19337 27928 19349 27931
rect 17736 27900 19349 27928
rect 17736 27888 17742 27900
rect 19337 27897 19349 27900
rect 19383 27928 19395 27931
rect 20364 27928 20392 28027
rect 21818 28024 21824 28036
rect 21876 28024 21882 28076
rect 22557 27999 22615 28005
rect 22557 27965 22569 27999
rect 22603 27965 22615 27999
rect 22557 27959 22615 27965
rect 22005 27931 22063 27937
rect 22005 27928 22017 27931
rect 19383 27900 20392 27928
rect 20456 27900 22017 27928
rect 19383 27897 19395 27900
rect 19337 27891 19395 27897
rect 18506 27860 18512 27872
rect 17328 27832 18512 27860
rect 18506 27820 18512 27832
rect 18564 27820 18570 27872
rect 18782 27820 18788 27872
rect 18840 27820 18846 27872
rect 19150 27820 19156 27872
rect 19208 27860 19214 27872
rect 20456 27860 20484 27900
rect 22005 27897 22017 27900
rect 22051 27897 22063 27931
rect 22005 27891 22063 27897
rect 22094 27888 22100 27940
rect 22152 27928 22158 27940
rect 22572 27928 22600 27959
rect 22830 27956 22836 28008
rect 22888 27996 22894 28008
rect 23201 27999 23259 28005
rect 23201 27996 23213 27999
rect 22888 27968 23213 27996
rect 22888 27956 22894 27968
rect 23201 27965 23213 27968
rect 23247 27965 23259 27999
rect 23201 27959 23259 27965
rect 23474 27956 23480 28008
rect 23532 27956 23538 28008
rect 23934 27956 23940 28008
rect 23992 27996 23998 28008
rect 24504 27996 24532 28118
rect 23992 27968 25268 27996
rect 23992 27956 23998 27968
rect 22152 27900 22600 27928
rect 22152 27888 22158 27900
rect 25240 27872 25268 27968
rect 19208 27832 20484 27860
rect 19208 27820 19214 27832
rect 22370 27820 22376 27872
rect 22428 27860 22434 27872
rect 22554 27860 22560 27872
rect 22428 27832 22560 27860
rect 22428 27820 22434 27832
rect 22554 27820 22560 27832
rect 22612 27860 22618 27872
rect 24949 27863 25007 27869
rect 24949 27860 24961 27863
rect 22612 27832 24961 27860
rect 22612 27820 22618 27832
rect 24949 27829 24961 27832
rect 24995 27829 25007 27863
rect 24949 27823 25007 27829
rect 25222 27820 25228 27872
rect 25280 27820 25286 27872
rect 25406 27820 25412 27872
rect 25464 27820 25470 27872
rect 1104 27770 25852 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 25852 27770
rect 1104 27696 25852 27718
rect 11422 27656 11428 27668
rect 10612 27628 11428 27656
rect 10505 27523 10563 27529
rect 10505 27489 10517 27523
rect 10551 27520 10563 27523
rect 10612 27520 10640 27628
rect 11422 27616 11428 27628
rect 11480 27616 11486 27668
rect 12621 27659 12679 27665
rect 12621 27656 12633 27659
rect 12406 27628 12633 27656
rect 12406 27588 12434 27628
rect 12621 27625 12633 27628
rect 12667 27656 12679 27659
rect 12710 27656 12716 27668
rect 12667 27628 12716 27656
rect 12667 27625 12679 27628
rect 12621 27619 12679 27625
rect 12710 27616 12716 27628
rect 12768 27616 12774 27668
rect 15102 27656 15108 27668
rect 13096 27628 15108 27656
rect 13096 27600 13124 27628
rect 15102 27616 15108 27628
rect 15160 27616 15166 27668
rect 18874 27616 18880 27668
rect 18932 27656 18938 27668
rect 19978 27656 19984 27668
rect 18932 27628 19984 27656
rect 18932 27616 18938 27628
rect 19978 27616 19984 27628
rect 20036 27616 20042 27668
rect 20152 27659 20210 27665
rect 20152 27625 20164 27659
rect 20198 27656 20210 27659
rect 23658 27656 23664 27668
rect 20198 27628 23664 27656
rect 20198 27625 20210 27628
rect 20152 27619 20210 27625
rect 23658 27616 23664 27628
rect 23716 27656 23722 27668
rect 23845 27659 23903 27665
rect 23845 27656 23857 27659
rect 23716 27628 23857 27656
rect 23716 27616 23722 27628
rect 23845 27625 23857 27628
rect 23891 27625 23903 27659
rect 23845 27619 23903 27625
rect 11900 27560 12434 27588
rect 10551 27492 10640 27520
rect 10551 27489 10563 27492
rect 10505 27483 10563 27489
rect 10778 27480 10784 27532
rect 10836 27480 10842 27532
rect 11900 27438 11928 27560
rect 13078 27548 13084 27600
rect 13136 27548 13142 27600
rect 16114 27548 16120 27600
rect 16172 27588 16178 27600
rect 17497 27591 17555 27597
rect 17497 27588 17509 27591
rect 16172 27560 17509 27588
rect 16172 27548 16178 27560
rect 17497 27557 17509 27560
rect 17543 27557 17555 27591
rect 17497 27551 17555 27557
rect 23474 27548 23480 27600
rect 23532 27588 23538 27600
rect 24762 27588 24768 27600
rect 23532 27560 24768 27588
rect 23532 27548 23538 27560
rect 24762 27548 24768 27560
rect 24820 27588 24826 27600
rect 24820 27560 25176 27588
rect 24820 27548 24826 27560
rect 13541 27523 13599 27529
rect 13541 27520 13553 27523
rect 12406 27492 13553 27520
rect 9306 27276 9312 27328
rect 9364 27316 9370 27328
rect 12253 27319 12311 27325
rect 12253 27316 12265 27319
rect 9364 27288 12265 27316
rect 9364 27276 9370 27288
rect 12253 27285 12265 27288
rect 12299 27316 12311 27319
rect 12406 27316 12434 27492
rect 13541 27489 13553 27492
rect 13587 27489 13599 27523
rect 13541 27483 13599 27489
rect 15102 27480 15108 27532
rect 15160 27520 15166 27532
rect 15749 27523 15807 27529
rect 15749 27520 15761 27523
rect 15160 27492 15761 27520
rect 15160 27480 15166 27492
rect 15749 27489 15761 27492
rect 15795 27489 15807 27523
rect 15749 27483 15807 27489
rect 17770 27480 17776 27532
rect 17828 27520 17834 27532
rect 18049 27523 18107 27529
rect 18049 27520 18061 27523
rect 17828 27492 18061 27520
rect 17828 27480 17834 27492
rect 18049 27489 18061 27492
rect 18095 27489 18107 27523
rect 18049 27483 18107 27489
rect 19889 27523 19947 27529
rect 19889 27489 19901 27523
rect 19935 27520 19947 27523
rect 22097 27523 22155 27529
rect 22097 27520 22109 27523
rect 19935 27492 22109 27520
rect 19935 27489 19947 27492
rect 19889 27483 19947 27489
rect 22097 27489 22109 27492
rect 22143 27520 22155 27523
rect 22830 27520 22836 27532
rect 22143 27492 22836 27520
rect 22143 27489 22155 27492
rect 22097 27483 22155 27489
rect 22830 27480 22836 27492
rect 22888 27480 22894 27532
rect 24118 27480 24124 27532
rect 24176 27480 24182 27532
rect 25038 27480 25044 27532
rect 25096 27480 25102 27532
rect 25148 27529 25176 27560
rect 25133 27523 25191 27529
rect 25133 27489 25145 27523
rect 25179 27489 25191 27523
rect 25133 27483 25191 27489
rect 13449 27455 13507 27461
rect 13449 27421 13461 27455
rect 13495 27452 13507 27455
rect 14826 27452 14832 27464
rect 13495 27424 14832 27452
rect 13495 27421 13507 27424
rect 13449 27415 13507 27421
rect 14826 27412 14832 27424
rect 14884 27412 14890 27464
rect 17865 27455 17923 27461
rect 17865 27421 17877 27455
rect 17911 27452 17923 27455
rect 17954 27452 17960 27464
rect 17911 27424 17960 27452
rect 17911 27421 17923 27424
rect 17865 27415 17923 27421
rect 17954 27412 17960 27424
rect 18012 27412 18018 27464
rect 23934 27452 23940 27464
rect 23506 27424 23940 27452
rect 23934 27412 23940 27424
rect 23992 27412 23998 27464
rect 24949 27455 25007 27461
rect 24949 27421 24961 27455
rect 24995 27452 25007 27455
rect 25406 27452 25412 27464
rect 24995 27424 25412 27452
rect 24995 27421 25007 27424
rect 24949 27415 25007 27421
rect 25406 27412 25412 27424
rect 25464 27412 25470 27464
rect 13357 27387 13415 27393
rect 13357 27353 13369 27387
rect 13403 27384 13415 27387
rect 13814 27384 13820 27396
rect 13403 27356 13820 27384
rect 13403 27353 13415 27356
rect 13357 27347 13415 27353
rect 13814 27344 13820 27356
rect 13872 27344 13878 27396
rect 16022 27384 16028 27396
rect 15580 27356 16028 27384
rect 12299 27288 12434 27316
rect 12299 27285 12311 27288
rect 12253 27279 12311 27285
rect 12618 27276 12624 27328
rect 12676 27316 12682 27328
rect 12989 27319 13047 27325
rect 12989 27316 13001 27319
rect 12676 27288 13001 27316
rect 12676 27276 12682 27288
rect 12989 27285 13001 27288
rect 13035 27285 13047 27319
rect 12989 27279 13047 27285
rect 13722 27276 13728 27328
rect 13780 27316 13786 27328
rect 15197 27319 15255 27325
rect 15197 27316 15209 27319
rect 13780 27288 15209 27316
rect 13780 27276 13786 27288
rect 15197 27285 15209 27288
rect 15243 27285 15255 27319
rect 15197 27279 15255 27285
rect 15470 27276 15476 27328
rect 15528 27316 15534 27328
rect 15580 27325 15608 27356
rect 16022 27344 16028 27356
rect 16080 27384 16086 27396
rect 16209 27387 16267 27393
rect 16209 27384 16221 27387
rect 16080 27356 16221 27384
rect 16080 27344 16086 27356
rect 16209 27353 16221 27356
rect 16255 27353 16267 27387
rect 16209 27347 16267 27353
rect 20070 27344 20076 27396
rect 20128 27384 20134 27396
rect 20128 27356 20654 27384
rect 20128 27344 20134 27356
rect 22370 27344 22376 27396
rect 22428 27344 22434 27396
rect 23658 27344 23664 27396
rect 23716 27384 23722 27396
rect 23716 27356 24624 27384
rect 23716 27344 23722 27356
rect 15565 27319 15623 27325
rect 15565 27316 15577 27319
rect 15528 27288 15577 27316
rect 15528 27276 15534 27288
rect 15565 27285 15577 27288
rect 15611 27285 15623 27319
rect 15565 27279 15623 27285
rect 15657 27319 15715 27325
rect 15657 27285 15669 27319
rect 15703 27316 15715 27319
rect 16482 27316 16488 27328
rect 15703 27288 16488 27316
rect 15703 27285 15715 27288
rect 15657 27279 15715 27285
rect 16482 27276 16488 27288
rect 16540 27276 16546 27328
rect 17586 27276 17592 27328
rect 17644 27316 17650 27328
rect 17957 27319 18015 27325
rect 17957 27316 17969 27319
rect 17644 27288 17969 27316
rect 17644 27276 17650 27288
rect 17957 27285 17969 27288
rect 18003 27285 18015 27319
rect 17957 27279 18015 27285
rect 21634 27276 21640 27328
rect 21692 27276 21698 27328
rect 24596 27325 24624 27356
rect 24581 27319 24639 27325
rect 24581 27285 24593 27319
rect 24627 27285 24639 27319
rect 24581 27279 24639 27285
rect 1104 27226 25852 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 25852 27226
rect 1104 27152 25852 27174
rect 9766 27112 9772 27124
rect 9324 27084 9772 27112
rect 9324 26985 9352 27084
rect 9766 27072 9772 27084
rect 9824 27112 9830 27124
rect 10870 27112 10876 27124
rect 9824 27084 10876 27112
rect 9824 27072 9830 27084
rect 10870 27072 10876 27084
rect 10928 27112 10934 27124
rect 11698 27112 11704 27124
rect 10928 27084 11704 27112
rect 10928 27072 10934 27084
rect 11698 27072 11704 27084
rect 11756 27072 11762 27124
rect 12710 27112 12716 27124
rect 12406 27084 12716 27112
rect 11146 27044 11152 27056
rect 10810 27016 11152 27044
rect 11146 27004 11152 27016
rect 11204 27044 11210 27056
rect 11609 27047 11667 27053
rect 11609 27044 11621 27047
rect 11204 27016 11621 27044
rect 11204 27004 11210 27016
rect 11609 27013 11621 27016
rect 11655 27044 11667 27047
rect 12406 27044 12434 27084
rect 12710 27072 12716 27084
rect 12768 27112 12774 27124
rect 15194 27112 15200 27124
rect 12768 27084 15200 27112
rect 12768 27072 12774 27084
rect 11655 27016 12434 27044
rect 13357 27047 13415 27053
rect 11655 27013 11667 27016
rect 11609 27007 11667 27013
rect 13357 27013 13369 27047
rect 13403 27044 13415 27047
rect 13630 27044 13636 27056
rect 13403 27016 13636 27044
rect 13403 27013 13415 27016
rect 13357 27007 13415 27013
rect 13630 27004 13636 27016
rect 13688 27004 13694 27056
rect 13740 27044 13768 27084
rect 15194 27072 15200 27084
rect 15252 27072 15258 27124
rect 15657 27115 15715 27121
rect 15657 27081 15669 27115
rect 15703 27112 15715 27115
rect 16850 27112 16856 27124
rect 15703 27084 16856 27112
rect 15703 27081 15715 27084
rect 15657 27075 15715 27081
rect 16850 27072 16856 27084
rect 16908 27072 16914 27124
rect 19242 27112 19248 27124
rect 18064 27084 19248 27112
rect 13740 27016 13846 27044
rect 15746 27004 15752 27056
rect 15804 27004 15810 27056
rect 18064 27044 18092 27084
rect 19242 27072 19248 27084
rect 19300 27072 19306 27124
rect 19978 27072 19984 27124
rect 20036 27072 20042 27124
rect 22738 27072 22744 27124
rect 22796 27112 22802 27124
rect 22833 27115 22891 27121
rect 22833 27112 22845 27115
rect 22796 27084 22845 27112
rect 22796 27072 22802 27084
rect 22833 27081 22845 27084
rect 22879 27081 22891 27115
rect 22833 27075 22891 27081
rect 24762 27072 24768 27124
rect 24820 27112 24826 27124
rect 25317 27115 25375 27121
rect 25317 27112 25329 27115
rect 24820 27084 25329 27112
rect 24820 27072 24826 27084
rect 25317 27081 25329 27084
rect 25363 27081 25375 27115
rect 25317 27075 25375 27081
rect 17972 27016 18092 27044
rect 9309 26979 9367 26985
rect 9309 26945 9321 26979
rect 9355 26945 9367 26979
rect 9309 26939 9367 26945
rect 11698 26936 11704 26988
rect 11756 26976 11762 26988
rect 12802 26976 12808 26988
rect 11756 26948 12808 26976
rect 11756 26936 11762 26948
rect 12802 26936 12808 26948
rect 12860 26976 12866 26988
rect 13078 26976 13084 26988
rect 12860 26948 13084 26976
rect 12860 26936 12866 26948
rect 13078 26936 13084 26948
rect 13136 26936 13142 26988
rect 14826 26936 14832 26988
rect 14884 26976 14890 26988
rect 16574 26976 16580 26988
rect 14884 26948 16580 26976
rect 14884 26936 14890 26948
rect 16574 26936 16580 26948
rect 16632 26936 16638 26988
rect 17972 26985 18000 27016
rect 18874 27004 18880 27056
rect 18932 27004 18938 27056
rect 22922 27004 22928 27056
rect 22980 27004 22986 27056
rect 25222 27044 25228 27056
rect 25070 27016 25228 27044
rect 25222 27004 25228 27016
rect 25280 27044 25286 27056
rect 26234 27044 26240 27056
rect 25280 27016 26240 27044
rect 25280 27004 25286 27016
rect 26234 27004 26240 27016
rect 26292 27004 26298 27056
rect 17957 26979 18015 26985
rect 17957 26945 17969 26979
rect 18003 26945 18015 26979
rect 17957 26939 18015 26945
rect 22646 26936 22652 26988
rect 22704 26976 22710 26988
rect 22741 26979 22799 26985
rect 22741 26976 22753 26979
rect 22704 26948 22753 26976
rect 22704 26936 22710 26948
rect 22741 26945 22753 26948
rect 22787 26945 22799 26979
rect 22940 26976 22968 27004
rect 23290 26976 23296 26988
rect 22940 26948 23296 26976
rect 22741 26939 22799 26945
rect 23290 26936 23296 26948
rect 23348 26976 23354 26988
rect 23569 26979 23627 26985
rect 23569 26976 23581 26979
rect 23348 26948 23581 26976
rect 23348 26936 23354 26948
rect 23569 26945 23581 26948
rect 23615 26945 23627 26979
rect 23569 26939 23627 26945
rect 9585 26911 9643 26917
rect 9585 26908 9597 26911
rect 9324 26880 9597 26908
rect 9324 26852 9352 26880
rect 9585 26877 9597 26880
rect 9631 26877 9643 26911
rect 9585 26871 9643 26877
rect 11057 26911 11115 26917
rect 11057 26877 11069 26911
rect 11103 26908 11115 26911
rect 11330 26908 11336 26920
rect 11103 26880 11336 26908
rect 11103 26877 11115 26880
rect 11057 26871 11115 26877
rect 11330 26868 11336 26880
rect 11388 26868 11394 26920
rect 13446 26908 13452 26920
rect 12406 26880 13452 26908
rect 9306 26800 9312 26852
rect 9364 26800 9370 26852
rect 12406 26840 12434 26880
rect 13446 26868 13452 26880
rect 13504 26868 13510 26920
rect 15841 26911 15899 26917
rect 15841 26877 15853 26911
rect 15887 26877 15899 26911
rect 15841 26871 15899 26877
rect 18233 26911 18291 26917
rect 18233 26877 18245 26911
rect 18279 26908 18291 26911
rect 22094 26908 22100 26920
rect 18279 26880 22100 26908
rect 18279 26877 18291 26880
rect 18233 26871 18291 26877
rect 15856 26840 15884 26871
rect 22094 26868 22100 26880
rect 22152 26868 22158 26920
rect 23017 26911 23075 26917
rect 23017 26877 23029 26911
rect 23063 26908 23075 26911
rect 23474 26908 23480 26920
rect 23063 26880 23480 26908
rect 23063 26877 23075 26880
rect 23017 26871 23075 26877
rect 23474 26868 23480 26880
rect 23532 26868 23538 26920
rect 23845 26911 23903 26917
rect 23845 26877 23857 26911
rect 23891 26908 23903 26911
rect 25590 26908 25596 26920
rect 23891 26880 25596 26908
rect 23891 26877 23903 26880
rect 23845 26871 23903 26877
rect 25590 26868 25596 26880
rect 25648 26868 25654 26920
rect 10612 26812 12434 26840
rect 14844 26812 15884 26840
rect 3418 26732 3424 26784
rect 3476 26772 3482 26784
rect 10612 26772 10640 26812
rect 3476 26744 10640 26772
rect 3476 26732 3482 26744
rect 11974 26732 11980 26784
rect 12032 26772 12038 26784
rect 14844 26781 14872 26812
rect 14829 26775 14887 26781
rect 14829 26772 14841 26775
rect 12032 26744 14841 26772
rect 12032 26732 12038 26744
rect 14829 26741 14841 26744
rect 14875 26741 14887 26775
rect 14829 26735 14887 26741
rect 14918 26732 14924 26784
rect 14976 26772 14982 26784
rect 15289 26775 15347 26781
rect 15289 26772 15301 26775
rect 14976 26744 15301 26772
rect 14976 26732 14982 26744
rect 15289 26741 15301 26744
rect 15335 26741 15347 26775
rect 15289 26735 15347 26741
rect 18966 26732 18972 26784
rect 19024 26772 19030 26784
rect 19705 26775 19763 26781
rect 19705 26772 19717 26775
rect 19024 26744 19717 26772
rect 19024 26732 19030 26744
rect 19705 26741 19717 26744
rect 19751 26741 19763 26775
rect 19705 26735 19763 26741
rect 21818 26732 21824 26784
rect 21876 26732 21882 26784
rect 22370 26732 22376 26784
rect 22428 26732 22434 26784
rect 24854 26732 24860 26784
rect 24912 26772 24918 26784
rect 25958 26772 25964 26784
rect 24912 26744 25964 26772
rect 24912 26732 24918 26744
rect 25958 26732 25964 26744
rect 26016 26732 26022 26784
rect 1104 26682 25852 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 25852 26682
rect 1104 26608 25852 26630
rect 11146 26528 11152 26580
rect 11204 26528 11210 26580
rect 13630 26528 13636 26580
rect 13688 26568 13694 26580
rect 15657 26571 15715 26577
rect 15657 26568 15669 26571
rect 13688 26540 15669 26568
rect 13688 26528 13694 26540
rect 15657 26537 15669 26540
rect 15703 26537 15715 26571
rect 15657 26531 15715 26537
rect 16022 26528 16028 26580
rect 16080 26568 16086 26580
rect 17034 26568 17040 26580
rect 16080 26540 17040 26568
rect 16080 26528 16086 26540
rect 17034 26528 17040 26540
rect 17092 26568 17098 26580
rect 17221 26571 17279 26577
rect 17221 26568 17233 26571
rect 17092 26540 17233 26568
rect 17092 26528 17098 26540
rect 17221 26537 17233 26540
rect 17267 26537 17279 26571
rect 17221 26531 17279 26537
rect 17586 26528 17592 26580
rect 17644 26568 17650 26580
rect 19886 26568 19892 26580
rect 17644 26540 19892 26568
rect 17644 26528 17650 26540
rect 19886 26528 19892 26540
rect 19944 26528 19950 26580
rect 20070 26528 20076 26580
rect 20128 26568 20134 26580
rect 21177 26571 21235 26577
rect 20128 26540 20760 26568
rect 20128 26528 20134 26540
rect 9125 26435 9183 26441
rect 9125 26401 9137 26435
rect 9171 26432 9183 26435
rect 9766 26432 9772 26444
rect 9171 26404 9772 26432
rect 9171 26401 9183 26404
rect 9125 26395 9183 26401
rect 9766 26392 9772 26404
rect 9824 26392 9830 26444
rect 10873 26435 10931 26441
rect 10873 26401 10885 26435
rect 10919 26432 10931 26435
rect 11054 26432 11060 26444
rect 10919 26404 11060 26432
rect 10919 26401 10931 26404
rect 10873 26395 10931 26401
rect 11054 26392 11060 26404
rect 11112 26392 11118 26444
rect 11164 26364 11192 26528
rect 11606 26460 11612 26512
rect 11664 26500 11670 26512
rect 14277 26503 14335 26509
rect 14277 26500 14289 26503
rect 11664 26472 14289 26500
rect 11664 26460 11670 26472
rect 14277 26469 14289 26472
rect 14323 26469 14335 26503
rect 20732 26500 20760 26540
rect 21177 26537 21189 26571
rect 21223 26568 21235 26571
rect 22094 26568 22100 26580
rect 21223 26540 22100 26568
rect 21223 26537 21235 26540
rect 21177 26531 21235 26537
rect 22094 26528 22100 26540
rect 22152 26528 22158 26580
rect 22278 26528 22284 26580
rect 22336 26528 22342 26580
rect 23845 26571 23903 26577
rect 23845 26537 23857 26571
rect 23891 26568 23903 26571
rect 24946 26568 24952 26580
rect 23891 26540 24952 26568
rect 23891 26537 23903 26540
rect 23845 26531 23903 26537
rect 24946 26528 24952 26540
rect 25004 26528 25010 26580
rect 21082 26500 21088 26512
rect 14277 26463 14335 26469
rect 14476 26472 16896 26500
rect 20732 26472 21088 26500
rect 10534 26336 11192 26364
rect 8570 26256 8576 26308
rect 8628 26296 8634 26308
rect 9401 26299 9459 26305
rect 9401 26296 9413 26299
rect 8628 26268 9413 26296
rect 8628 26256 8634 26268
rect 9401 26265 9413 26268
rect 9447 26296 9459 26299
rect 11333 26299 11391 26305
rect 11333 26296 11345 26299
rect 9447 26268 9812 26296
rect 9447 26265 9459 26268
rect 9401 26259 9459 26265
rect 9784 26228 9812 26268
rect 10704 26268 11345 26296
rect 10704 26228 10732 26268
rect 11333 26265 11345 26268
rect 11379 26296 11391 26299
rect 11790 26296 11796 26308
rect 11379 26268 11796 26296
rect 11379 26265 11391 26268
rect 11333 26259 11391 26265
rect 11790 26256 11796 26268
rect 11848 26256 11854 26308
rect 14476 26296 14504 26472
rect 14921 26435 14979 26441
rect 14921 26401 14933 26435
rect 14967 26432 14979 26435
rect 15010 26432 15016 26444
rect 14967 26404 15016 26432
rect 14967 26401 14979 26404
rect 14921 26395 14979 26401
rect 15010 26392 15016 26404
rect 15068 26392 15074 26444
rect 15194 26392 15200 26444
rect 15252 26432 15258 26444
rect 15289 26435 15347 26441
rect 15289 26432 15301 26435
rect 15252 26404 15301 26432
rect 15252 26392 15258 26404
rect 15289 26401 15301 26404
rect 15335 26401 15347 26435
rect 15289 26395 15347 26401
rect 16209 26435 16267 26441
rect 16209 26401 16221 26435
rect 16255 26401 16267 26435
rect 16209 26395 16267 26401
rect 14550 26324 14556 26376
rect 14608 26364 14614 26376
rect 15102 26364 15108 26376
rect 14608 26336 15108 26364
rect 14608 26324 14614 26336
rect 15102 26324 15108 26336
rect 15160 26364 15166 26376
rect 16224 26364 16252 26395
rect 16574 26392 16580 26444
rect 16632 26432 16638 26444
rect 16669 26435 16727 26441
rect 16669 26432 16681 26435
rect 16632 26404 16681 26432
rect 16632 26392 16638 26404
rect 16669 26401 16681 26404
rect 16715 26401 16727 26435
rect 16669 26395 16727 26401
rect 16868 26373 16896 26472
rect 21082 26460 21088 26472
rect 21140 26500 21146 26512
rect 21453 26503 21511 26509
rect 21453 26500 21465 26503
rect 21140 26472 21465 26500
rect 21140 26460 21146 26472
rect 21453 26469 21465 26472
rect 21499 26500 21511 26503
rect 21818 26500 21824 26512
rect 21499 26472 21824 26500
rect 21499 26469 21511 26472
rect 21453 26463 21511 26469
rect 21818 26460 21824 26472
rect 21876 26460 21882 26512
rect 22296 26500 22324 26528
rect 22204 26472 22324 26500
rect 17402 26432 17408 26444
rect 17039 26404 17408 26432
rect 15160 26336 16252 26364
rect 16853 26367 16911 26373
rect 15160 26324 15166 26336
rect 16853 26333 16865 26367
rect 16899 26364 16911 26367
rect 16942 26364 16948 26376
rect 16899 26336 16948 26364
rect 16899 26333 16911 26336
rect 16853 26327 16911 26333
rect 16942 26324 16948 26336
rect 17000 26364 17006 26376
rect 17039 26364 17067 26404
rect 17402 26392 17408 26404
rect 17460 26392 17466 26444
rect 19426 26392 19432 26444
rect 19484 26392 19490 26444
rect 19705 26435 19763 26441
rect 19705 26401 19717 26435
rect 19751 26432 19763 26435
rect 20990 26432 20996 26444
rect 19751 26404 20996 26432
rect 19751 26401 19763 26404
rect 19705 26395 19763 26401
rect 20990 26392 20996 26404
rect 21048 26432 21054 26444
rect 21634 26432 21640 26444
rect 21048 26404 21640 26432
rect 21048 26392 21054 26404
rect 21634 26392 21640 26404
rect 21692 26392 21698 26444
rect 17000 26336 17067 26364
rect 17129 26367 17187 26373
rect 17000 26324 17006 26336
rect 17129 26333 17141 26367
rect 17175 26364 17187 26367
rect 17218 26364 17224 26376
rect 17175 26336 17224 26364
rect 17175 26333 17187 26336
rect 17129 26327 17187 26333
rect 14645 26299 14703 26305
rect 14645 26296 14657 26299
rect 14476 26268 14657 26296
rect 14645 26265 14657 26268
rect 14691 26265 14703 26299
rect 14645 26259 14703 26265
rect 14737 26299 14795 26305
rect 14737 26265 14749 26299
rect 14783 26296 14795 26299
rect 14826 26296 14832 26308
rect 14783 26268 14832 26296
rect 14783 26265 14795 26268
rect 14737 26259 14795 26265
rect 14826 26256 14832 26268
rect 14884 26256 14890 26308
rect 15562 26256 15568 26308
rect 15620 26296 15626 26308
rect 16022 26296 16028 26308
rect 15620 26268 16028 26296
rect 15620 26256 15626 26268
rect 16022 26256 16028 26268
rect 16080 26256 16086 26308
rect 16117 26299 16175 26305
rect 16117 26265 16129 26299
rect 16163 26296 16175 26299
rect 16298 26296 16304 26308
rect 16163 26268 16304 26296
rect 16163 26265 16175 26268
rect 16117 26259 16175 26265
rect 16298 26256 16304 26268
rect 16356 26296 16362 26308
rect 17144 26296 17172 26327
rect 17218 26324 17224 26336
rect 17276 26324 17282 26376
rect 22204 26364 22232 26472
rect 22554 26460 22560 26512
rect 22612 26500 22618 26512
rect 22649 26503 22707 26509
rect 22649 26500 22661 26503
rect 22612 26472 22661 26500
rect 22612 26460 22618 26472
rect 22649 26469 22661 26472
rect 22695 26469 22707 26503
rect 22649 26463 22707 26469
rect 24581 26503 24639 26509
rect 24581 26469 24593 26503
rect 24627 26500 24639 26503
rect 25038 26500 25044 26512
rect 24627 26472 25044 26500
rect 24627 26469 24639 26472
rect 24581 26463 24639 26469
rect 25038 26460 25044 26472
rect 25096 26460 25102 26512
rect 22278 26392 22284 26444
rect 22336 26432 22342 26444
rect 23201 26435 23259 26441
rect 23201 26432 23213 26435
rect 22336 26404 23213 26432
rect 22336 26392 22342 26404
rect 23201 26401 23213 26404
rect 23247 26401 23259 26435
rect 25130 26432 25136 26444
rect 23201 26395 23259 26401
rect 25056 26404 25136 26432
rect 22738 26364 22744 26376
rect 22204 26336 22744 26364
rect 22738 26324 22744 26336
rect 22796 26364 22802 26376
rect 23017 26367 23075 26373
rect 23017 26364 23029 26367
rect 22796 26336 23029 26364
rect 22796 26324 22802 26336
rect 23017 26333 23029 26336
rect 23063 26333 23075 26367
rect 23017 26327 23075 26333
rect 23109 26367 23167 26373
rect 23109 26333 23121 26367
rect 23155 26364 23167 26367
rect 23382 26364 23388 26376
rect 23155 26336 23388 26364
rect 23155 26333 23167 26336
rect 23109 26327 23167 26333
rect 23382 26324 23388 26336
rect 23440 26324 23446 26376
rect 24026 26324 24032 26376
rect 24084 26324 24090 26376
rect 24854 26324 24860 26376
rect 24912 26364 24918 26376
rect 25056 26373 25084 26404
rect 25130 26392 25136 26404
rect 25188 26392 25194 26444
rect 25222 26392 25228 26444
rect 25280 26392 25286 26444
rect 25406 26392 25412 26444
rect 25464 26392 25470 26444
rect 24949 26367 25007 26373
rect 24949 26364 24961 26367
rect 24912 26336 24961 26364
rect 24912 26324 24918 26336
rect 24949 26333 24961 26336
rect 24995 26333 25007 26367
rect 24949 26327 25007 26333
rect 25041 26367 25099 26373
rect 25041 26333 25053 26367
rect 25087 26333 25099 26367
rect 25041 26327 25099 26333
rect 16356 26268 17172 26296
rect 16356 26256 16362 26268
rect 19978 26256 19984 26308
rect 20036 26296 20042 26308
rect 20036 26268 20194 26296
rect 20036 26256 20042 26268
rect 25130 26256 25136 26308
rect 25188 26296 25194 26308
rect 25424 26296 25452 26392
rect 25866 26324 25872 26376
rect 25924 26324 25930 26376
rect 25188 26268 25452 26296
rect 25188 26256 25194 26268
rect 25590 26256 25596 26308
rect 25648 26296 25654 26308
rect 25884 26296 25912 26324
rect 25648 26268 25912 26296
rect 25648 26256 25654 26268
rect 9784 26200 10732 26228
rect 18233 26231 18291 26237
rect 18233 26197 18245 26231
rect 18279 26228 18291 26231
rect 18322 26228 18328 26240
rect 18279 26200 18328 26228
rect 18279 26197 18291 26200
rect 18233 26191 18291 26197
rect 18322 26188 18328 26200
rect 18380 26188 18386 26240
rect 1104 26138 25852 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 25852 26138
rect 1104 26064 25852 26086
rect 12618 25984 12624 26036
rect 12676 25984 12682 26036
rect 14001 26027 14059 26033
rect 14001 25993 14013 26027
rect 14047 26024 14059 26027
rect 14642 26024 14648 26036
rect 14047 25996 14648 26024
rect 14047 25993 14059 25996
rect 14001 25987 14059 25993
rect 14642 25984 14648 25996
rect 14700 25984 14706 26036
rect 14829 26027 14887 26033
rect 14829 25993 14841 26027
rect 14875 25993 14887 26027
rect 14829 25987 14887 25993
rect 15289 26027 15347 26033
rect 15289 25993 15301 26027
rect 15335 26024 15347 26027
rect 15335 25996 16252 26024
rect 15335 25993 15347 25996
rect 15289 25987 15347 25993
rect 10686 25916 10692 25968
rect 10744 25956 10750 25968
rect 13909 25959 13967 25965
rect 13909 25956 13921 25959
rect 10744 25928 13921 25956
rect 10744 25916 10750 25928
rect 13909 25925 13921 25928
rect 13955 25925 13967 25959
rect 13909 25919 13967 25925
rect 14182 25916 14188 25968
rect 14240 25956 14246 25968
rect 14844 25956 14872 25987
rect 14240 25928 14872 25956
rect 16224 25956 16252 25996
rect 16298 25984 16304 26036
rect 16356 26024 16362 26036
rect 17773 26027 17831 26033
rect 17773 26024 17785 26027
rect 16356 25996 17785 26024
rect 16356 25984 16362 25996
rect 17773 25993 17785 25996
rect 17819 25993 17831 26027
rect 17773 25987 17831 25993
rect 18141 26027 18199 26033
rect 18141 25993 18153 26027
rect 18187 26024 18199 26027
rect 18322 26024 18328 26036
rect 18187 25996 18328 26024
rect 18187 25993 18199 25996
rect 18141 25987 18199 25993
rect 18322 25984 18328 25996
rect 18380 25984 18386 26036
rect 18874 25984 18880 26036
rect 18932 26024 18938 26036
rect 19153 26027 19211 26033
rect 19153 26024 19165 26027
rect 18932 25996 19165 26024
rect 18932 25984 18938 25996
rect 19153 25993 19165 25996
rect 19199 26024 19211 26027
rect 20162 26024 20168 26036
rect 19199 25996 20168 26024
rect 19199 25993 19211 25996
rect 19153 25987 19211 25993
rect 20162 25984 20168 25996
rect 20220 25984 20226 26036
rect 22462 25984 22468 26036
rect 22520 25984 22526 26036
rect 25130 26024 25136 26036
rect 23400 25996 25136 26024
rect 17405 25959 17463 25965
rect 17405 25956 17417 25959
rect 16224 25928 17417 25956
rect 14240 25916 14246 25928
rect 17405 25925 17417 25928
rect 17451 25956 17463 25959
rect 17586 25956 17592 25968
rect 17451 25928 17592 25956
rect 17451 25925 17463 25928
rect 17405 25919 17463 25925
rect 17586 25916 17592 25928
rect 17644 25916 17650 25968
rect 18233 25959 18291 25965
rect 18233 25925 18245 25959
rect 18279 25956 18291 25959
rect 18414 25956 18420 25968
rect 18279 25928 18420 25956
rect 18279 25925 18291 25928
rect 18233 25919 18291 25925
rect 18414 25916 18420 25928
rect 18472 25916 18478 25968
rect 23400 25956 23428 25996
rect 25130 25984 25136 25996
rect 25188 25984 25194 26036
rect 24854 25956 24860 25968
rect 22388 25928 23428 25956
rect 23492 25928 24860 25956
rect 12526 25848 12532 25900
rect 12584 25848 12590 25900
rect 22388 25897 22416 25928
rect 23492 25897 23520 25928
rect 24854 25916 24860 25928
rect 24912 25916 24918 25968
rect 15197 25891 15255 25897
rect 12820 25860 14228 25888
rect 11330 25780 11336 25832
rect 11388 25820 11394 25832
rect 12713 25823 12771 25829
rect 11388 25792 12572 25820
rect 11388 25780 11394 25792
rect 12544 25752 12572 25792
rect 12713 25789 12725 25823
rect 12759 25789 12771 25823
rect 12713 25783 12771 25789
rect 12728 25752 12756 25783
rect 12544 25724 12756 25752
rect 12161 25687 12219 25693
rect 12161 25653 12173 25687
rect 12207 25684 12219 25687
rect 12820 25684 12848 25860
rect 14090 25780 14096 25832
rect 14148 25780 14154 25832
rect 14200 25820 14228 25860
rect 15197 25857 15209 25891
rect 15243 25888 15255 25891
rect 16025 25891 16083 25897
rect 16025 25888 16037 25891
rect 15243 25860 16037 25888
rect 15243 25857 15255 25860
rect 15197 25851 15255 25857
rect 16025 25857 16037 25860
rect 16071 25857 16083 25891
rect 17037 25891 17095 25897
rect 17037 25888 17049 25891
rect 16025 25851 16083 25857
rect 16132 25860 17049 25888
rect 14200 25792 15332 25820
rect 13541 25755 13599 25761
rect 13541 25721 13553 25755
rect 13587 25752 13599 25755
rect 15304 25752 15332 25792
rect 15378 25780 15384 25832
rect 15436 25780 15442 25832
rect 16132 25752 16160 25860
rect 17037 25857 17049 25860
rect 17083 25857 17095 25891
rect 22373 25891 22431 25897
rect 22373 25888 22385 25891
rect 17037 25851 17095 25857
rect 21560 25860 22385 25888
rect 18417 25823 18475 25829
rect 18417 25789 18429 25823
rect 18463 25820 18475 25823
rect 18598 25820 18604 25832
rect 18463 25792 18604 25820
rect 18463 25789 18475 25792
rect 18417 25783 18475 25789
rect 18598 25780 18604 25792
rect 18656 25780 18662 25832
rect 17770 25752 17776 25764
rect 13587 25724 15240 25752
rect 15304 25724 16160 25752
rect 16500 25724 17776 25752
rect 13587 25721 13599 25724
rect 13541 25715 13599 25721
rect 12207 25656 12848 25684
rect 12207 25653 12219 25656
rect 12161 25647 12219 25653
rect 14826 25644 14832 25696
rect 14884 25684 14890 25696
rect 15010 25684 15016 25696
rect 14884 25656 15016 25684
rect 14884 25644 14890 25656
rect 15010 25644 15016 25656
rect 15068 25644 15074 25696
rect 15212 25684 15240 25724
rect 16500 25684 16528 25724
rect 17770 25712 17776 25724
rect 17828 25712 17834 25764
rect 15212 25656 16528 25684
rect 16850 25644 16856 25696
rect 16908 25644 16914 25696
rect 21174 25644 21180 25696
rect 21232 25684 21238 25696
rect 21560 25693 21588 25860
rect 22373 25857 22385 25860
rect 22419 25857 22431 25891
rect 22373 25851 22431 25857
rect 23477 25891 23535 25897
rect 23477 25857 23489 25891
rect 23523 25857 23535 25891
rect 23477 25851 23535 25857
rect 23934 25848 23940 25900
rect 23992 25848 23998 25900
rect 22649 25823 22707 25829
rect 22649 25789 22661 25823
rect 22695 25820 22707 25823
rect 23382 25820 23388 25832
rect 22695 25792 23388 25820
rect 22695 25789 22707 25792
rect 22649 25783 22707 25789
rect 23382 25780 23388 25792
rect 23440 25780 23446 25832
rect 25130 25780 25136 25832
rect 25188 25780 25194 25832
rect 22370 25712 22376 25764
rect 22428 25752 22434 25764
rect 22830 25752 22836 25764
rect 22428 25724 22836 25752
rect 22428 25712 22434 25724
rect 22830 25712 22836 25724
rect 22888 25712 22894 25764
rect 21545 25687 21603 25693
rect 21545 25684 21557 25687
rect 21232 25656 21557 25684
rect 21232 25644 21238 25656
rect 21545 25653 21557 25656
rect 21591 25653 21603 25687
rect 21545 25647 21603 25653
rect 21634 25644 21640 25696
rect 21692 25684 21698 25696
rect 22005 25687 22063 25693
rect 22005 25684 22017 25687
rect 21692 25656 22017 25684
rect 21692 25644 21698 25656
rect 22005 25653 22017 25656
rect 22051 25653 22063 25687
rect 22005 25647 22063 25653
rect 22462 25644 22468 25696
rect 22520 25684 22526 25696
rect 23293 25687 23351 25693
rect 23293 25684 23305 25687
rect 22520 25656 23305 25684
rect 22520 25644 22526 25656
rect 23293 25653 23305 25656
rect 23339 25653 23351 25687
rect 23293 25647 23351 25653
rect 1104 25594 25852 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 25852 25594
rect 1104 25520 25852 25542
rect 11698 25440 11704 25492
rect 11756 25480 11762 25492
rect 14277 25483 14335 25489
rect 14277 25480 14289 25483
rect 11756 25452 14289 25480
rect 11756 25440 11762 25452
rect 14277 25449 14289 25452
rect 14323 25449 14335 25483
rect 14277 25443 14335 25449
rect 16482 25440 16488 25492
rect 16540 25480 16546 25492
rect 18325 25483 18383 25489
rect 18325 25480 18337 25483
rect 16540 25452 18337 25480
rect 16540 25440 16546 25452
rect 18325 25449 18337 25452
rect 18371 25480 18383 25483
rect 18874 25480 18880 25492
rect 18371 25452 18880 25480
rect 18371 25449 18383 25452
rect 18325 25443 18383 25449
rect 18874 25440 18880 25452
rect 18932 25440 18938 25492
rect 20254 25440 20260 25492
rect 20312 25440 20318 25492
rect 21545 25483 21603 25489
rect 21545 25449 21557 25483
rect 21591 25480 21603 25483
rect 23934 25480 23940 25492
rect 21591 25452 23940 25480
rect 21591 25449 21603 25452
rect 21545 25443 21603 25449
rect 23934 25440 23940 25452
rect 23992 25440 23998 25492
rect 24026 25440 24032 25492
rect 24084 25480 24090 25492
rect 24581 25483 24639 25489
rect 24581 25480 24593 25483
rect 24084 25452 24593 25480
rect 24084 25440 24090 25452
rect 24581 25449 24593 25452
rect 24627 25449 24639 25483
rect 24581 25443 24639 25449
rect 12710 25372 12716 25424
rect 12768 25412 12774 25424
rect 12897 25415 12955 25421
rect 12897 25412 12909 25415
rect 12768 25384 12909 25412
rect 12768 25372 12774 25384
rect 12897 25381 12909 25384
rect 12943 25381 12955 25415
rect 12897 25375 12955 25381
rect 16945 25415 17003 25421
rect 16945 25381 16957 25415
rect 16991 25412 17003 25415
rect 24489 25415 24547 25421
rect 16991 25384 21772 25412
rect 16991 25381 17003 25384
rect 16945 25375 17003 25381
rect 10870 25304 10876 25356
rect 10928 25304 10934 25356
rect 11149 25347 11207 25353
rect 11149 25313 11161 25347
rect 11195 25344 11207 25347
rect 14550 25344 14556 25356
rect 11195 25316 14556 25344
rect 11195 25313 11207 25316
rect 11149 25307 11207 25313
rect 14550 25304 14556 25316
rect 14608 25304 14614 25356
rect 14642 25304 14648 25356
rect 14700 25344 14706 25356
rect 14737 25347 14795 25353
rect 14737 25344 14749 25347
rect 14700 25316 14749 25344
rect 14700 25304 14706 25316
rect 14737 25313 14749 25316
rect 14783 25313 14795 25347
rect 14737 25307 14795 25313
rect 14826 25304 14832 25356
rect 14884 25304 14890 25356
rect 16301 25347 16359 25353
rect 16301 25344 16313 25347
rect 14936 25316 16313 25344
rect 12710 25276 12716 25288
rect 12282 25248 12716 25276
rect 12710 25236 12716 25248
rect 12768 25236 12774 25288
rect 13354 25236 13360 25288
rect 13412 25276 13418 25288
rect 14936 25276 14964 25316
rect 16301 25313 16313 25316
rect 16347 25313 16359 25347
rect 16301 25307 16359 25313
rect 16850 25304 16856 25356
rect 16908 25344 16914 25356
rect 16908 25316 21036 25344
rect 16908 25304 16914 25316
rect 13412 25248 14964 25276
rect 13412 25236 13418 25248
rect 15194 25236 15200 25288
rect 15252 25276 15258 25288
rect 17129 25279 17187 25285
rect 17129 25276 17141 25279
rect 15252 25272 16804 25276
rect 16868 25272 17141 25276
rect 15252 25248 17141 25272
rect 15252 25236 15258 25248
rect 16776 25244 16896 25248
rect 17129 25245 17141 25248
rect 17175 25245 17187 25279
rect 17129 25239 17187 25245
rect 17770 25236 17776 25288
rect 17828 25236 17834 25288
rect 18141 25279 18199 25285
rect 18141 25245 18153 25279
rect 18187 25276 18199 25279
rect 18322 25276 18328 25288
rect 18187 25248 18328 25276
rect 18187 25245 18199 25248
rect 18141 25239 18199 25245
rect 18322 25236 18328 25248
rect 18380 25236 18386 25288
rect 19797 25279 19855 25285
rect 19797 25245 19809 25279
rect 19843 25276 19855 25279
rect 20254 25276 20260 25288
rect 19843 25248 20260 25276
rect 19843 25245 19855 25248
rect 19797 25239 19855 25245
rect 20254 25236 20260 25248
rect 20312 25236 20318 25288
rect 21008 25285 21036 25316
rect 21744 25285 21772 25384
rect 24489 25381 24501 25415
rect 24535 25412 24547 25415
rect 24854 25412 24860 25424
rect 24535 25384 24860 25412
rect 24535 25381 24547 25384
rect 24489 25375 24547 25381
rect 24854 25372 24860 25384
rect 24912 25372 24918 25424
rect 25133 25415 25191 25421
rect 25133 25381 25145 25415
rect 25179 25381 25191 25415
rect 25133 25375 25191 25381
rect 22370 25304 22376 25356
rect 22428 25344 22434 25356
rect 25148 25344 25176 25375
rect 22428 25316 25176 25344
rect 22428 25304 22434 25316
rect 20993 25279 21051 25285
rect 20993 25245 21005 25279
rect 21039 25245 21051 25279
rect 20993 25239 21051 25245
rect 21729 25279 21787 25285
rect 21729 25245 21741 25279
rect 21775 25245 21787 25279
rect 21729 25239 21787 25245
rect 22649 25279 22707 25285
rect 22649 25245 22661 25279
rect 22695 25245 22707 25279
rect 22649 25239 22707 25245
rect 15289 25211 15347 25217
rect 15289 25208 15301 25211
rect 12544 25180 15301 25208
rect 10318 25100 10324 25152
rect 10376 25140 10382 25152
rect 12544 25140 12572 25180
rect 15289 25177 15301 25180
rect 15335 25208 15347 25211
rect 15378 25208 15384 25220
rect 15335 25180 15384 25208
rect 15335 25177 15347 25180
rect 15289 25171 15347 25177
rect 15378 25168 15384 25180
rect 15436 25168 15442 25220
rect 16117 25211 16175 25217
rect 16117 25177 16129 25211
rect 16163 25208 16175 25211
rect 16390 25208 16396 25220
rect 16163 25180 16396 25208
rect 16163 25177 16175 25180
rect 16117 25171 16175 25177
rect 16390 25168 16396 25180
rect 16448 25168 16454 25220
rect 19058 25208 19064 25220
rect 17604 25180 19064 25208
rect 10376 25112 12572 25140
rect 10376 25100 10382 25112
rect 12618 25100 12624 25152
rect 12676 25100 12682 25152
rect 14645 25143 14703 25149
rect 14645 25109 14657 25143
rect 14691 25140 14703 25143
rect 15654 25140 15660 25152
rect 14691 25112 15660 25140
rect 14691 25109 14703 25112
rect 14645 25103 14703 25109
rect 15654 25100 15660 25112
rect 15712 25100 15718 25152
rect 15746 25100 15752 25152
rect 15804 25100 15810 25152
rect 16209 25143 16267 25149
rect 16209 25109 16221 25143
rect 16255 25140 16267 25143
rect 16482 25140 16488 25152
rect 16255 25112 16488 25140
rect 16255 25109 16267 25112
rect 16209 25103 16267 25109
rect 16482 25100 16488 25112
rect 16540 25100 16546 25152
rect 17604 25149 17632 25180
rect 19058 25168 19064 25180
rect 19116 25168 19122 25220
rect 19334 25168 19340 25220
rect 19392 25208 19398 25220
rect 20070 25208 20076 25220
rect 19392 25180 20076 25208
rect 19392 25168 19398 25180
rect 20070 25168 20076 25180
rect 20128 25168 20134 25220
rect 22664 25208 22692 25239
rect 25314 25236 25320 25288
rect 25372 25236 25378 25288
rect 20824 25180 22692 25208
rect 17589 25143 17647 25149
rect 17589 25109 17601 25143
rect 17635 25109 17647 25143
rect 17589 25103 17647 25109
rect 18506 25100 18512 25152
rect 18564 25140 18570 25152
rect 18693 25143 18751 25149
rect 18693 25140 18705 25143
rect 18564 25112 18705 25140
rect 18564 25100 18570 25112
rect 18693 25109 18705 25112
rect 18739 25109 18751 25143
rect 18693 25103 18751 25109
rect 19886 25100 19892 25152
rect 19944 25100 19950 25152
rect 20824 25149 20852 25180
rect 23842 25168 23848 25220
rect 23900 25168 23906 25220
rect 24857 25211 24915 25217
rect 24857 25177 24869 25211
rect 24903 25208 24915 25211
rect 26050 25208 26056 25220
rect 24903 25180 26056 25208
rect 24903 25177 24915 25180
rect 24857 25171 24915 25177
rect 25148 25152 25176 25180
rect 26050 25168 26056 25180
rect 26108 25168 26114 25220
rect 20809 25143 20867 25149
rect 20809 25109 20821 25143
rect 20855 25109 20867 25143
rect 20809 25103 20867 25109
rect 25130 25100 25136 25152
rect 25188 25100 25194 25152
rect 1104 25050 25852 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 25852 25050
rect 1104 24976 25852 24998
rect 7558 24896 7564 24948
rect 7616 24936 7622 24948
rect 7616 24908 11008 24936
rect 7616 24896 7622 24908
rect 9398 24828 9404 24880
rect 9456 24868 9462 24880
rect 10980 24868 11008 24908
rect 11146 24896 11152 24948
rect 11204 24936 11210 24948
rect 14826 24936 14832 24948
rect 11204 24908 14832 24936
rect 11204 24896 11210 24908
rect 14826 24896 14832 24908
rect 14884 24896 14890 24948
rect 15105 24939 15163 24945
rect 15105 24905 15117 24939
rect 15151 24936 15163 24939
rect 15654 24936 15660 24948
rect 15151 24908 15660 24936
rect 15151 24905 15163 24908
rect 15105 24899 15163 24905
rect 15654 24896 15660 24908
rect 15712 24896 15718 24948
rect 16390 24896 16396 24948
rect 16448 24936 16454 24948
rect 18322 24936 18328 24948
rect 16448 24908 18328 24936
rect 16448 24896 16454 24908
rect 18322 24896 18328 24908
rect 18380 24936 18386 24948
rect 18417 24939 18475 24945
rect 18417 24936 18429 24939
rect 18380 24908 18429 24936
rect 18380 24896 18386 24908
rect 18417 24905 18429 24908
rect 18463 24936 18475 24939
rect 18782 24936 18788 24948
rect 18463 24908 18788 24936
rect 18463 24905 18475 24908
rect 18417 24899 18475 24905
rect 18782 24896 18788 24908
rect 18840 24936 18846 24948
rect 19334 24936 19340 24948
rect 18840 24908 19340 24936
rect 18840 24896 18846 24908
rect 19334 24896 19340 24908
rect 19392 24896 19398 24948
rect 12069 24871 12127 24877
rect 12069 24868 12081 24871
rect 9456 24840 10166 24868
rect 10980 24840 12081 24868
rect 9456 24828 9462 24840
rect 12069 24837 12081 24840
rect 12115 24837 12127 24871
rect 12069 24831 12127 24837
rect 12710 24828 12716 24880
rect 12768 24868 12774 24880
rect 13538 24868 13544 24880
rect 12768 24840 13544 24868
rect 12768 24828 12774 24840
rect 13538 24828 13544 24840
rect 13596 24868 13602 24880
rect 13596 24840 13754 24868
rect 13596 24828 13602 24840
rect 14642 24828 14648 24880
rect 14700 24868 14706 24880
rect 15381 24871 15439 24877
rect 15381 24868 15393 24871
rect 14700 24840 15393 24868
rect 14700 24828 14706 24840
rect 15381 24837 15393 24840
rect 15427 24868 15439 24871
rect 15930 24868 15936 24880
rect 15427 24840 15936 24868
rect 15427 24837 15439 24840
rect 15381 24831 15439 24837
rect 15930 24828 15936 24840
rect 15988 24828 15994 24880
rect 17034 24828 17040 24880
rect 17092 24868 17098 24880
rect 17221 24871 17279 24877
rect 17221 24868 17233 24871
rect 17092 24840 17233 24868
rect 17092 24828 17098 24840
rect 17221 24837 17233 24840
rect 17267 24868 17279 24871
rect 18509 24871 18567 24877
rect 17267 24840 18000 24868
rect 17267 24837 17279 24840
rect 17221 24831 17279 24837
rect 12158 24760 12164 24812
rect 12216 24760 12222 24812
rect 12802 24760 12808 24812
rect 12860 24800 12866 24812
rect 12989 24803 13047 24809
rect 12989 24800 13001 24803
rect 12860 24772 13001 24800
rect 12860 24760 12866 24772
rect 12989 24769 13001 24772
rect 13035 24769 13047 24803
rect 15948 24800 15976 24828
rect 17313 24803 17371 24809
rect 17313 24800 17325 24803
rect 15948 24772 17325 24800
rect 12989 24763 13047 24769
rect 17313 24769 17325 24772
rect 17359 24800 17371 24803
rect 17972 24800 18000 24840
rect 18509 24837 18521 24871
rect 18555 24868 18567 24871
rect 18874 24868 18880 24880
rect 18555 24840 18880 24868
rect 18555 24837 18567 24840
rect 18509 24831 18567 24837
rect 18874 24828 18880 24840
rect 18932 24828 18938 24880
rect 22465 24871 22523 24877
rect 22465 24837 22477 24871
rect 22511 24868 22523 24871
rect 24118 24868 24124 24880
rect 22511 24840 24124 24868
rect 22511 24837 22523 24840
rect 22465 24831 22523 24837
rect 24118 24828 24124 24840
rect 24176 24828 24182 24880
rect 25130 24868 25136 24880
rect 25070 24840 25136 24868
rect 25130 24828 25136 24840
rect 25188 24828 25194 24880
rect 18322 24800 18328 24812
rect 17359 24772 17908 24800
rect 17972 24772 18328 24800
rect 17359 24769 17371 24772
rect 17313 24763 17371 24769
rect 9401 24735 9459 24741
rect 9401 24701 9413 24735
rect 9447 24701 9459 24735
rect 9401 24695 9459 24701
rect 9677 24735 9735 24741
rect 9677 24701 9689 24735
rect 9723 24732 9735 24735
rect 10870 24732 10876 24744
rect 9723 24704 10876 24732
rect 9723 24701 9735 24704
rect 9677 24695 9735 24701
rect 9416 24596 9444 24695
rect 10870 24692 10876 24704
rect 10928 24692 10934 24744
rect 11054 24692 11060 24744
rect 11112 24732 11118 24744
rect 12253 24735 12311 24741
rect 12253 24732 12265 24735
rect 11112 24704 12265 24732
rect 11112 24692 11118 24704
rect 12253 24701 12265 24704
rect 12299 24701 12311 24735
rect 12253 24695 12311 24701
rect 13265 24735 13323 24741
rect 13265 24701 13277 24735
rect 13311 24732 13323 24735
rect 13906 24732 13912 24744
rect 13311 24704 13912 24732
rect 13311 24701 13323 24704
rect 13265 24695 13323 24701
rect 13906 24692 13912 24704
rect 13964 24692 13970 24744
rect 14550 24692 14556 24744
rect 14608 24732 14614 24744
rect 14737 24735 14795 24741
rect 14737 24732 14749 24735
rect 14608 24704 14749 24732
rect 14608 24692 14614 24704
rect 14737 24701 14749 24704
rect 14783 24701 14795 24735
rect 14737 24695 14795 24701
rect 15010 24692 15016 24744
rect 15068 24732 15074 24744
rect 17405 24735 17463 24741
rect 17405 24732 17417 24735
rect 15068 24704 17417 24732
rect 15068 24692 15074 24704
rect 17405 24701 17417 24704
rect 17451 24701 17463 24735
rect 17880 24732 17908 24772
rect 18322 24760 18328 24772
rect 18380 24800 18386 24812
rect 19061 24803 19119 24809
rect 19061 24800 19073 24803
rect 18380 24772 19073 24800
rect 18380 24760 18386 24772
rect 19061 24769 19073 24772
rect 19107 24769 19119 24803
rect 19061 24763 19119 24769
rect 19426 24760 19432 24812
rect 19484 24800 19490 24812
rect 19705 24803 19763 24809
rect 19705 24800 19717 24803
rect 19484 24772 19717 24800
rect 19484 24760 19490 24772
rect 19705 24769 19717 24772
rect 19751 24769 19763 24803
rect 19705 24763 19763 24769
rect 21082 24760 21088 24812
rect 21140 24760 21146 24812
rect 23290 24760 23296 24812
rect 23348 24800 23354 24812
rect 23569 24803 23627 24809
rect 23569 24800 23581 24803
rect 23348 24772 23581 24800
rect 23348 24760 23354 24772
rect 23569 24769 23581 24772
rect 23615 24769 23627 24803
rect 23569 24763 23627 24769
rect 18138 24732 18144 24744
rect 17880 24704 18144 24732
rect 17405 24695 17463 24701
rect 18138 24692 18144 24704
rect 18196 24692 18202 24744
rect 18601 24735 18659 24741
rect 18601 24701 18613 24735
rect 18647 24701 18659 24735
rect 18601 24695 18659 24701
rect 19981 24735 20039 24741
rect 19981 24701 19993 24735
rect 20027 24732 20039 24735
rect 20438 24732 20444 24744
rect 20027 24704 20444 24732
rect 20027 24701 20039 24704
rect 19981 24695 20039 24701
rect 15194 24664 15200 24676
rect 14752 24636 15200 24664
rect 11054 24596 11060 24608
rect 9416 24568 11060 24596
rect 11054 24556 11060 24568
rect 11112 24556 11118 24608
rect 11146 24556 11152 24608
rect 11204 24556 11210 24608
rect 11701 24599 11759 24605
rect 11701 24565 11713 24599
rect 11747 24596 11759 24599
rect 14752 24596 14780 24636
rect 15194 24624 15200 24636
rect 15252 24624 15258 24676
rect 17034 24624 17040 24676
rect 17092 24664 17098 24676
rect 18616 24664 18644 24695
rect 20438 24692 20444 24704
rect 20496 24692 20502 24744
rect 21453 24735 21511 24741
rect 21453 24701 21465 24735
rect 21499 24732 21511 24735
rect 22278 24732 22284 24744
rect 21499 24704 22284 24732
rect 21499 24701 21511 24704
rect 21453 24695 21511 24701
rect 22278 24692 22284 24704
rect 22336 24692 22342 24744
rect 22557 24735 22615 24741
rect 22557 24701 22569 24735
rect 22603 24701 22615 24735
rect 22557 24695 22615 24701
rect 17092 24636 18644 24664
rect 22572 24664 22600 24695
rect 22646 24692 22652 24744
rect 22704 24692 22710 24744
rect 23845 24735 23903 24741
rect 23845 24701 23857 24735
rect 23891 24732 23903 24735
rect 25130 24732 25136 24744
rect 23891 24704 25136 24732
rect 23891 24701 23903 24704
rect 23845 24695 23903 24701
rect 25130 24692 25136 24704
rect 25188 24692 25194 24744
rect 23566 24664 23572 24676
rect 22572 24636 23572 24664
rect 17092 24624 17098 24636
rect 23566 24624 23572 24636
rect 23624 24624 23630 24676
rect 11747 24568 14780 24596
rect 11747 24565 11759 24568
rect 11701 24559 11759 24565
rect 15102 24556 15108 24608
rect 15160 24596 15166 24608
rect 15473 24599 15531 24605
rect 15473 24596 15485 24599
rect 15160 24568 15485 24596
rect 15160 24556 15166 24568
rect 15473 24565 15485 24568
rect 15519 24565 15531 24599
rect 15473 24559 15531 24565
rect 15562 24556 15568 24608
rect 15620 24596 15626 24608
rect 16853 24599 16911 24605
rect 16853 24596 16865 24599
rect 15620 24568 16865 24596
rect 15620 24556 15626 24568
rect 16853 24565 16865 24568
rect 16899 24565 16911 24599
rect 16853 24559 16911 24565
rect 17862 24556 17868 24608
rect 17920 24596 17926 24608
rect 18049 24599 18107 24605
rect 18049 24596 18061 24599
rect 17920 24568 18061 24596
rect 17920 24556 17926 24568
rect 18049 24565 18061 24568
rect 18095 24565 18107 24599
rect 18049 24559 18107 24565
rect 18138 24556 18144 24608
rect 18196 24596 18202 24608
rect 18690 24596 18696 24608
rect 18196 24568 18696 24596
rect 18196 24556 18202 24568
rect 18690 24556 18696 24568
rect 18748 24596 18754 24608
rect 19337 24599 19395 24605
rect 19337 24596 19349 24599
rect 18748 24568 19349 24596
rect 18748 24556 18754 24568
rect 19337 24565 19349 24568
rect 19383 24565 19395 24599
rect 19337 24559 19395 24565
rect 22094 24556 22100 24608
rect 22152 24556 22158 24608
rect 25222 24556 25228 24608
rect 25280 24596 25286 24608
rect 25317 24599 25375 24605
rect 25317 24596 25329 24599
rect 25280 24568 25329 24596
rect 25280 24556 25286 24568
rect 25317 24565 25329 24568
rect 25363 24596 25375 24599
rect 25406 24596 25412 24608
rect 25363 24568 25412 24596
rect 25363 24565 25375 24568
rect 25317 24559 25375 24565
rect 25406 24556 25412 24568
rect 25464 24556 25470 24608
rect 1104 24506 25852 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 25852 24506
rect 1104 24432 25852 24454
rect 12618 24392 12624 24404
rect 10428 24364 12624 24392
rect 9401 24259 9459 24265
rect 9401 24225 9413 24259
rect 9447 24256 9459 24259
rect 9490 24256 9496 24268
rect 9447 24228 9496 24256
rect 9447 24225 9459 24228
rect 9401 24219 9459 24225
rect 9490 24216 9496 24228
rect 9548 24256 9554 24268
rect 10428 24256 10456 24364
rect 12618 24352 12624 24364
rect 12676 24392 12682 24404
rect 12894 24392 12900 24404
rect 12676 24364 12900 24392
rect 12676 24352 12682 24364
rect 12894 24352 12900 24364
rect 12952 24352 12958 24404
rect 13538 24352 13544 24404
rect 13596 24392 13602 24404
rect 14185 24395 14243 24401
rect 14185 24392 14197 24395
rect 13596 24364 14197 24392
rect 13596 24352 13602 24364
rect 14185 24361 14197 24364
rect 14231 24392 14243 24395
rect 15102 24392 15108 24404
rect 14231 24364 15108 24392
rect 14231 24361 14243 24364
rect 14185 24355 14243 24361
rect 15102 24352 15108 24364
rect 15160 24352 15166 24404
rect 20438 24352 20444 24404
rect 20496 24392 20502 24404
rect 21177 24395 21235 24401
rect 21177 24392 21189 24395
rect 20496 24364 21189 24392
rect 20496 24352 20502 24364
rect 21177 24361 21189 24364
rect 21223 24361 21235 24395
rect 21177 24355 21235 24361
rect 25314 24352 25320 24404
rect 25372 24352 25378 24404
rect 25501 24395 25559 24401
rect 25501 24361 25513 24395
rect 25547 24392 25559 24395
rect 26050 24392 26056 24404
rect 25547 24364 26056 24392
rect 25547 24361 25559 24364
rect 25501 24355 25559 24361
rect 26050 24352 26056 24364
rect 26108 24352 26114 24404
rect 18141 24327 18199 24333
rect 18141 24293 18153 24327
rect 18187 24324 18199 24327
rect 19150 24324 19156 24336
rect 18187 24296 19156 24324
rect 18187 24293 18199 24296
rect 18141 24287 18199 24293
rect 19150 24284 19156 24296
rect 19208 24284 19214 24336
rect 21082 24284 21088 24336
rect 21140 24324 21146 24336
rect 21450 24324 21456 24336
rect 21140 24296 21456 24324
rect 21140 24284 21146 24296
rect 21450 24284 21456 24296
rect 21508 24324 21514 24336
rect 21545 24327 21603 24333
rect 21545 24324 21557 24327
rect 21508 24296 21557 24324
rect 21508 24284 21514 24296
rect 21545 24293 21557 24296
rect 21591 24293 21603 24327
rect 21545 24287 21603 24293
rect 23290 24284 23296 24336
rect 23348 24284 23354 24336
rect 25133 24327 25191 24333
rect 25133 24293 25145 24327
rect 25179 24324 25191 24327
rect 25406 24324 25412 24336
rect 25179 24296 25412 24324
rect 25179 24293 25191 24296
rect 25133 24287 25191 24293
rect 25406 24284 25412 24296
rect 25464 24324 25470 24336
rect 25958 24324 25964 24336
rect 25464 24296 25964 24324
rect 25464 24284 25470 24296
rect 25958 24284 25964 24296
rect 26016 24284 26022 24336
rect 9548 24228 10456 24256
rect 9548 24216 9554 24228
rect 11054 24216 11060 24268
rect 11112 24256 11118 24268
rect 11977 24259 12035 24265
rect 11977 24256 11989 24259
rect 11112 24228 11989 24256
rect 11112 24216 11118 24228
rect 11977 24225 11989 24228
rect 12023 24256 12035 24259
rect 12342 24256 12348 24268
rect 12023 24228 12348 24256
rect 12023 24225 12035 24228
rect 11977 24219 12035 24225
rect 12342 24216 12348 24228
rect 12400 24216 12406 24268
rect 18785 24259 18843 24265
rect 18785 24225 18797 24259
rect 18831 24256 18843 24259
rect 18966 24256 18972 24268
rect 18831 24228 18972 24256
rect 18831 24225 18843 24228
rect 18785 24219 18843 24225
rect 18966 24216 18972 24228
rect 19024 24216 19030 24268
rect 19426 24216 19432 24268
rect 19484 24216 19490 24268
rect 7834 24148 7840 24200
rect 7892 24188 7898 24200
rect 9125 24191 9183 24197
rect 9125 24188 9137 24191
rect 7892 24160 9137 24188
rect 7892 24148 7898 24160
rect 9125 24157 9137 24160
rect 9171 24157 9183 24191
rect 9125 24151 9183 24157
rect 17678 24148 17684 24200
rect 17736 24148 17742 24200
rect 18506 24148 18512 24200
rect 18564 24148 18570 24200
rect 18601 24191 18659 24197
rect 18601 24157 18613 24191
rect 18647 24188 18659 24191
rect 19242 24188 19248 24200
rect 18647 24160 19248 24188
rect 18647 24157 18659 24160
rect 18601 24151 18659 24157
rect 19242 24148 19248 24160
rect 19300 24148 19306 24200
rect 21100 24188 21128 24284
rect 21913 24259 21971 24265
rect 21913 24225 21925 24259
rect 21959 24256 21971 24259
rect 22186 24256 22192 24268
rect 21959 24228 22192 24256
rect 21959 24225 21971 24228
rect 21913 24219 21971 24225
rect 22186 24216 22192 24228
rect 22244 24256 22250 24268
rect 23308 24256 23336 24284
rect 22244 24228 23336 24256
rect 22244 24216 22250 24228
rect 24118 24216 24124 24268
rect 24176 24256 24182 24268
rect 24581 24259 24639 24265
rect 24581 24256 24593 24259
rect 24176 24228 24593 24256
rect 24176 24216 24182 24228
rect 24581 24225 24593 24228
rect 24627 24225 24639 24259
rect 24581 24219 24639 24225
rect 20838 24160 21128 24188
rect 9398 24080 9404 24132
rect 9456 24120 9462 24132
rect 11241 24123 11299 24129
rect 11241 24120 11253 24123
rect 9456 24092 9890 24120
rect 10704 24092 11253 24120
rect 9456 24080 9462 24092
rect 9784 24052 9812 24092
rect 10704 24052 10732 24092
rect 11241 24089 11253 24092
rect 11287 24120 11299 24123
rect 11425 24123 11483 24129
rect 11425 24120 11437 24123
rect 11287 24092 11437 24120
rect 11287 24089 11299 24092
rect 11241 24083 11299 24089
rect 11425 24089 11437 24092
rect 11471 24089 11483 24123
rect 11425 24083 11483 24089
rect 9784 24024 10732 24052
rect 10870 24012 10876 24064
rect 10928 24012 10934 24064
rect 11440 24052 11468 24083
rect 11974 24080 11980 24132
rect 12032 24120 12038 24132
rect 12253 24123 12311 24129
rect 12253 24120 12265 24123
rect 12032 24092 12265 24120
rect 12032 24080 12038 24092
rect 12253 24089 12265 24092
rect 12299 24089 12311 24123
rect 12710 24120 12716 24132
rect 12253 24083 12311 24089
rect 12406 24092 12716 24120
rect 12406 24052 12434 24092
rect 12710 24080 12716 24092
rect 12768 24080 12774 24132
rect 15933 24123 15991 24129
rect 15933 24089 15945 24123
rect 15979 24120 15991 24123
rect 18874 24120 18880 24132
rect 15979 24092 18880 24120
rect 15979 24089 15991 24092
rect 15933 24083 15991 24089
rect 18874 24080 18880 24092
rect 18932 24080 18938 24132
rect 19705 24123 19763 24129
rect 19705 24089 19717 24123
rect 19751 24089 19763 24123
rect 19705 24083 19763 24089
rect 22189 24123 22247 24129
rect 22189 24089 22201 24123
rect 22235 24120 22247 24123
rect 22278 24120 22284 24132
rect 22235 24092 22284 24120
rect 22235 24089 22247 24092
rect 22189 24083 22247 24089
rect 11440 24024 12434 24052
rect 13725 24055 13783 24061
rect 13725 24021 13737 24055
rect 13771 24052 13783 24055
rect 13906 24052 13912 24064
rect 13771 24024 13912 24052
rect 13771 24021 13783 24024
rect 13725 24015 13783 24021
rect 13906 24012 13912 24024
rect 13964 24012 13970 24064
rect 16574 24012 16580 24064
rect 16632 24052 16638 24064
rect 18782 24052 18788 24064
rect 16632 24024 18788 24052
rect 16632 24012 16638 24024
rect 18782 24012 18788 24024
rect 18840 24012 18846 24064
rect 19720 24052 19748 24083
rect 22278 24080 22284 24092
rect 22336 24080 22342 24132
rect 23414 24092 24072 24120
rect 19886 24052 19892 24064
rect 19720 24024 19892 24052
rect 19886 24012 19892 24024
rect 19944 24012 19950 24064
rect 23566 24012 23572 24064
rect 23624 24052 23630 24064
rect 24044 24061 24072 24092
rect 23661 24055 23719 24061
rect 23661 24052 23673 24055
rect 23624 24024 23673 24052
rect 23624 24012 23630 24024
rect 23661 24021 23673 24024
rect 23707 24021 23719 24055
rect 23661 24015 23719 24021
rect 24029 24055 24087 24061
rect 24029 24021 24041 24055
rect 24075 24052 24087 24055
rect 24946 24052 24952 24064
rect 24075 24024 24952 24052
rect 24075 24021 24087 24024
rect 24029 24015 24087 24021
rect 24946 24012 24952 24024
rect 25004 24012 25010 24064
rect 1104 23962 25852 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 25852 23962
rect 1104 23888 25852 23910
rect 9674 23808 9680 23860
rect 9732 23848 9738 23860
rect 9769 23851 9827 23857
rect 9769 23848 9781 23851
rect 9732 23820 9781 23848
rect 9732 23808 9738 23820
rect 9769 23817 9781 23820
rect 9815 23817 9827 23851
rect 9769 23811 9827 23817
rect 7834 23672 7840 23724
rect 7892 23712 7898 23724
rect 8021 23715 8079 23721
rect 8021 23712 8033 23715
rect 7892 23684 8033 23712
rect 7892 23672 7898 23684
rect 8021 23681 8033 23684
rect 8067 23681 8079 23715
rect 8021 23675 8079 23681
rect 9398 23672 9404 23724
rect 9456 23672 9462 23724
rect 9784 23712 9812 23811
rect 10410 23808 10416 23860
rect 10468 23808 10474 23860
rect 10781 23851 10839 23857
rect 10781 23817 10793 23851
rect 10827 23848 10839 23851
rect 14182 23848 14188 23860
rect 10827 23820 14188 23848
rect 10827 23817 10839 23820
rect 10781 23811 10839 23817
rect 14182 23808 14188 23820
rect 14240 23808 14246 23860
rect 14918 23808 14924 23860
rect 14976 23808 14982 23860
rect 16574 23808 16580 23860
rect 16632 23848 16638 23860
rect 17221 23851 17279 23857
rect 17221 23848 17233 23851
rect 16632 23820 17233 23848
rect 16632 23808 16638 23820
rect 17221 23817 17233 23820
rect 17267 23817 17279 23851
rect 17221 23811 17279 23817
rect 17313 23851 17371 23857
rect 17313 23817 17325 23851
rect 17359 23848 17371 23851
rect 17770 23848 17776 23860
rect 17359 23820 17776 23848
rect 17359 23817 17371 23820
rect 17313 23811 17371 23817
rect 17770 23808 17776 23820
rect 17828 23808 17834 23860
rect 18049 23851 18107 23857
rect 18049 23817 18061 23851
rect 18095 23817 18107 23851
rect 18049 23811 18107 23817
rect 18601 23851 18659 23857
rect 18601 23817 18613 23851
rect 18647 23848 18659 23851
rect 18782 23848 18788 23860
rect 18647 23820 18788 23848
rect 18647 23817 18659 23820
rect 18601 23811 18659 23817
rect 13630 23740 13636 23792
rect 13688 23740 13694 23792
rect 13722 23740 13728 23792
rect 13780 23740 13786 23792
rect 15838 23740 15844 23792
rect 15896 23780 15902 23792
rect 18064 23780 18092 23811
rect 18782 23808 18788 23820
rect 18840 23808 18846 23860
rect 18874 23808 18880 23860
rect 18932 23808 18938 23860
rect 19058 23808 19064 23860
rect 19116 23848 19122 23860
rect 24949 23851 25007 23857
rect 19116 23820 22094 23848
rect 19116 23808 19122 23820
rect 22066 23780 22094 23820
rect 24949 23817 24961 23851
rect 24995 23848 25007 23851
rect 25130 23848 25136 23860
rect 24995 23820 25136 23848
rect 24995 23817 25007 23820
rect 24949 23811 25007 23817
rect 25130 23808 25136 23820
rect 25188 23808 25194 23860
rect 25406 23808 25412 23860
rect 25464 23808 25470 23860
rect 23382 23780 23388 23792
rect 15896 23752 17448 23780
rect 18064 23752 21956 23780
rect 22066 23752 22416 23780
rect 15896 23740 15902 23752
rect 9784 23684 11008 23712
rect 10980 23656 11008 23684
rect 13998 23672 14004 23724
rect 14056 23712 14062 23724
rect 14829 23715 14887 23721
rect 14829 23712 14841 23715
rect 14056 23684 14841 23712
rect 14056 23672 14062 23684
rect 14829 23681 14841 23684
rect 14875 23681 14887 23715
rect 14829 23675 14887 23681
rect 8297 23647 8355 23653
rect 8297 23613 8309 23647
rect 8343 23644 8355 23647
rect 8343 23616 9996 23644
rect 8343 23613 8355 23616
rect 8297 23607 8355 23613
rect 9968 23576 9996 23616
rect 10042 23604 10048 23656
rect 10100 23644 10106 23656
rect 10873 23647 10931 23653
rect 10873 23644 10885 23647
rect 10100 23616 10885 23644
rect 10100 23604 10106 23616
rect 10873 23613 10885 23616
rect 10919 23613 10931 23647
rect 10873 23607 10931 23613
rect 10962 23604 10968 23656
rect 11020 23604 11026 23656
rect 13817 23647 13875 23653
rect 13817 23613 13829 23647
rect 13863 23613 13875 23647
rect 13817 23607 13875 23613
rect 10318 23576 10324 23588
rect 9968 23548 10324 23576
rect 10318 23536 10324 23548
rect 10376 23536 10382 23588
rect 12894 23536 12900 23588
rect 12952 23576 12958 23588
rect 13832 23576 13860 23607
rect 13906 23604 13912 23656
rect 13964 23644 13970 23656
rect 15013 23647 15071 23653
rect 15013 23644 15025 23647
rect 13964 23616 15025 23644
rect 13964 23604 13970 23616
rect 15013 23613 15025 23616
rect 15059 23613 15071 23647
rect 15013 23607 15071 23613
rect 15654 23604 15660 23656
rect 15712 23604 15718 23656
rect 17420 23653 17448 23752
rect 18233 23715 18291 23721
rect 18233 23681 18245 23715
rect 18279 23681 18291 23715
rect 18233 23675 18291 23681
rect 17405 23647 17463 23653
rect 17405 23613 17417 23647
rect 17451 23613 17463 23647
rect 17405 23607 17463 23613
rect 12952 23548 13860 23576
rect 14461 23579 14519 23585
rect 12952 23536 12958 23548
rect 14461 23545 14473 23579
rect 14507 23576 14519 23579
rect 18248 23576 18276 23675
rect 19610 23672 19616 23724
rect 19668 23672 19674 23724
rect 19705 23715 19763 23721
rect 19705 23681 19717 23715
rect 19751 23712 19763 23715
rect 20346 23712 20352 23724
rect 19751 23684 20352 23712
rect 19751 23681 19763 23684
rect 19705 23675 19763 23681
rect 19518 23604 19524 23656
rect 19576 23644 19582 23656
rect 19720 23644 19748 23675
rect 20346 23672 20352 23684
rect 20404 23672 20410 23724
rect 20806 23672 20812 23724
rect 20864 23672 20870 23724
rect 20901 23715 20959 23721
rect 20901 23681 20913 23715
rect 20947 23712 20959 23715
rect 21358 23712 21364 23724
rect 20947 23684 21364 23712
rect 20947 23681 20959 23684
rect 20901 23675 20959 23681
rect 21358 23672 21364 23684
rect 21416 23672 21422 23724
rect 21450 23672 21456 23724
rect 21508 23672 21514 23724
rect 21928 23712 21956 23752
rect 22002 23712 22008 23724
rect 21928 23684 22008 23712
rect 22002 23672 22008 23684
rect 22060 23672 22066 23724
rect 22388 23721 22416 23752
rect 22480 23752 23388 23780
rect 22373 23715 22431 23721
rect 22373 23681 22385 23715
rect 22419 23681 22431 23715
rect 22373 23675 22431 23681
rect 19576 23616 19748 23644
rect 19576 23604 19582 23616
rect 19886 23604 19892 23656
rect 19944 23604 19950 23656
rect 20990 23604 20996 23656
rect 21048 23604 21054 23656
rect 22480 23644 22508 23752
rect 23382 23740 23388 23752
rect 23440 23740 23446 23792
rect 25317 23783 25375 23789
rect 25317 23780 25329 23783
rect 24702 23752 25329 23780
rect 24964 23724 24992 23752
rect 25317 23749 25329 23752
rect 25363 23780 25375 23783
rect 26050 23780 26056 23792
rect 25363 23752 26056 23780
rect 25363 23749 25375 23752
rect 25317 23743 25375 23749
rect 26050 23740 26056 23752
rect 26108 23740 26114 23792
rect 23198 23672 23204 23724
rect 23256 23672 23262 23724
rect 24946 23672 24952 23724
rect 25004 23672 25010 23724
rect 21100 23616 22508 23644
rect 23477 23647 23535 23653
rect 14507 23548 18276 23576
rect 19904 23576 19932 23604
rect 21100 23576 21128 23616
rect 23477 23613 23489 23647
rect 23523 23644 23535 23647
rect 23566 23644 23572 23656
rect 23523 23616 23572 23644
rect 23523 23613 23535 23616
rect 23477 23607 23535 23613
rect 23566 23604 23572 23616
rect 23624 23604 23630 23656
rect 19904 23548 21128 23576
rect 14507 23545 14519 23548
rect 14461 23539 14519 23545
rect 22094 23536 22100 23588
rect 22152 23576 22158 23588
rect 22278 23576 22284 23588
rect 22152 23548 22284 23576
rect 22152 23536 22158 23548
rect 22278 23536 22284 23548
rect 22336 23536 22342 23588
rect 9398 23468 9404 23520
rect 9456 23508 9462 23520
rect 10045 23511 10103 23517
rect 10045 23508 10057 23511
rect 9456 23480 10057 23508
rect 9456 23468 9462 23480
rect 10045 23477 10057 23480
rect 10091 23477 10103 23511
rect 10045 23471 10103 23477
rect 10870 23468 10876 23520
rect 10928 23508 10934 23520
rect 12618 23508 12624 23520
rect 10928 23480 12624 23508
rect 10928 23468 10934 23480
rect 12618 23468 12624 23480
rect 12676 23468 12682 23520
rect 12802 23468 12808 23520
rect 12860 23508 12866 23520
rect 13265 23511 13323 23517
rect 13265 23508 13277 23511
rect 12860 23480 13277 23508
rect 12860 23468 12866 23480
rect 13265 23477 13277 23480
rect 13311 23477 13323 23511
rect 13265 23471 13323 23477
rect 16853 23511 16911 23517
rect 16853 23477 16865 23511
rect 16899 23508 16911 23511
rect 17310 23508 17316 23520
rect 16899 23480 17316 23508
rect 16899 23477 16911 23480
rect 16853 23471 16911 23477
rect 17310 23468 17316 23480
rect 17368 23468 17374 23520
rect 17770 23468 17776 23520
rect 17828 23508 17834 23520
rect 18785 23511 18843 23517
rect 18785 23508 18797 23511
rect 17828 23480 18797 23508
rect 17828 23468 17834 23480
rect 18785 23477 18797 23480
rect 18831 23508 18843 23511
rect 19058 23508 19064 23520
rect 18831 23480 19064 23508
rect 18831 23477 18843 23480
rect 18785 23471 18843 23477
rect 19058 23468 19064 23480
rect 19116 23468 19122 23520
rect 19242 23468 19248 23520
rect 19300 23468 19306 23520
rect 19334 23468 19340 23520
rect 19392 23508 19398 23520
rect 20441 23511 20499 23517
rect 20441 23508 20453 23511
rect 19392 23480 20453 23508
rect 19392 23468 19398 23480
rect 20441 23477 20453 23480
rect 20487 23477 20499 23511
rect 20441 23471 20499 23477
rect 22189 23511 22247 23517
rect 22189 23477 22201 23511
rect 22235 23508 22247 23511
rect 23934 23508 23940 23520
rect 22235 23480 23940 23508
rect 22235 23477 22247 23480
rect 22189 23471 22247 23477
rect 23934 23468 23940 23480
rect 23992 23468 23998 23520
rect 1104 23418 25852 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 25852 23418
rect 1104 23344 25852 23366
rect 9125 23307 9183 23313
rect 9125 23273 9137 23307
rect 9171 23304 9183 23307
rect 9214 23304 9220 23316
rect 9171 23276 9220 23304
rect 9171 23273 9183 23276
rect 9125 23267 9183 23273
rect 9214 23264 9220 23276
rect 9272 23264 9278 23316
rect 10134 23264 10140 23316
rect 10192 23304 10198 23316
rect 15194 23304 15200 23316
rect 10192 23276 15200 23304
rect 10192 23264 10198 23276
rect 15194 23264 15200 23276
rect 15252 23264 15258 23316
rect 15841 23307 15899 23313
rect 15841 23273 15853 23307
rect 15887 23304 15899 23307
rect 17126 23304 17132 23316
rect 15887 23276 17132 23304
rect 15887 23273 15899 23276
rect 15841 23267 15899 23273
rect 9398 23196 9404 23248
rect 9456 23236 9462 23248
rect 9456 23208 12434 23236
rect 9456 23196 9462 23208
rect 8662 23128 8668 23180
rect 8720 23168 8726 23180
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 8720 23140 9689 23168
rect 8720 23128 8726 23140
rect 9677 23137 9689 23140
rect 9723 23137 9735 23171
rect 9677 23131 9735 23137
rect 10229 23171 10287 23177
rect 10229 23137 10241 23171
rect 10275 23168 10287 23171
rect 10318 23168 10324 23180
rect 10275 23140 10324 23168
rect 10275 23137 10287 23140
rect 10229 23131 10287 23137
rect 10318 23128 10324 23140
rect 10376 23168 10382 23180
rect 10594 23168 10600 23180
rect 10376 23140 10600 23168
rect 10376 23128 10382 23140
rect 10594 23128 10600 23140
rect 10652 23128 10658 23180
rect 11698 23128 11704 23180
rect 11756 23128 11762 23180
rect 11790 23128 11796 23180
rect 11848 23128 11854 23180
rect 12406 23168 12434 23208
rect 12710 23196 12716 23248
rect 12768 23236 12774 23248
rect 14737 23239 14795 23245
rect 14737 23236 14749 23239
rect 12768 23208 14749 23236
rect 12768 23196 12774 23208
rect 14737 23205 14749 23208
rect 14783 23205 14795 23239
rect 14737 23199 14795 23205
rect 13541 23171 13599 23177
rect 13541 23168 13553 23171
rect 12406 23140 13553 23168
rect 13541 23137 13553 23140
rect 13587 23137 13599 23171
rect 15289 23171 15347 23177
rect 15289 23168 15301 23171
rect 13541 23131 13599 23137
rect 14476 23140 15301 23168
rect 9585 23103 9643 23109
rect 9585 23069 9597 23103
rect 9631 23100 9643 23103
rect 10778 23100 10784 23112
rect 9631 23072 10784 23100
rect 9631 23069 9643 23072
rect 9585 23063 9643 23069
rect 10778 23060 10784 23072
rect 10836 23060 10842 23112
rect 11606 23060 11612 23112
rect 11664 23060 11670 23112
rect 13357 23103 13415 23109
rect 13357 23069 13369 23103
rect 13403 23100 13415 23103
rect 14182 23100 14188 23112
rect 13403 23072 14188 23100
rect 13403 23069 13415 23072
rect 13357 23063 13415 23069
rect 14182 23060 14188 23072
rect 14240 23060 14246 23112
rect 9493 23035 9551 23041
rect 9493 23001 9505 23035
rect 9539 23032 9551 23035
rect 10410 23032 10416 23044
rect 9539 23004 10416 23032
rect 9539 23001 9551 23004
rect 9493 22995 9551 23001
rect 10410 22992 10416 23004
rect 10468 22992 10474 23044
rect 14090 22992 14096 23044
rect 14148 23032 14154 23044
rect 14476 23041 14504 23140
rect 15289 23137 15301 23140
rect 15335 23137 15347 23171
rect 15289 23131 15347 23137
rect 15105 23103 15163 23109
rect 15105 23069 15117 23103
rect 15151 23100 15163 23103
rect 15654 23100 15660 23112
rect 15151 23072 15660 23100
rect 15151 23069 15163 23072
rect 15105 23063 15163 23069
rect 15654 23060 15660 23072
rect 15712 23060 15718 23112
rect 14461 23035 14519 23041
rect 14461 23032 14473 23035
rect 14148 23004 14473 23032
rect 14148 22992 14154 23004
rect 14461 23001 14473 23004
rect 14507 23001 14519 23035
rect 14461 22995 14519 23001
rect 15197 23035 15255 23041
rect 15197 23001 15209 23035
rect 15243 23032 15255 23035
rect 15856 23032 15884 23267
rect 17126 23264 17132 23276
rect 17184 23264 17190 23316
rect 18969 23307 19027 23313
rect 18969 23273 18981 23307
rect 19015 23304 19027 23307
rect 19518 23304 19524 23316
rect 19015 23276 19524 23304
rect 19015 23273 19027 23276
rect 18969 23267 19027 23273
rect 19518 23264 19524 23276
rect 19576 23264 19582 23316
rect 17865 23239 17923 23245
rect 17865 23205 17877 23239
rect 17911 23236 17923 23239
rect 18874 23236 18880 23248
rect 17911 23208 18880 23236
rect 17911 23205 17923 23208
rect 17865 23199 17923 23205
rect 18874 23196 18880 23208
rect 18932 23196 18938 23248
rect 25866 23236 25872 23248
rect 25056 23208 25872 23236
rect 18414 23128 18420 23180
rect 18472 23128 18478 23180
rect 20165 23171 20223 23177
rect 20165 23137 20177 23171
rect 20211 23168 20223 23171
rect 20438 23168 20444 23180
rect 20211 23140 20444 23168
rect 20211 23137 20223 23140
rect 20165 23131 20223 23137
rect 20438 23128 20444 23140
rect 20496 23128 20502 23180
rect 20717 23171 20775 23177
rect 20717 23137 20729 23171
rect 20763 23168 20775 23171
rect 20806 23168 20812 23180
rect 20763 23140 20812 23168
rect 20763 23137 20775 23140
rect 20717 23131 20775 23137
rect 20806 23128 20812 23140
rect 20864 23128 20870 23180
rect 25056 23177 25084 23208
rect 25866 23196 25872 23208
rect 25924 23196 25930 23248
rect 25041 23171 25099 23177
rect 25041 23137 25053 23171
rect 25087 23137 25099 23171
rect 25041 23131 25099 23137
rect 25225 23171 25283 23177
rect 25225 23137 25237 23171
rect 25271 23168 25283 23171
rect 25314 23168 25320 23180
rect 25271 23140 25320 23168
rect 25271 23137 25283 23140
rect 25225 23131 25283 23137
rect 25314 23128 25320 23140
rect 25372 23128 25378 23180
rect 18233 23103 18291 23109
rect 18233 23069 18245 23103
rect 18279 23100 18291 23103
rect 18322 23100 18328 23112
rect 18279 23072 18328 23100
rect 18279 23069 18291 23072
rect 18233 23063 18291 23069
rect 18322 23060 18328 23072
rect 18380 23060 18386 23112
rect 19242 23060 19248 23112
rect 19300 23100 19306 23112
rect 19889 23103 19947 23109
rect 19889 23100 19901 23103
rect 19300 23072 19901 23100
rect 19300 23060 19306 23072
rect 19889 23069 19901 23072
rect 19935 23069 19947 23103
rect 19889 23063 19947 23069
rect 19981 23103 20039 23109
rect 19981 23069 19993 23103
rect 20027 23100 20039 23103
rect 21634 23100 21640 23112
rect 20027 23072 21640 23100
rect 20027 23069 20039 23072
rect 19981 23063 20039 23069
rect 21634 23060 21640 23072
rect 21692 23060 21698 23112
rect 21821 23103 21879 23109
rect 21821 23069 21833 23103
rect 21867 23069 21879 23103
rect 21821 23063 21879 23069
rect 22833 23103 22891 23109
rect 22833 23069 22845 23103
rect 22879 23100 22891 23103
rect 23750 23100 23756 23112
rect 22879 23072 23756 23100
rect 22879 23069 22891 23072
rect 22833 23063 22891 23069
rect 15243 23004 15884 23032
rect 15243 23001 15255 23004
rect 15197 22995 15255 23001
rect 16850 22992 16856 23044
rect 16908 23032 16914 23044
rect 21836 23032 21864 23063
rect 23750 23060 23756 23072
rect 23808 23060 23814 23112
rect 24949 23103 25007 23109
rect 24949 23069 24961 23103
rect 24995 23100 25007 23103
rect 25406 23100 25412 23112
rect 24995 23072 25412 23100
rect 24995 23069 25007 23072
rect 24949 23063 25007 23069
rect 25406 23060 25412 23072
rect 25464 23060 25470 23112
rect 16908 23004 21864 23032
rect 23845 23035 23903 23041
rect 16908 22992 16914 23004
rect 23845 23001 23857 23035
rect 23891 23032 23903 23035
rect 25866 23032 25872 23044
rect 23891 23004 25872 23032
rect 23891 23001 23903 23004
rect 23845 22995 23903 23001
rect 25866 22992 25872 23004
rect 25924 22992 25930 23044
rect 10502 22924 10508 22976
rect 10560 22964 10566 22976
rect 11241 22967 11299 22973
rect 11241 22964 11253 22967
rect 10560 22936 11253 22964
rect 10560 22924 10566 22936
rect 11241 22933 11253 22936
rect 11287 22933 11299 22967
rect 11241 22927 11299 22933
rect 12158 22924 12164 22976
rect 12216 22964 12222 22976
rect 12989 22967 13047 22973
rect 12989 22964 13001 22967
rect 12216 22936 13001 22964
rect 12216 22924 12222 22936
rect 12989 22933 13001 22936
rect 13035 22933 13047 22967
rect 12989 22927 13047 22933
rect 13449 22967 13507 22973
rect 13449 22933 13461 22967
rect 13495 22964 13507 22967
rect 14185 22967 14243 22973
rect 14185 22964 14197 22967
rect 13495 22936 14197 22964
rect 13495 22933 13507 22936
rect 13449 22927 13507 22933
rect 14185 22933 14197 22936
rect 14231 22964 14243 22967
rect 17770 22964 17776 22976
rect 14231 22936 17776 22964
rect 14231 22933 14243 22936
rect 14185 22927 14243 22933
rect 17770 22924 17776 22936
rect 17828 22924 17834 22976
rect 18325 22967 18383 22973
rect 18325 22933 18337 22967
rect 18371 22964 18383 22967
rect 18690 22964 18696 22976
rect 18371 22936 18696 22964
rect 18371 22933 18383 22936
rect 18325 22927 18383 22933
rect 18690 22924 18696 22936
rect 18748 22924 18754 22976
rect 18966 22924 18972 22976
rect 19024 22964 19030 22976
rect 19521 22967 19579 22973
rect 19521 22964 19533 22967
rect 19024 22936 19533 22964
rect 19024 22924 19030 22936
rect 19521 22933 19533 22936
rect 19567 22933 19579 22967
rect 19521 22927 19579 22933
rect 21637 22967 21695 22973
rect 21637 22933 21649 22967
rect 21683 22964 21695 22967
rect 22094 22964 22100 22976
rect 21683 22936 22100 22964
rect 21683 22933 21695 22936
rect 21637 22927 21695 22933
rect 22094 22924 22100 22936
rect 22152 22924 22158 22976
rect 24578 22924 24584 22976
rect 24636 22924 24642 22976
rect 1104 22874 25852 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 25852 22874
rect 1104 22800 25852 22822
rect 11330 22720 11336 22772
rect 11388 22760 11394 22772
rect 14090 22760 14096 22772
rect 11388 22732 14096 22760
rect 11388 22720 11394 22732
rect 14090 22720 14096 22732
rect 14148 22720 14154 22772
rect 14182 22720 14188 22772
rect 14240 22760 14246 22772
rect 14461 22763 14519 22769
rect 14461 22760 14473 22763
rect 14240 22732 14473 22760
rect 14240 22720 14246 22732
rect 14461 22729 14473 22732
rect 14507 22760 14519 22763
rect 14734 22760 14740 22772
rect 14507 22732 14740 22760
rect 14507 22729 14519 22732
rect 14461 22723 14519 22729
rect 14734 22720 14740 22732
rect 14792 22720 14798 22772
rect 16850 22720 16856 22772
rect 16908 22720 16914 22772
rect 18322 22720 18328 22772
rect 18380 22760 18386 22772
rect 18693 22763 18751 22769
rect 18693 22760 18705 22763
rect 18380 22732 18705 22760
rect 18380 22720 18386 22732
rect 18693 22729 18705 22732
rect 18739 22729 18751 22763
rect 18693 22723 18751 22729
rect 14553 22695 14611 22701
rect 14553 22692 14565 22695
rect 13846 22664 14565 22692
rect 14553 22661 14565 22664
rect 14599 22692 14611 22695
rect 15102 22692 15108 22704
rect 14599 22664 15108 22692
rect 14599 22661 14611 22664
rect 14553 22655 14611 22661
rect 15102 22652 15108 22664
rect 15160 22652 15166 22704
rect 18708 22692 18736 22723
rect 19058 22720 19064 22772
rect 19116 22760 19122 22772
rect 19242 22760 19248 22772
rect 19116 22732 19248 22760
rect 19116 22720 19122 22732
rect 19242 22720 19248 22732
rect 19300 22720 19306 22772
rect 19610 22720 19616 22772
rect 19668 22760 19674 22772
rect 19705 22763 19763 22769
rect 19705 22760 19717 22763
rect 19668 22732 19717 22760
rect 19668 22720 19674 22732
rect 19705 22729 19717 22732
rect 19751 22729 19763 22763
rect 19705 22723 19763 22729
rect 21177 22763 21235 22769
rect 21177 22729 21189 22763
rect 21223 22760 21235 22763
rect 22370 22760 22376 22772
rect 21223 22732 22376 22760
rect 21223 22729 21235 22732
rect 21177 22723 21235 22729
rect 22370 22720 22376 22732
rect 22428 22720 22434 22772
rect 20806 22692 20812 22704
rect 18708 22664 20812 22692
rect 20806 22652 20812 22664
rect 20864 22652 20870 22704
rect 7834 22584 7840 22636
rect 7892 22624 7898 22636
rect 8113 22627 8171 22633
rect 8113 22624 8125 22627
rect 7892 22596 8125 22624
rect 7892 22584 7898 22596
rect 8113 22593 8125 22596
rect 8159 22593 8171 22627
rect 8113 22587 8171 22593
rect 9490 22584 9496 22636
rect 9548 22624 9554 22636
rect 10137 22627 10195 22633
rect 10137 22624 10149 22627
rect 9548 22596 10149 22624
rect 9548 22584 9554 22596
rect 10137 22593 10149 22596
rect 10183 22593 10195 22627
rect 10137 22587 10195 22593
rect 12342 22584 12348 22636
rect 12400 22584 12406 22636
rect 13906 22584 13912 22636
rect 13964 22624 13970 22636
rect 17037 22627 17095 22633
rect 17037 22624 17049 22627
rect 13964 22596 17049 22624
rect 13964 22584 13970 22596
rect 17037 22593 17049 22596
rect 17083 22593 17095 22627
rect 17037 22587 17095 22593
rect 18690 22584 18696 22636
rect 18748 22624 18754 22636
rect 18877 22627 18935 22633
rect 18877 22624 18889 22627
rect 18748 22596 18889 22624
rect 18748 22584 18754 22596
rect 18877 22593 18889 22596
rect 18923 22624 18935 22627
rect 20898 22624 20904 22636
rect 18923 22596 20904 22624
rect 18923 22593 18935 22596
rect 18877 22587 18935 22593
rect 20898 22584 20904 22596
rect 20956 22584 20962 22636
rect 21082 22584 21088 22636
rect 21140 22584 21146 22636
rect 22094 22584 22100 22636
rect 22152 22584 22158 22636
rect 23934 22584 23940 22636
rect 23992 22584 23998 22636
rect 8389 22559 8447 22565
rect 8389 22525 8401 22559
rect 8435 22556 8447 22559
rect 11146 22556 11152 22568
rect 8435 22528 11152 22556
rect 8435 22525 8447 22528
rect 8389 22519 8447 22525
rect 11146 22516 11152 22528
rect 11204 22516 11210 22568
rect 12621 22559 12679 22565
rect 12621 22525 12633 22559
rect 12667 22556 12679 22559
rect 13354 22556 13360 22568
rect 12667 22528 13360 22556
rect 12667 22525 12679 22528
rect 12621 22519 12679 22525
rect 13354 22516 13360 22528
rect 13412 22516 13418 22568
rect 20162 22516 20168 22568
rect 20220 22556 20226 22568
rect 21269 22559 21327 22565
rect 21269 22556 21281 22559
rect 20220 22528 21281 22556
rect 20220 22516 20226 22528
rect 21269 22525 21281 22528
rect 21315 22525 21327 22559
rect 21269 22519 21327 22525
rect 23290 22516 23296 22568
rect 23348 22516 23354 22568
rect 24762 22516 24768 22568
rect 24820 22516 24826 22568
rect 11790 22488 11796 22500
rect 9876 22460 11796 22488
rect 6914 22380 6920 22432
rect 6972 22420 6978 22432
rect 9876 22429 9904 22460
rect 11790 22448 11796 22460
rect 11848 22448 11854 22500
rect 15194 22448 15200 22500
rect 15252 22488 15258 22500
rect 20349 22491 20407 22497
rect 20349 22488 20361 22491
rect 15252 22460 20361 22488
rect 15252 22448 15258 22460
rect 20349 22457 20361 22460
rect 20395 22488 20407 22491
rect 21082 22488 21088 22500
rect 20395 22460 21088 22488
rect 20395 22457 20407 22460
rect 20349 22451 20407 22457
rect 21082 22448 21088 22460
rect 21140 22448 21146 22500
rect 9861 22423 9919 22429
rect 9861 22420 9873 22423
rect 6972 22392 9873 22420
rect 6972 22380 6978 22392
rect 9861 22389 9873 22392
rect 9907 22389 9919 22423
rect 9861 22383 9919 22389
rect 14090 22380 14096 22432
rect 14148 22380 14154 22432
rect 20714 22380 20720 22432
rect 20772 22380 20778 22432
rect 1104 22330 25852 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 25852 22330
rect 1104 22256 25852 22278
rect 11977 22219 12035 22225
rect 11977 22185 11989 22219
rect 12023 22216 12035 22219
rect 13906 22216 13912 22228
rect 12023 22188 13912 22216
rect 12023 22185 12035 22188
rect 11977 22179 12035 22185
rect 13906 22176 13912 22188
rect 13964 22176 13970 22228
rect 22002 22176 22008 22228
rect 22060 22216 22066 22228
rect 23293 22219 23351 22225
rect 22060 22188 22876 22216
rect 22060 22176 22066 22188
rect 11514 22148 11520 22160
rect 11348 22120 11520 22148
rect 11348 22089 11376 22120
rect 11514 22108 11520 22120
rect 11572 22108 11578 22160
rect 12802 22148 12808 22160
rect 12452 22120 12808 22148
rect 11333 22083 11391 22089
rect 11333 22049 11345 22083
rect 11379 22080 11391 22083
rect 11379 22052 11413 22080
rect 11379 22049 11391 22052
rect 11333 22043 11391 22049
rect 9214 21972 9220 22024
rect 9272 22012 9278 22024
rect 12452 22021 12480 22120
rect 12802 22108 12808 22120
rect 12860 22108 12866 22160
rect 15746 22148 15752 22160
rect 15304 22120 15752 22148
rect 12618 22040 12624 22092
rect 12676 22040 12682 22092
rect 15304 22089 15332 22120
rect 15746 22108 15752 22120
rect 15804 22108 15810 22160
rect 15289 22083 15347 22089
rect 15289 22049 15301 22083
rect 15335 22080 15347 22083
rect 15473 22083 15531 22089
rect 15335 22052 15369 22080
rect 15335 22049 15347 22052
rect 15289 22043 15347 22049
rect 15473 22049 15485 22083
rect 15519 22049 15531 22083
rect 15473 22043 15531 22049
rect 12437 22015 12495 22021
rect 9272 21984 11284 22012
rect 9272 21972 9278 21984
rect 11149 21947 11207 21953
rect 11149 21944 11161 21947
rect 10336 21916 11161 21944
rect 10336 21888 10364 21916
rect 11149 21913 11161 21916
rect 11195 21913 11207 21947
rect 11149 21907 11207 21913
rect 8294 21836 8300 21888
rect 8352 21876 8358 21888
rect 8941 21879 8999 21885
rect 8941 21876 8953 21879
rect 8352 21848 8953 21876
rect 8352 21836 8358 21848
rect 8941 21845 8953 21848
rect 8987 21876 8999 21879
rect 9490 21876 9496 21888
rect 8987 21848 9496 21876
rect 8987 21845 8999 21848
rect 8941 21839 8999 21845
rect 9490 21836 9496 21848
rect 9548 21836 9554 21888
rect 10318 21836 10324 21888
rect 10376 21836 10382 21888
rect 10686 21836 10692 21888
rect 10744 21836 10750 21888
rect 11054 21836 11060 21888
rect 11112 21836 11118 21888
rect 11256 21876 11284 21984
rect 12437 21981 12449 22015
rect 12483 21981 12495 22015
rect 12437 21975 12495 21981
rect 14090 21972 14096 22024
rect 14148 22012 14154 22024
rect 15488 22012 15516 22043
rect 16942 22040 16948 22092
rect 17000 22080 17006 22092
rect 18141 22083 18199 22089
rect 18141 22080 18153 22083
rect 17000 22052 18153 22080
rect 17000 22040 17006 22052
rect 18141 22049 18153 22052
rect 18187 22049 18199 22083
rect 18141 22043 18199 22049
rect 20346 22040 20352 22092
rect 20404 22040 20410 22092
rect 21545 22083 21603 22089
rect 21545 22049 21557 22083
rect 21591 22080 21603 22083
rect 22186 22080 22192 22092
rect 21591 22052 22192 22080
rect 21591 22049 21603 22052
rect 21545 22043 21603 22049
rect 22186 22040 22192 22052
rect 22244 22040 22250 22092
rect 22848 22080 22876 22188
rect 23293 22185 23305 22219
rect 23339 22216 23351 22219
rect 23382 22216 23388 22228
rect 23339 22188 23388 22216
rect 23339 22185 23351 22188
rect 23293 22179 23351 22185
rect 23382 22176 23388 22188
rect 23440 22176 23446 22228
rect 23750 22176 23756 22228
rect 23808 22176 23814 22228
rect 25222 22176 25228 22228
rect 25280 22176 25286 22228
rect 23198 22108 23204 22160
rect 23256 22148 23262 22160
rect 23256 22120 24992 22148
rect 23256 22108 23262 22120
rect 22848 22052 23980 22080
rect 23952 22021 23980 22052
rect 24964 22021 24992 22120
rect 25038 22040 25044 22092
rect 25096 22040 25102 22092
rect 25240 22089 25268 22176
rect 25225 22083 25283 22089
rect 25225 22049 25237 22083
rect 25271 22049 25283 22083
rect 25225 22043 25283 22049
rect 14148 21984 15516 22012
rect 16117 22015 16175 22021
rect 14148 21972 14154 21984
rect 16117 21981 16129 22015
rect 16163 21981 16175 22015
rect 16117 21975 16175 21981
rect 23937 22015 23995 22021
rect 23937 21981 23949 22015
rect 23983 21981 23995 22015
rect 23937 21975 23995 21981
rect 24949 22015 25007 22021
rect 24949 21981 24961 22015
rect 24995 21981 25007 22015
rect 24949 21975 25007 21981
rect 12345 21879 12403 21885
rect 12345 21876 12357 21879
rect 11256 21848 12357 21876
rect 12345 21845 12357 21848
rect 12391 21845 12403 21879
rect 12345 21839 12403 21845
rect 14826 21836 14832 21888
rect 14884 21836 14890 21888
rect 15194 21836 15200 21888
rect 15252 21836 15258 21888
rect 16132 21876 16160 21975
rect 16393 21947 16451 21953
rect 16393 21913 16405 21947
rect 16439 21944 16451 21947
rect 16482 21944 16488 21956
rect 16439 21916 16488 21944
rect 16439 21913 16451 21916
rect 16393 21907 16451 21913
rect 16482 21904 16488 21916
rect 16540 21944 16546 21956
rect 16540 21916 16804 21944
rect 16540 21904 16546 21916
rect 16574 21876 16580 21888
rect 16132 21848 16580 21876
rect 16574 21836 16580 21848
rect 16632 21836 16638 21888
rect 16776 21876 16804 21916
rect 16942 21904 16948 21956
rect 17000 21904 17006 21956
rect 21174 21944 21180 21956
rect 19720 21916 21180 21944
rect 17034 21876 17040 21888
rect 16776 21848 17040 21876
rect 17034 21836 17040 21848
rect 17092 21836 17098 21888
rect 17126 21836 17132 21888
rect 17184 21876 17190 21888
rect 19720 21885 19748 21916
rect 21174 21904 21180 21916
rect 21232 21904 21238 21956
rect 21821 21947 21879 21953
rect 21821 21913 21833 21947
rect 21867 21944 21879 21947
rect 22094 21944 22100 21956
rect 21867 21916 22100 21944
rect 21867 21913 21879 21916
rect 21821 21907 21879 21913
rect 22094 21904 22100 21916
rect 22152 21904 22158 21956
rect 22278 21904 22284 21956
rect 22336 21904 22342 21956
rect 17865 21879 17923 21885
rect 17865 21876 17877 21879
rect 17184 21848 17877 21876
rect 17184 21836 17190 21848
rect 17865 21845 17877 21848
rect 17911 21845 17923 21879
rect 17865 21839 17923 21845
rect 19705 21879 19763 21885
rect 19705 21845 19717 21879
rect 19751 21845 19763 21879
rect 19705 21839 19763 21845
rect 20070 21836 20076 21888
rect 20128 21836 20134 21888
rect 20165 21879 20223 21885
rect 20165 21845 20177 21879
rect 20211 21876 20223 21879
rect 20254 21876 20260 21888
rect 20211 21848 20260 21876
rect 20211 21845 20223 21848
rect 20165 21839 20223 21845
rect 20254 21836 20260 21848
rect 20312 21836 20318 21888
rect 20901 21879 20959 21885
rect 20901 21845 20913 21879
rect 20947 21876 20959 21879
rect 23198 21876 23204 21888
rect 20947 21848 23204 21876
rect 20947 21845 20959 21848
rect 20901 21839 20959 21845
rect 23198 21836 23204 21848
rect 23256 21836 23262 21888
rect 23290 21836 23296 21888
rect 23348 21876 23354 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 23348 21848 24593 21876
rect 23348 21836 23354 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 1104 21786 25852 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 25852 21786
rect 1104 21712 25852 21734
rect 10226 21632 10232 21684
rect 10284 21672 10290 21684
rect 10413 21675 10471 21681
rect 10413 21672 10425 21675
rect 10284 21644 10425 21672
rect 10284 21632 10290 21644
rect 10413 21641 10425 21644
rect 10459 21641 10471 21675
rect 10413 21635 10471 21641
rect 11054 21632 11060 21684
rect 11112 21672 11118 21684
rect 11701 21675 11759 21681
rect 11701 21672 11713 21675
rect 11112 21644 11713 21672
rect 11112 21632 11118 21644
rect 11701 21641 11713 21644
rect 11747 21641 11759 21675
rect 11701 21635 11759 21641
rect 20254 21632 20260 21684
rect 20312 21672 20318 21684
rect 21361 21675 21419 21681
rect 21361 21672 21373 21675
rect 20312 21644 21373 21672
rect 20312 21632 20318 21644
rect 21361 21641 21373 21644
rect 21407 21641 21419 21675
rect 21361 21635 21419 21641
rect 21450 21632 21456 21684
rect 21508 21672 21514 21684
rect 21545 21675 21603 21681
rect 21545 21672 21557 21675
rect 21508 21644 21557 21672
rect 21508 21632 21514 21644
rect 21545 21641 21557 21644
rect 21591 21672 21603 21675
rect 22278 21672 22284 21684
rect 21591 21644 22284 21672
rect 21591 21641 21603 21644
rect 21545 21635 21603 21641
rect 22278 21632 22284 21644
rect 22336 21632 22342 21684
rect 22465 21675 22523 21681
rect 22465 21641 22477 21675
rect 22511 21672 22523 21675
rect 22554 21672 22560 21684
rect 22511 21644 22560 21672
rect 22511 21641 22523 21644
rect 22465 21635 22523 21641
rect 22554 21632 22560 21644
rect 22612 21632 22618 21684
rect 24210 21632 24216 21684
rect 24268 21672 24274 21684
rect 24946 21672 24952 21684
rect 24268 21644 24952 21672
rect 24268 21632 24274 21644
rect 24946 21632 24952 21644
rect 25004 21672 25010 21684
rect 25317 21675 25375 21681
rect 25317 21672 25329 21675
rect 25004 21644 25329 21672
rect 25004 21632 25010 21644
rect 25317 21641 25329 21644
rect 25363 21641 25375 21675
rect 25317 21635 25375 21641
rect 9030 21564 9036 21616
rect 9088 21604 9094 21616
rect 9677 21607 9735 21613
rect 9677 21604 9689 21607
rect 9088 21576 9689 21604
rect 9088 21564 9094 21576
rect 9677 21573 9689 21576
rect 9723 21573 9735 21607
rect 9677 21567 9735 21573
rect 10873 21607 10931 21613
rect 10873 21573 10885 21607
rect 10919 21604 10931 21607
rect 12066 21604 12072 21616
rect 10919 21576 12072 21604
rect 10919 21573 10931 21576
rect 10873 21567 10931 21573
rect 12066 21564 12072 21576
rect 12124 21564 12130 21616
rect 15102 21604 15108 21616
rect 14582 21576 15108 21604
rect 15102 21564 15108 21576
rect 15160 21564 15166 21616
rect 15378 21564 15384 21616
rect 15436 21604 15442 21616
rect 15657 21607 15715 21613
rect 15657 21604 15669 21607
rect 15436 21576 15669 21604
rect 15436 21564 15442 21576
rect 15657 21573 15669 21576
rect 15703 21573 15715 21607
rect 15657 21567 15715 21573
rect 20070 21564 20076 21616
rect 20128 21604 20134 21616
rect 21177 21607 21235 21613
rect 21177 21604 21189 21607
rect 20128 21576 21189 21604
rect 20128 21564 20134 21576
rect 21177 21573 21189 21576
rect 21223 21573 21235 21607
rect 21177 21567 21235 21573
rect 22186 21564 22192 21616
rect 22244 21604 22250 21616
rect 22244 21576 23336 21604
rect 22244 21564 22250 21576
rect 8294 21496 8300 21548
rect 8352 21496 8358 21548
rect 9585 21539 9643 21545
rect 9585 21505 9597 21539
rect 9631 21536 9643 21539
rect 9950 21536 9956 21548
rect 9631 21508 9956 21536
rect 9631 21505 9643 21508
rect 9585 21499 9643 21505
rect 9950 21496 9956 21508
rect 10008 21496 10014 21548
rect 10781 21539 10839 21545
rect 10781 21505 10793 21539
rect 10827 21536 10839 21539
rect 11146 21536 11152 21548
rect 10827 21508 11152 21536
rect 10827 21505 10839 21508
rect 10781 21499 10839 21505
rect 11146 21496 11152 21508
rect 11204 21496 11210 21548
rect 14826 21496 14832 21548
rect 14884 21536 14890 21548
rect 18877 21539 18935 21545
rect 18877 21536 18889 21539
rect 14884 21508 18889 21536
rect 14884 21496 14890 21508
rect 18877 21505 18889 21508
rect 18923 21505 18935 21539
rect 18877 21499 18935 21505
rect 19889 21539 19947 21545
rect 19889 21505 19901 21539
rect 19935 21536 19947 21539
rect 20717 21539 20775 21545
rect 20717 21536 20729 21539
rect 19935 21508 20729 21536
rect 19935 21505 19947 21508
rect 19889 21499 19947 21505
rect 20717 21505 20729 21508
rect 20763 21505 20775 21539
rect 20717 21499 20775 21505
rect 22002 21496 22008 21548
rect 22060 21536 22066 21548
rect 23308 21545 23336 21576
rect 24118 21564 24124 21616
rect 24176 21564 24182 21616
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 22060 21508 22385 21536
rect 22060 21496 22066 21508
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 22373 21499 22431 21505
rect 23293 21539 23351 21545
rect 23293 21505 23305 21539
rect 23339 21505 23351 21539
rect 23293 21499 23351 21505
rect 6917 21471 6975 21477
rect 6917 21437 6929 21471
rect 6963 21437 6975 21471
rect 6917 21431 6975 21437
rect 7193 21471 7251 21477
rect 7193 21437 7205 21471
rect 7239 21468 7251 21471
rect 8478 21468 8484 21480
rect 7239 21440 8484 21468
rect 7239 21437 7251 21440
rect 7193 21431 7251 21437
rect 6932 21332 6960 21431
rect 8478 21428 8484 21440
rect 8536 21428 8542 21480
rect 9306 21428 9312 21480
rect 9364 21468 9370 21480
rect 9769 21471 9827 21477
rect 9769 21468 9781 21471
rect 9364 21440 9781 21468
rect 9364 21428 9370 21440
rect 9769 21437 9781 21440
rect 9815 21437 9827 21471
rect 9769 21431 9827 21437
rect 10962 21428 10968 21480
rect 11020 21428 11026 21480
rect 12434 21428 12440 21480
rect 12492 21468 12498 21480
rect 12710 21468 12716 21480
rect 12492 21440 12716 21468
rect 12492 21428 12498 21440
rect 12710 21428 12716 21440
rect 12768 21468 12774 21480
rect 13081 21471 13139 21477
rect 13081 21468 13093 21471
rect 12768 21440 13093 21468
rect 12768 21428 12774 21440
rect 13081 21437 13093 21440
rect 13127 21437 13139 21471
rect 13081 21431 13139 21437
rect 13357 21471 13415 21477
rect 13357 21437 13369 21471
rect 13403 21468 13415 21471
rect 14090 21468 14096 21480
rect 13403 21440 14096 21468
rect 13403 21437 13415 21440
rect 13357 21431 13415 21437
rect 14090 21428 14096 21440
rect 14148 21428 14154 21480
rect 19058 21428 19064 21480
rect 19116 21468 19122 21480
rect 19981 21471 20039 21477
rect 19981 21468 19993 21471
rect 19116 21440 19993 21468
rect 19116 21428 19122 21440
rect 19981 21437 19993 21440
rect 20027 21437 20039 21471
rect 19981 21431 20039 21437
rect 20162 21428 20168 21480
rect 20220 21428 20226 21480
rect 22649 21471 22707 21477
rect 22649 21437 22661 21471
rect 22695 21437 22707 21471
rect 22649 21431 22707 21437
rect 23569 21471 23627 21477
rect 23569 21437 23581 21471
rect 23615 21468 23627 21471
rect 25314 21468 25320 21480
rect 23615 21440 25320 21468
rect 23615 21437 23627 21440
rect 23569 21431 23627 21437
rect 9217 21403 9275 21409
rect 9217 21369 9229 21403
rect 9263 21400 9275 21403
rect 9263 21372 12434 21400
rect 9263 21369 9275 21372
rect 9217 21363 9275 21369
rect 7742 21332 7748 21344
rect 6932 21304 7748 21332
rect 7742 21292 7748 21304
rect 7800 21292 7806 21344
rect 8294 21292 8300 21344
rect 8352 21332 8358 21344
rect 8662 21332 8668 21344
rect 8352 21304 8668 21332
rect 8352 21292 8358 21304
rect 8662 21292 8668 21304
rect 8720 21292 8726 21344
rect 12406 21332 12434 21372
rect 14550 21360 14556 21412
rect 14608 21400 14614 21412
rect 15841 21403 15899 21409
rect 15841 21400 15853 21403
rect 14608 21372 15853 21400
rect 14608 21360 14614 21372
rect 15841 21369 15853 21372
rect 15887 21369 15899 21403
rect 15841 21363 15899 21369
rect 18693 21403 18751 21409
rect 18693 21369 18705 21403
rect 18739 21400 18751 21403
rect 22462 21400 22468 21412
rect 18739 21372 22468 21400
rect 18739 21369 18751 21372
rect 18693 21363 18751 21369
rect 22462 21360 22468 21372
rect 22520 21360 22526 21412
rect 12526 21332 12532 21344
rect 12406 21304 12532 21332
rect 12526 21292 12532 21304
rect 12584 21292 12590 21344
rect 14366 21292 14372 21344
rect 14424 21332 14430 21344
rect 14829 21335 14887 21341
rect 14829 21332 14841 21335
rect 14424 21304 14841 21332
rect 14424 21292 14430 21304
rect 14829 21301 14841 21304
rect 14875 21332 14887 21335
rect 15010 21332 15016 21344
rect 14875 21304 15016 21332
rect 14875 21301 14887 21304
rect 14829 21295 14887 21301
rect 15010 21292 15016 21304
rect 15068 21292 15074 21344
rect 15102 21292 15108 21344
rect 15160 21292 15166 21344
rect 19058 21292 19064 21344
rect 19116 21332 19122 21344
rect 19153 21335 19211 21341
rect 19153 21332 19165 21335
rect 19116 21304 19165 21332
rect 19116 21292 19122 21304
rect 19153 21301 19165 21304
rect 19199 21301 19211 21335
rect 19153 21295 19211 21301
rect 19518 21292 19524 21344
rect 19576 21292 19582 21344
rect 21726 21292 21732 21344
rect 21784 21332 21790 21344
rect 22005 21335 22063 21341
rect 22005 21332 22017 21335
rect 21784 21304 22017 21332
rect 21784 21292 21790 21304
rect 22005 21301 22017 21304
rect 22051 21301 22063 21335
rect 22664 21332 22692 21431
rect 25314 21428 25320 21440
rect 25372 21428 25378 21480
rect 23566 21332 23572 21344
rect 22664 21304 23572 21332
rect 22005 21295 22063 21301
rect 23566 21292 23572 21304
rect 23624 21292 23630 21344
rect 25038 21292 25044 21344
rect 25096 21292 25102 21344
rect 1104 21242 25852 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 25852 21242
rect 1104 21168 25852 21190
rect 4798 21088 4804 21140
rect 4856 21128 4862 21140
rect 19058 21128 19064 21140
rect 4856 21100 19064 21128
rect 4856 21088 4862 21100
rect 19058 21088 19064 21100
rect 19116 21088 19122 21140
rect 20898 21088 20904 21140
rect 20956 21128 20962 21140
rect 21453 21131 21511 21137
rect 21453 21128 21465 21131
rect 20956 21100 21465 21128
rect 20956 21088 20962 21100
rect 21453 21097 21465 21100
rect 21499 21097 21511 21131
rect 21453 21091 21511 21097
rect 22094 21088 22100 21140
rect 22152 21128 22158 21140
rect 25038 21128 25044 21140
rect 22152 21100 25044 21128
rect 22152 21088 22158 21100
rect 25038 21088 25044 21100
rect 25096 21088 25102 21140
rect 12437 21063 12495 21069
rect 12437 21029 12449 21063
rect 12483 21060 12495 21063
rect 13354 21060 13360 21072
rect 12483 21032 13360 21060
rect 12483 21029 12495 21032
rect 12437 21023 12495 21029
rect 13354 21020 13360 21032
rect 13412 21020 13418 21072
rect 16574 21020 16580 21072
rect 16632 21020 16638 21072
rect 20809 21063 20867 21069
rect 20809 21029 20821 21063
rect 20855 21060 20867 21063
rect 20855 21032 22692 21060
rect 20855 21029 20867 21032
rect 20809 21023 20867 21029
rect 9950 20952 9956 21004
rect 10008 20952 10014 21004
rect 15197 20995 15255 21001
rect 15197 20961 15209 20995
rect 15243 20992 15255 20995
rect 16592 20992 16620 21020
rect 15243 20964 16620 20992
rect 15243 20961 15255 20964
rect 15197 20955 15255 20961
rect 19702 20952 19708 21004
rect 19760 20992 19766 21004
rect 19981 20995 20039 21001
rect 19981 20992 19993 20995
rect 19760 20964 19993 20992
rect 19760 20952 19766 20964
rect 19981 20961 19993 20964
rect 20027 20961 20039 20995
rect 19981 20955 20039 20961
rect 22002 20952 22008 21004
rect 22060 20952 22066 21004
rect 9766 20884 9772 20936
rect 9824 20924 9830 20936
rect 10689 20927 10747 20933
rect 10689 20924 10701 20927
rect 9824 20896 10701 20924
rect 9824 20884 9830 20896
rect 10689 20893 10701 20896
rect 10735 20893 10747 20927
rect 10689 20887 10747 20893
rect 18690 20884 18696 20936
rect 18748 20884 18754 20936
rect 19242 20884 19248 20936
rect 19300 20924 19306 20936
rect 19889 20927 19947 20933
rect 19889 20924 19901 20927
rect 19300 20896 19901 20924
rect 19300 20884 19306 20896
rect 19889 20893 19901 20896
rect 19935 20893 19947 20927
rect 19889 20887 19947 20893
rect 3510 20816 3516 20868
rect 3568 20856 3574 20868
rect 10134 20856 10140 20868
rect 3568 20828 10140 20856
rect 3568 20816 3574 20828
rect 10134 20816 10140 20828
rect 10192 20816 10198 20868
rect 10870 20816 10876 20868
rect 10928 20856 10934 20868
rect 10965 20859 11023 20865
rect 10965 20856 10977 20859
rect 10928 20828 10977 20856
rect 10928 20816 10934 20828
rect 10965 20825 10977 20828
rect 11011 20825 11023 20859
rect 12434 20856 12440 20868
rect 12190 20828 12440 20856
rect 10965 20819 11023 20825
rect 12434 20816 12440 20828
rect 12492 20856 12498 20868
rect 12713 20859 12771 20865
rect 12713 20856 12725 20859
rect 12492 20828 12725 20856
rect 12492 20816 12498 20828
rect 12713 20825 12725 20828
rect 12759 20856 12771 20859
rect 14553 20859 14611 20865
rect 14553 20856 14565 20859
rect 12759 20828 14565 20856
rect 12759 20825 12771 20828
rect 12713 20819 12771 20825
rect 14553 20825 14565 20828
rect 14599 20856 14611 20859
rect 14642 20856 14648 20868
rect 14599 20828 14648 20856
rect 14599 20825 14611 20828
rect 14553 20819 14611 20825
rect 14642 20816 14648 20828
rect 14700 20816 14706 20868
rect 15473 20859 15531 20865
rect 15473 20825 15485 20859
rect 15519 20856 15531 20859
rect 15746 20856 15752 20868
rect 15519 20828 15752 20856
rect 15519 20825 15531 20828
rect 15473 20819 15531 20825
rect 15746 20816 15752 20828
rect 15804 20816 15810 20868
rect 18708 20856 18736 20884
rect 19797 20859 19855 20865
rect 19797 20856 19809 20859
rect 15856 20828 15962 20856
rect 18708 20828 19809 20856
rect 8662 20748 8668 20800
rect 8720 20788 8726 20800
rect 9030 20788 9036 20800
rect 8720 20760 9036 20788
rect 8720 20748 8726 20760
rect 9030 20748 9036 20760
rect 9088 20748 9094 20800
rect 14660 20788 14688 20816
rect 15102 20788 15108 20800
rect 14660 20760 15108 20788
rect 15102 20748 15108 20760
rect 15160 20788 15166 20800
rect 15856 20788 15884 20828
rect 19797 20825 19809 20828
rect 19843 20825 19855 20859
rect 19904 20856 19932 20887
rect 20990 20884 20996 20936
rect 21048 20884 21054 20936
rect 22664 20933 22692 21032
rect 23845 20995 23903 21001
rect 23845 20961 23857 20995
rect 23891 20992 23903 20995
rect 24854 20992 24860 21004
rect 23891 20964 24860 20992
rect 23891 20961 23903 20964
rect 23845 20955 23903 20961
rect 24854 20952 24860 20964
rect 24912 20952 24918 21004
rect 24946 20952 24952 21004
rect 25004 20992 25010 21004
rect 25041 20995 25099 21001
rect 25041 20992 25053 20995
rect 25004 20964 25053 20992
rect 25004 20952 25010 20964
rect 25041 20961 25053 20964
rect 25087 20961 25099 20995
rect 25041 20955 25099 20961
rect 25133 20995 25191 21001
rect 25133 20961 25145 20995
rect 25179 20961 25191 20995
rect 25133 20955 25191 20961
rect 22649 20927 22707 20933
rect 22649 20893 22661 20927
rect 22695 20893 22707 20927
rect 22649 20887 22707 20893
rect 23934 20884 23940 20936
rect 23992 20924 23998 20936
rect 25148 20924 25176 20955
rect 23992 20896 25176 20924
rect 23992 20884 23998 20896
rect 21269 20859 21327 20865
rect 21269 20856 21281 20859
rect 19904 20828 21281 20856
rect 19797 20819 19855 20825
rect 21269 20825 21281 20828
rect 21315 20825 21327 20859
rect 21269 20819 21327 20825
rect 15160 20760 15884 20788
rect 15160 20748 15166 20760
rect 16482 20748 16488 20800
rect 16540 20788 16546 20800
rect 16945 20791 17003 20797
rect 16945 20788 16957 20791
rect 16540 20760 16957 20788
rect 16540 20748 16546 20760
rect 16945 20757 16957 20760
rect 16991 20757 17003 20791
rect 16945 20751 17003 20757
rect 17034 20748 17040 20800
rect 17092 20788 17098 20800
rect 17221 20791 17279 20797
rect 17221 20788 17233 20791
rect 17092 20760 17233 20788
rect 17092 20748 17098 20760
rect 17221 20757 17233 20760
rect 17267 20788 17279 20791
rect 17586 20788 17592 20800
rect 17267 20760 17592 20788
rect 17267 20757 17279 20760
rect 17221 20751 17279 20757
rect 17586 20748 17592 20760
rect 17644 20788 17650 20800
rect 18693 20791 18751 20797
rect 18693 20788 18705 20791
rect 17644 20760 18705 20788
rect 17644 20748 17650 20760
rect 18693 20757 18705 20760
rect 18739 20757 18751 20791
rect 18693 20751 18751 20757
rect 19429 20791 19487 20797
rect 19429 20757 19441 20791
rect 19475 20788 19487 20791
rect 19610 20788 19616 20800
rect 19475 20760 19616 20788
rect 19475 20757 19487 20760
rect 19429 20751 19487 20757
rect 19610 20748 19616 20760
rect 19668 20748 19674 20800
rect 19812 20788 19840 20819
rect 20441 20791 20499 20797
rect 20441 20788 20453 20791
rect 19812 20760 20453 20788
rect 20441 20757 20453 20760
rect 20487 20757 20499 20791
rect 20441 20751 20499 20757
rect 24581 20791 24639 20797
rect 24581 20757 24593 20791
rect 24627 20788 24639 20791
rect 24854 20788 24860 20800
rect 24627 20760 24860 20788
rect 24627 20757 24639 20760
rect 24581 20751 24639 20757
rect 24854 20748 24860 20760
rect 24912 20748 24918 20800
rect 24946 20748 24952 20800
rect 25004 20748 25010 20800
rect 1104 20698 25852 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 25852 20698
rect 1104 20624 25852 20646
rect 10410 20544 10416 20596
rect 10468 20544 10474 20596
rect 10781 20587 10839 20593
rect 10781 20553 10793 20587
rect 10827 20584 10839 20587
rect 12618 20584 12624 20596
rect 10827 20556 12624 20584
rect 10827 20553 10839 20556
rect 10781 20547 10839 20553
rect 12618 20544 12624 20556
rect 12676 20544 12682 20596
rect 13630 20544 13636 20596
rect 13688 20584 13694 20596
rect 15381 20587 15439 20593
rect 15381 20584 15393 20587
rect 13688 20556 15393 20584
rect 13688 20544 13694 20556
rect 15381 20553 15393 20556
rect 15427 20553 15439 20587
rect 15381 20547 15439 20553
rect 15473 20587 15531 20593
rect 15473 20553 15485 20587
rect 15519 20584 15531 20587
rect 15562 20584 15568 20596
rect 15519 20556 15568 20584
rect 15519 20553 15531 20556
rect 15473 20547 15531 20553
rect 15562 20544 15568 20556
rect 15620 20544 15626 20596
rect 19426 20584 19432 20596
rect 16868 20556 19432 20584
rect 8021 20519 8079 20525
rect 8021 20485 8033 20519
rect 8067 20516 8079 20519
rect 8294 20516 8300 20528
rect 8067 20488 8300 20516
rect 8067 20485 8079 20488
rect 8021 20479 8079 20485
rect 8294 20476 8300 20488
rect 8352 20476 8358 20528
rect 9306 20516 9312 20528
rect 9246 20488 9312 20516
rect 9306 20476 9312 20488
rect 9364 20476 9370 20528
rect 14642 20448 14648 20460
rect 14122 20420 14648 20448
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 16868 20457 16896 20556
rect 19426 20544 19432 20556
rect 19484 20544 19490 20596
rect 20806 20544 20812 20596
rect 20864 20544 20870 20596
rect 20898 20544 20904 20596
rect 20956 20544 20962 20596
rect 25314 20544 25320 20596
rect 25372 20544 25378 20596
rect 17126 20476 17132 20528
rect 17184 20476 17190 20528
rect 17586 20476 17592 20528
rect 17644 20476 17650 20528
rect 20824 20516 20852 20544
rect 21453 20519 21511 20525
rect 21453 20516 21465 20519
rect 20824 20488 21465 20516
rect 21453 20485 21465 20488
rect 21499 20485 21511 20519
rect 21453 20479 21511 20485
rect 22738 20476 22744 20528
rect 22796 20516 22802 20528
rect 23382 20516 23388 20528
rect 22796 20488 23388 20516
rect 22796 20476 22802 20488
rect 23382 20476 23388 20488
rect 23440 20476 23446 20528
rect 24118 20476 24124 20528
rect 24176 20516 24182 20528
rect 24176 20488 24334 20516
rect 24176 20476 24182 20488
rect 16853 20451 16911 20457
rect 16853 20417 16865 20451
rect 16899 20417 16911 20451
rect 16853 20411 16911 20417
rect 18414 20408 18420 20460
rect 18472 20448 18478 20460
rect 18690 20448 18696 20460
rect 18472 20420 18696 20448
rect 18472 20408 18478 20420
rect 18690 20408 18696 20420
rect 18748 20408 18754 20460
rect 18782 20408 18788 20460
rect 18840 20448 18846 20460
rect 19150 20448 19156 20460
rect 18840 20420 19156 20448
rect 18840 20408 18846 20420
rect 19150 20408 19156 20420
rect 19208 20408 19214 20460
rect 19245 20451 19303 20457
rect 19245 20417 19257 20451
rect 19291 20448 19303 20451
rect 19794 20448 19800 20460
rect 19291 20420 19800 20448
rect 19291 20417 19303 20420
rect 19245 20411 19303 20417
rect 19794 20408 19800 20420
rect 19852 20408 19858 20460
rect 19889 20451 19947 20457
rect 19889 20417 19901 20451
rect 19935 20448 19947 20451
rect 21818 20448 21824 20460
rect 19935 20420 21824 20448
rect 19935 20417 19947 20420
rect 19889 20411 19947 20417
rect 21818 20408 21824 20420
rect 21876 20408 21882 20460
rect 22186 20408 22192 20460
rect 22244 20408 22250 20460
rect 22462 20408 22468 20460
rect 22520 20448 22526 20460
rect 22925 20451 22983 20457
rect 22925 20448 22937 20451
rect 22520 20420 22937 20448
rect 22520 20408 22526 20420
rect 22925 20417 22937 20420
rect 22971 20417 22983 20451
rect 22925 20411 22983 20417
rect 7742 20340 7748 20392
rect 7800 20340 7806 20392
rect 8478 20340 8484 20392
rect 8536 20380 8542 20392
rect 9490 20380 9496 20392
rect 8536 20352 9496 20380
rect 8536 20340 8542 20352
rect 9490 20340 9496 20352
rect 9548 20380 9554 20392
rect 9769 20383 9827 20389
rect 9548 20352 9720 20380
rect 9548 20340 9554 20352
rect 9692 20312 9720 20352
rect 9769 20349 9781 20383
rect 9815 20380 9827 20383
rect 9950 20380 9956 20392
rect 9815 20352 9956 20380
rect 9815 20349 9827 20352
rect 9769 20343 9827 20349
rect 9950 20340 9956 20352
rect 10008 20340 10014 20392
rect 10226 20340 10232 20392
rect 10284 20380 10290 20392
rect 10873 20383 10931 20389
rect 10873 20380 10885 20383
rect 10284 20352 10885 20380
rect 10284 20340 10290 20352
rect 10873 20349 10885 20352
rect 10919 20349 10931 20383
rect 10873 20343 10931 20349
rect 10965 20383 11023 20389
rect 10965 20349 10977 20383
rect 11011 20349 11023 20383
rect 10965 20343 11023 20349
rect 10980 20312 11008 20343
rect 12710 20340 12716 20392
rect 12768 20340 12774 20392
rect 12989 20383 13047 20389
rect 12989 20349 13001 20383
rect 13035 20380 13047 20383
rect 13446 20380 13452 20392
rect 13035 20352 13452 20380
rect 13035 20349 13047 20352
rect 12989 20343 13047 20349
rect 13446 20340 13452 20352
rect 13504 20380 13510 20392
rect 14366 20380 14372 20392
rect 13504 20352 14372 20380
rect 13504 20340 13510 20352
rect 14366 20340 14372 20352
rect 14424 20340 14430 20392
rect 15565 20383 15623 20389
rect 15565 20380 15577 20383
rect 14476 20352 15577 20380
rect 9692 20284 11008 20312
rect 8478 20204 8484 20256
rect 8536 20244 8542 20256
rect 9306 20244 9312 20256
rect 8536 20216 9312 20244
rect 8536 20204 8542 20216
rect 9306 20204 9312 20216
rect 9364 20244 9370 20256
rect 10137 20247 10195 20253
rect 10137 20244 10149 20247
rect 9364 20216 10149 20244
rect 9364 20204 9370 20216
rect 10137 20213 10149 20216
rect 10183 20244 10195 20247
rect 10410 20244 10416 20256
rect 10183 20216 10416 20244
rect 10183 20213 10195 20216
rect 10137 20207 10195 20213
rect 10410 20204 10416 20216
rect 10468 20204 10474 20256
rect 13538 20204 13544 20256
rect 13596 20244 13602 20256
rect 14476 20253 14504 20352
rect 15565 20349 15577 20352
rect 15611 20349 15623 20383
rect 20990 20380 20996 20392
rect 15565 20343 15623 20349
rect 15672 20352 20996 20380
rect 15102 20272 15108 20324
rect 15160 20312 15166 20324
rect 15672 20312 15700 20352
rect 20990 20340 20996 20352
rect 21048 20340 21054 20392
rect 21085 20383 21143 20389
rect 21085 20349 21097 20383
rect 21131 20380 21143 20383
rect 22278 20380 22284 20392
rect 21131 20352 22284 20380
rect 21131 20349 21143 20352
rect 21085 20343 21143 20349
rect 22278 20340 22284 20352
rect 22336 20340 22342 20392
rect 23566 20340 23572 20392
rect 23624 20340 23630 20392
rect 23845 20383 23903 20389
rect 23845 20349 23857 20383
rect 23891 20380 23903 20383
rect 25130 20380 25136 20392
rect 23891 20352 25136 20380
rect 23891 20349 23903 20352
rect 23845 20343 23903 20349
rect 25130 20340 25136 20352
rect 25188 20340 25194 20392
rect 19150 20312 19156 20324
rect 15160 20284 15700 20312
rect 18524 20284 19156 20312
rect 15160 20272 15166 20284
rect 14461 20247 14519 20253
rect 14461 20244 14473 20247
rect 13596 20216 14473 20244
rect 13596 20204 13602 20216
rect 14461 20213 14473 20216
rect 14507 20213 14519 20247
rect 14461 20207 14519 20213
rect 15013 20247 15071 20253
rect 15013 20213 15025 20247
rect 15059 20244 15071 20247
rect 18524 20244 18552 20284
rect 19150 20272 19156 20284
rect 19208 20272 19214 20324
rect 22005 20315 22063 20321
rect 22005 20281 22017 20315
rect 22051 20312 22063 20315
rect 23474 20312 23480 20324
rect 22051 20284 23480 20312
rect 22051 20281 22063 20284
rect 22005 20275 22063 20281
rect 23474 20272 23480 20284
rect 23532 20272 23538 20324
rect 15059 20216 18552 20244
rect 18601 20247 18659 20253
rect 15059 20213 15071 20216
rect 15013 20207 15071 20213
rect 18601 20213 18613 20247
rect 18647 20244 18659 20247
rect 18690 20244 18696 20256
rect 18647 20216 18696 20244
rect 18647 20213 18659 20216
rect 18601 20207 18659 20213
rect 18690 20204 18696 20216
rect 18748 20204 18754 20256
rect 19058 20204 19064 20256
rect 19116 20204 19122 20256
rect 19705 20247 19763 20253
rect 19705 20213 19717 20247
rect 19751 20244 19763 20247
rect 19794 20244 19800 20256
rect 19751 20216 19800 20244
rect 19751 20213 19763 20216
rect 19705 20207 19763 20213
rect 19794 20204 19800 20216
rect 19852 20204 19858 20256
rect 20441 20247 20499 20253
rect 20441 20213 20453 20247
rect 20487 20244 20499 20247
rect 20530 20244 20536 20256
rect 20487 20216 20536 20244
rect 20487 20213 20499 20216
rect 20441 20207 20499 20213
rect 20530 20204 20536 20216
rect 20588 20204 20594 20256
rect 22738 20204 22744 20256
rect 22796 20204 22802 20256
rect 1104 20154 25852 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 25852 20154
rect 1104 20080 25852 20102
rect 8478 20000 8484 20052
rect 8536 20000 8542 20052
rect 11333 20043 11391 20049
rect 11333 20009 11345 20043
rect 11379 20040 11391 20043
rect 13998 20040 14004 20052
rect 11379 20012 14004 20040
rect 11379 20009 11391 20012
rect 11333 20003 11391 20009
rect 13998 20000 14004 20012
rect 14056 20000 14062 20052
rect 15746 20000 15752 20052
rect 15804 20040 15810 20052
rect 16025 20043 16083 20049
rect 16025 20040 16037 20043
rect 15804 20012 16037 20040
rect 15804 20000 15810 20012
rect 16025 20009 16037 20012
rect 16071 20009 16083 20043
rect 16025 20003 16083 20009
rect 16485 20043 16543 20049
rect 16485 20009 16497 20043
rect 16531 20040 16543 20043
rect 22186 20040 22192 20052
rect 16531 20012 22192 20040
rect 16531 20009 16543 20012
rect 16485 20003 16543 20009
rect 22186 20000 22192 20012
rect 22244 20000 22250 20052
rect 23845 20043 23903 20049
rect 23845 20009 23857 20043
rect 23891 20040 23903 20043
rect 23934 20040 23940 20052
rect 23891 20012 23940 20040
rect 23891 20009 23903 20012
rect 23845 20003 23903 20009
rect 23934 20000 23940 20012
rect 23992 20000 23998 20052
rect 17126 19932 17132 19984
rect 17184 19972 17190 19984
rect 17184 19944 18092 19972
rect 17184 19932 17190 19944
rect 7742 19864 7748 19916
rect 7800 19904 7806 19916
rect 9125 19907 9183 19913
rect 9125 19904 9137 19907
rect 7800 19876 9137 19904
rect 7800 19864 7806 19876
rect 9125 19873 9137 19876
rect 9171 19904 9183 19907
rect 9766 19904 9772 19916
rect 9171 19876 9772 19904
rect 9171 19873 9183 19876
rect 9125 19867 9183 19873
rect 9766 19864 9772 19876
rect 9824 19864 9830 19916
rect 11974 19864 11980 19916
rect 12032 19864 12038 19916
rect 14553 19907 14611 19913
rect 14553 19873 14565 19907
rect 14599 19904 14611 19907
rect 15838 19904 15844 19916
rect 14599 19876 15844 19904
rect 14599 19873 14611 19876
rect 14553 19867 14611 19873
rect 15838 19864 15844 19876
rect 15896 19864 15902 19916
rect 17862 19864 17868 19916
rect 17920 19904 17926 19916
rect 18064 19913 18092 19944
rect 17957 19907 18015 19913
rect 17957 19904 17969 19907
rect 17920 19876 17969 19904
rect 17920 19864 17926 19876
rect 17957 19873 17969 19876
rect 18003 19873 18015 19907
rect 17957 19867 18015 19873
rect 18049 19907 18107 19913
rect 18049 19873 18061 19907
rect 18095 19873 18107 19907
rect 18049 19867 18107 19873
rect 19889 19907 19947 19913
rect 19889 19873 19901 19907
rect 19935 19904 19947 19907
rect 20254 19904 20260 19916
rect 19935 19876 20260 19904
rect 19935 19873 19947 19876
rect 19889 19867 19947 19873
rect 20254 19864 20260 19876
rect 20312 19904 20318 19916
rect 22097 19907 22155 19913
rect 22097 19904 22109 19907
rect 20312 19876 22109 19904
rect 20312 19864 20318 19876
rect 22097 19873 22109 19876
rect 22143 19873 22155 19907
rect 22097 19867 22155 19873
rect 12710 19796 12716 19848
rect 12768 19836 12774 19848
rect 14277 19839 14335 19845
rect 14277 19836 14289 19839
rect 12768 19808 14289 19836
rect 12768 19796 12774 19808
rect 14277 19805 14289 19808
rect 14323 19805 14335 19839
rect 14277 19799 14335 19805
rect 16666 19796 16672 19848
rect 16724 19796 16730 19848
rect 18598 19796 18604 19848
rect 18656 19836 18662 19848
rect 18877 19839 18935 19845
rect 18877 19836 18889 19839
rect 18656 19808 18889 19836
rect 18656 19796 18662 19808
rect 18877 19805 18889 19808
rect 18923 19805 18935 19839
rect 21450 19836 21456 19848
rect 21298 19808 21456 19836
rect 18877 19799 18935 19805
rect 21450 19796 21456 19808
rect 21508 19796 21514 19848
rect 8478 19728 8484 19780
rect 8536 19768 8542 19780
rect 9398 19768 9404 19780
rect 8536 19740 9404 19768
rect 8536 19728 8542 19740
rect 9398 19728 9404 19740
rect 9456 19728 9462 19780
rect 10410 19728 10416 19780
rect 10468 19728 10474 19780
rect 11054 19728 11060 19780
rect 11112 19768 11118 19780
rect 11793 19771 11851 19777
rect 11793 19768 11805 19771
rect 11112 19740 11805 19768
rect 11112 19728 11118 19740
rect 11793 19737 11805 19740
rect 11839 19737 11851 19771
rect 11793 19731 11851 19737
rect 14642 19728 14648 19780
rect 14700 19768 14706 19780
rect 14700 19740 15042 19768
rect 14700 19728 14706 19740
rect 10870 19660 10876 19712
rect 10928 19660 10934 19712
rect 11698 19660 11704 19712
rect 11756 19660 11762 19712
rect 14936 19700 14964 19740
rect 15838 19728 15844 19780
rect 15896 19768 15902 19780
rect 17865 19771 17923 19777
rect 17865 19768 17877 19771
rect 15896 19740 17877 19768
rect 15896 19728 15902 19740
rect 17865 19737 17877 19740
rect 17911 19737 17923 19771
rect 17865 19731 17923 19737
rect 18340 19740 20116 19768
rect 16945 19703 17003 19709
rect 16945 19700 16957 19703
rect 14936 19672 16957 19700
rect 16945 19669 16957 19672
rect 16991 19700 17003 19703
rect 17034 19700 17040 19712
rect 16991 19672 17040 19700
rect 16991 19669 17003 19672
rect 16945 19663 17003 19669
rect 17034 19660 17040 19672
rect 17092 19660 17098 19712
rect 17497 19703 17555 19709
rect 17497 19669 17509 19703
rect 17543 19700 17555 19703
rect 18340 19700 18368 19740
rect 17543 19672 18368 19700
rect 17543 19669 17555 19672
rect 17497 19663 17555 19669
rect 18414 19660 18420 19712
rect 18472 19700 18478 19712
rect 18693 19703 18751 19709
rect 18693 19700 18705 19703
rect 18472 19672 18705 19700
rect 18472 19660 18478 19672
rect 18693 19669 18705 19672
rect 18739 19669 18751 19703
rect 20088 19700 20116 19740
rect 20162 19728 20168 19780
rect 20220 19728 20226 19780
rect 22373 19771 22431 19777
rect 22373 19768 22385 19771
rect 22066 19740 22385 19768
rect 21450 19700 21456 19712
rect 20088 19672 21456 19700
rect 18693 19663 18751 19669
rect 21450 19660 21456 19672
rect 21508 19660 21514 19712
rect 21634 19660 21640 19712
rect 21692 19700 21698 19712
rect 22066 19700 22094 19740
rect 22373 19737 22385 19740
rect 22419 19737 22431 19771
rect 24118 19768 24124 19780
rect 23598 19740 24124 19768
rect 22373 19731 22431 19737
rect 24118 19728 24124 19740
rect 24176 19768 24182 19780
rect 25406 19768 25412 19780
rect 24176 19740 25412 19768
rect 24176 19728 24182 19740
rect 25406 19728 25412 19740
rect 25464 19728 25470 19780
rect 21692 19672 22094 19700
rect 21692 19660 21698 19672
rect 23382 19660 23388 19712
rect 23440 19700 23446 19712
rect 24397 19703 24455 19709
rect 24397 19700 24409 19703
rect 23440 19672 24409 19700
rect 23440 19660 23446 19672
rect 24397 19669 24409 19672
rect 24443 19700 24455 19703
rect 24946 19700 24952 19712
rect 24443 19672 24952 19700
rect 24443 19669 24455 19672
rect 24397 19663 24455 19669
rect 24946 19660 24952 19672
rect 25004 19660 25010 19712
rect 1104 19610 25852 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 25852 19610
rect 1104 19536 25852 19558
rect 8754 19456 8760 19508
rect 8812 19456 8818 19508
rect 11698 19456 11704 19508
rect 11756 19456 11762 19508
rect 11790 19456 11796 19508
rect 11848 19496 11854 19508
rect 16853 19499 16911 19505
rect 11848 19468 15240 19496
rect 11848 19456 11854 19468
rect 8386 19428 8392 19440
rect 8050 19400 8392 19428
rect 8386 19388 8392 19400
rect 8444 19388 8450 19440
rect 9030 19320 9036 19372
rect 9088 19360 9094 19372
rect 9125 19363 9183 19369
rect 9125 19360 9137 19363
rect 9088 19332 9137 19360
rect 9088 19320 9094 19332
rect 9125 19329 9137 19332
rect 9171 19329 9183 19363
rect 9125 19323 9183 19329
rect 9217 19363 9275 19369
rect 9217 19329 9229 19363
rect 9263 19360 9275 19363
rect 10134 19360 10140 19372
rect 9263 19332 10140 19360
rect 9263 19329 9275 19332
rect 9217 19323 9275 19329
rect 10134 19320 10140 19332
rect 10192 19320 10198 19372
rect 10410 19320 10416 19372
rect 10468 19360 10474 19372
rect 15212 19369 15240 19468
rect 16853 19465 16865 19499
rect 16899 19465 16911 19499
rect 16853 19459 16911 19465
rect 16868 19428 16896 19459
rect 17310 19456 17316 19508
rect 17368 19456 17374 19508
rect 18969 19499 19027 19505
rect 18969 19465 18981 19499
rect 19015 19465 19027 19499
rect 18969 19459 19027 19465
rect 18984 19428 19012 19459
rect 19518 19456 19524 19508
rect 19576 19496 19582 19508
rect 20441 19499 20499 19505
rect 20441 19496 20453 19499
rect 19576 19468 20453 19496
rect 19576 19456 19582 19468
rect 20441 19465 20453 19468
rect 20487 19465 20499 19499
rect 20441 19459 20499 19465
rect 20533 19499 20591 19505
rect 20533 19465 20545 19499
rect 20579 19496 20591 19499
rect 20714 19496 20720 19508
rect 20579 19468 20720 19496
rect 20579 19465 20591 19468
rect 20533 19459 20591 19465
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 22649 19499 22707 19505
rect 22649 19465 22661 19499
rect 22695 19496 22707 19499
rect 24578 19496 24584 19508
rect 22695 19468 24584 19496
rect 22695 19465 22707 19468
rect 22649 19459 22707 19465
rect 24578 19456 24584 19468
rect 24636 19456 24642 19508
rect 25130 19456 25136 19508
rect 25188 19456 25194 19508
rect 25406 19456 25412 19508
rect 25464 19456 25470 19508
rect 22186 19428 22192 19440
rect 16868 19400 18920 19428
rect 18984 19400 22192 19428
rect 15197 19363 15255 19369
rect 10468 19332 10916 19360
rect 13938 19332 14688 19360
rect 10468 19320 10474 19332
rect 6546 19252 6552 19304
rect 6604 19252 6610 19304
rect 6825 19295 6883 19301
rect 6825 19261 6837 19295
rect 6871 19292 6883 19295
rect 6914 19292 6920 19304
rect 6871 19264 6920 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 6914 19252 6920 19264
rect 6972 19252 6978 19304
rect 9306 19252 9312 19304
rect 9364 19252 9370 19304
rect 10888 19224 10916 19332
rect 10962 19252 10968 19304
rect 11020 19292 11026 19304
rect 11149 19295 11207 19301
rect 11149 19292 11161 19295
rect 11020 19264 11161 19292
rect 11020 19252 11026 19264
rect 11149 19261 11161 19264
rect 11195 19261 11207 19295
rect 12434 19292 12440 19304
rect 11149 19255 11207 19261
rect 11256 19264 12440 19292
rect 11057 19227 11115 19233
rect 11057 19224 11069 19227
rect 10888 19196 11069 19224
rect 11057 19193 11069 19196
rect 11103 19224 11115 19227
rect 11256 19224 11284 19264
rect 12434 19252 12440 19264
rect 12492 19252 12498 19304
rect 12529 19295 12587 19301
rect 12529 19261 12541 19295
rect 12575 19261 12587 19295
rect 12529 19255 12587 19261
rect 12805 19295 12863 19301
rect 12805 19261 12817 19295
rect 12851 19292 12863 19295
rect 13538 19292 13544 19304
rect 12851 19264 13544 19292
rect 12851 19261 12863 19264
rect 12805 19255 12863 19261
rect 11103 19196 11284 19224
rect 11103 19193 11115 19196
rect 11057 19187 11115 19193
rect 8294 19116 8300 19168
rect 8352 19156 8358 19168
rect 9122 19156 9128 19168
rect 8352 19128 9128 19156
rect 8352 19116 8358 19128
rect 9122 19116 9128 19128
rect 9180 19116 9186 19168
rect 12544 19156 12572 19255
rect 13538 19252 13544 19264
rect 13596 19252 13602 19304
rect 14660 19168 14688 19332
rect 15197 19329 15209 19363
rect 15243 19329 15255 19363
rect 15197 19323 15255 19329
rect 16114 19320 16120 19372
rect 16172 19320 16178 19372
rect 16206 19320 16212 19372
rect 16264 19360 16270 19372
rect 17221 19363 17279 19369
rect 17221 19360 17233 19363
rect 16264 19332 17233 19360
rect 16264 19320 16270 19332
rect 17221 19329 17233 19332
rect 17267 19329 17279 19363
rect 18892 19360 18920 19400
rect 22186 19388 22192 19400
rect 22244 19388 22250 19440
rect 23566 19428 23572 19440
rect 23400 19400 23572 19428
rect 18892 19332 19104 19360
rect 17221 19323 17279 19329
rect 15746 19252 15752 19304
rect 15804 19292 15810 19304
rect 17405 19295 17463 19301
rect 17405 19292 17417 19295
rect 15804 19264 17417 19292
rect 15804 19252 15810 19264
rect 17405 19261 17417 19264
rect 17451 19261 17463 19295
rect 19076 19292 19104 19332
rect 19150 19320 19156 19372
rect 19208 19320 19214 19372
rect 19242 19320 19248 19372
rect 19300 19360 19306 19372
rect 23400 19369 23428 19400
rect 23566 19388 23572 19400
rect 23624 19388 23630 19440
rect 23661 19431 23719 19437
rect 23661 19397 23673 19431
rect 23707 19428 23719 19431
rect 23934 19428 23940 19440
rect 23707 19400 23940 19428
rect 23707 19397 23719 19400
rect 23661 19391 23719 19397
rect 23934 19388 23940 19400
rect 23992 19388 23998 19440
rect 24118 19388 24124 19440
rect 24176 19388 24182 19440
rect 21269 19363 21327 19369
rect 19300 19332 20116 19360
rect 19300 19320 19306 19332
rect 19334 19292 19340 19304
rect 19076 19264 19340 19292
rect 17405 19255 17463 19261
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 14826 19184 14832 19236
rect 14884 19224 14890 19236
rect 20088 19233 20116 19332
rect 21269 19329 21281 19363
rect 21315 19360 21327 19363
rect 22557 19363 22615 19369
rect 22557 19360 22569 19363
rect 21315 19332 22569 19360
rect 21315 19329 21327 19332
rect 21269 19323 21327 19329
rect 22557 19329 22569 19332
rect 22603 19329 22615 19363
rect 22557 19323 22615 19329
rect 23385 19363 23443 19369
rect 23385 19329 23397 19363
rect 23431 19329 23443 19363
rect 23385 19323 23443 19329
rect 20717 19295 20775 19301
rect 20717 19261 20729 19295
rect 20763 19292 20775 19295
rect 21634 19292 21640 19304
rect 20763 19264 21640 19292
rect 20763 19261 20775 19264
rect 20717 19255 20775 19261
rect 21634 19252 21640 19264
rect 21692 19252 21698 19304
rect 22094 19252 22100 19304
rect 22152 19292 22158 19304
rect 22741 19295 22799 19301
rect 22741 19292 22753 19295
rect 22152 19264 22753 19292
rect 22152 19252 22158 19264
rect 22741 19261 22753 19264
rect 22787 19261 22799 19295
rect 22741 19255 22799 19261
rect 15933 19227 15991 19233
rect 15933 19224 15945 19227
rect 14884 19196 15945 19224
rect 14884 19184 14890 19196
rect 15933 19193 15945 19196
rect 15979 19193 15991 19227
rect 15933 19187 15991 19193
rect 20073 19227 20131 19233
rect 20073 19193 20085 19227
rect 20119 19193 20131 19227
rect 20073 19187 20131 19193
rect 21542 19184 21548 19236
rect 21600 19224 21606 19236
rect 21818 19224 21824 19236
rect 21600 19196 21824 19224
rect 21600 19184 21606 19196
rect 21818 19184 21824 19196
rect 21876 19184 21882 19236
rect 21910 19184 21916 19236
rect 21968 19224 21974 19236
rect 22189 19227 22247 19233
rect 22189 19224 22201 19227
rect 21968 19196 22201 19224
rect 21968 19184 21974 19196
rect 22189 19193 22201 19196
rect 22235 19193 22247 19227
rect 22189 19187 22247 19193
rect 12802 19156 12808 19168
rect 12544 19128 12808 19156
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 14277 19159 14335 19165
rect 14277 19125 14289 19159
rect 14323 19156 14335 19159
rect 14366 19156 14372 19168
rect 14323 19128 14372 19156
rect 14323 19125 14335 19128
rect 14277 19119 14335 19125
rect 14366 19116 14372 19128
rect 14424 19116 14430 19168
rect 14642 19116 14648 19168
rect 14700 19116 14706 19168
rect 15013 19159 15071 19165
rect 15013 19125 15025 19159
rect 15059 19156 15071 19159
rect 15102 19156 15108 19168
rect 15059 19128 15108 19156
rect 15059 19125 15071 19128
rect 15013 19119 15071 19125
rect 15102 19116 15108 19128
rect 15160 19116 15166 19168
rect 1104 19066 25852 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 25852 19066
rect 1104 18992 25852 19014
rect 10042 18912 10048 18964
rect 10100 18912 10106 18964
rect 10778 18912 10784 18964
rect 10836 18952 10842 18964
rect 12713 18955 12771 18961
rect 12713 18952 12725 18955
rect 10836 18924 12725 18952
rect 10836 18912 10842 18924
rect 12713 18921 12725 18924
rect 12759 18921 12771 18955
rect 12713 18915 12771 18921
rect 25225 18955 25283 18961
rect 25225 18921 25237 18955
rect 25271 18952 25283 18955
rect 25590 18952 25596 18964
rect 25271 18924 25596 18952
rect 25271 18921 25283 18924
rect 25225 18915 25283 18921
rect 7926 18844 7932 18896
rect 7984 18884 7990 18896
rect 11054 18884 11060 18896
rect 7984 18856 11060 18884
rect 7984 18844 7990 18856
rect 11054 18844 11060 18856
rect 11112 18844 11118 18896
rect 11517 18887 11575 18893
rect 11517 18853 11529 18887
rect 11563 18884 11575 18887
rect 16666 18884 16672 18896
rect 11563 18856 16672 18884
rect 11563 18853 11575 18856
rect 11517 18847 11575 18853
rect 16666 18844 16672 18856
rect 16724 18844 16730 18896
rect 24394 18884 24400 18896
rect 22066 18856 24400 18884
rect 6917 18819 6975 18825
rect 6917 18785 6929 18819
rect 6963 18816 6975 18819
rect 8294 18816 8300 18828
rect 6963 18788 8300 18816
rect 6963 18785 6975 18788
rect 6917 18779 6975 18785
rect 8294 18776 8300 18788
rect 8352 18776 8358 18828
rect 10594 18776 10600 18828
rect 10652 18776 10658 18828
rect 10870 18776 10876 18828
rect 10928 18816 10934 18828
rect 12069 18819 12127 18825
rect 12069 18816 12081 18819
rect 10928 18788 12081 18816
rect 10928 18776 10934 18788
rect 12069 18785 12081 18788
rect 12115 18785 12127 18819
rect 13265 18819 13323 18825
rect 13265 18816 13277 18819
rect 12069 18779 12127 18785
rect 12268 18788 13277 18816
rect 6638 18708 6644 18760
rect 6696 18708 6702 18760
rect 8662 18708 8668 18760
rect 8720 18748 8726 18760
rect 9677 18751 9735 18757
rect 9677 18748 9689 18751
rect 8720 18720 9689 18748
rect 8720 18708 8726 18720
rect 9677 18717 9689 18720
rect 9723 18748 9735 18751
rect 10413 18751 10471 18757
rect 10413 18748 10425 18751
rect 9723 18720 10425 18748
rect 9723 18717 9735 18720
rect 9677 18711 9735 18717
rect 10413 18717 10425 18720
rect 10459 18717 10471 18751
rect 10612 18748 10640 18776
rect 11057 18751 11115 18757
rect 11057 18748 11069 18751
rect 10612 18720 11069 18748
rect 10413 18711 10471 18717
rect 11057 18717 11069 18720
rect 11103 18748 11115 18751
rect 11698 18748 11704 18760
rect 11103 18720 11704 18748
rect 11103 18717 11115 18720
rect 11057 18711 11115 18717
rect 11698 18708 11704 18720
rect 11756 18708 11762 18760
rect 11977 18751 12035 18757
rect 11977 18717 11989 18751
rect 12023 18748 12035 18751
rect 12158 18748 12164 18760
rect 12023 18720 12164 18748
rect 12023 18717 12035 18720
rect 11977 18711 12035 18717
rect 12158 18708 12164 18720
rect 12216 18708 12222 18760
rect 8294 18680 8300 18692
rect 8142 18652 8300 18680
rect 8294 18640 8300 18652
rect 8352 18680 8358 18692
rect 8757 18683 8815 18689
rect 8757 18680 8769 18683
rect 8352 18652 8769 18680
rect 8352 18640 8358 18652
rect 8757 18649 8769 18652
rect 8803 18649 8815 18683
rect 8757 18643 8815 18649
rect 9490 18640 9496 18692
rect 9548 18680 9554 18692
rect 12268 18680 12296 18788
rect 13265 18785 13277 18788
rect 13311 18785 13323 18819
rect 13265 18779 13323 18785
rect 17494 18776 17500 18828
rect 17552 18776 17558 18828
rect 17221 18751 17279 18757
rect 17221 18717 17233 18751
rect 17267 18748 17279 18751
rect 17310 18748 17316 18760
rect 17267 18720 17316 18748
rect 17267 18717 17279 18720
rect 17221 18711 17279 18717
rect 17310 18708 17316 18720
rect 17368 18748 17374 18760
rect 17770 18748 17776 18760
rect 17368 18720 17776 18748
rect 17368 18708 17374 18720
rect 17770 18708 17776 18720
rect 17828 18748 17834 18760
rect 17865 18751 17923 18757
rect 17865 18748 17877 18751
rect 17828 18720 17877 18748
rect 17828 18708 17834 18720
rect 17865 18717 17877 18720
rect 17911 18717 17923 18751
rect 17865 18711 17923 18717
rect 21453 18751 21511 18757
rect 21453 18717 21465 18751
rect 21499 18748 21511 18751
rect 22066 18748 22094 18856
rect 24394 18844 24400 18856
rect 24452 18844 24458 18896
rect 23842 18776 23848 18828
rect 23900 18776 23906 18828
rect 21499 18720 22094 18748
rect 21499 18717 21511 18720
rect 21453 18711 21511 18717
rect 22186 18708 22192 18760
rect 22244 18708 22250 18760
rect 22738 18708 22744 18760
rect 22796 18708 22802 18760
rect 24673 18751 24731 18757
rect 24673 18717 24685 18751
rect 24719 18748 24731 18751
rect 25240 18748 25268 18915
rect 25590 18912 25596 18924
rect 25648 18912 25654 18964
rect 24719 18720 25268 18748
rect 24719 18717 24731 18720
rect 24673 18711 24731 18717
rect 9548 18652 12296 18680
rect 9548 18640 9554 18652
rect 12342 18640 12348 18692
rect 12400 18680 12406 18692
rect 23382 18680 23388 18692
rect 12400 18652 23388 18680
rect 12400 18640 12406 18652
rect 23382 18640 23388 18652
rect 23440 18640 23446 18692
rect 24857 18683 24915 18689
rect 24857 18649 24869 18683
rect 24903 18680 24915 18683
rect 25222 18680 25228 18692
rect 24903 18652 25228 18680
rect 24903 18649 24915 18652
rect 24857 18643 24915 18649
rect 25222 18640 25228 18652
rect 25280 18640 25286 18692
rect 8389 18615 8447 18621
rect 8389 18581 8401 18615
rect 8435 18612 8447 18615
rect 8478 18612 8484 18624
rect 8435 18584 8484 18612
rect 8435 18581 8447 18584
rect 8389 18575 8447 18581
rect 8478 18572 8484 18584
rect 8536 18572 8542 18624
rect 10505 18615 10563 18621
rect 10505 18581 10517 18615
rect 10551 18612 10563 18615
rect 10870 18612 10876 18624
rect 10551 18584 10876 18612
rect 10551 18581 10563 18584
rect 10505 18575 10563 18581
rect 10870 18572 10876 18584
rect 10928 18572 10934 18624
rect 11054 18572 11060 18624
rect 11112 18612 11118 18624
rect 11885 18615 11943 18621
rect 11885 18612 11897 18615
rect 11112 18584 11897 18612
rect 11112 18572 11118 18584
rect 11885 18581 11897 18584
rect 11931 18581 11943 18615
rect 11885 18575 11943 18581
rect 12618 18572 12624 18624
rect 12676 18612 12682 18624
rect 13081 18615 13139 18621
rect 13081 18612 13093 18615
rect 12676 18584 13093 18612
rect 12676 18572 12682 18584
rect 13081 18581 13093 18584
rect 13127 18581 13139 18615
rect 13081 18575 13139 18581
rect 13173 18615 13231 18621
rect 13173 18581 13185 18615
rect 13219 18612 13231 18615
rect 13446 18612 13452 18624
rect 13219 18584 13452 18612
rect 13219 18581 13231 18584
rect 13173 18575 13231 18581
rect 13446 18572 13452 18584
rect 13504 18572 13510 18624
rect 13814 18572 13820 18624
rect 13872 18572 13878 18624
rect 14274 18572 14280 18624
rect 14332 18572 14338 18624
rect 16853 18615 16911 18621
rect 16853 18581 16865 18615
rect 16899 18612 16911 18615
rect 17034 18612 17040 18624
rect 16899 18584 17040 18612
rect 16899 18581 16911 18584
rect 16853 18575 16911 18581
rect 17034 18572 17040 18584
rect 17092 18572 17098 18624
rect 17126 18572 17132 18624
rect 17184 18612 17190 18624
rect 17313 18615 17371 18621
rect 17313 18612 17325 18615
rect 17184 18584 17325 18612
rect 17184 18572 17190 18584
rect 17313 18581 17325 18584
rect 17359 18612 17371 18615
rect 17586 18612 17592 18624
rect 17359 18584 17592 18612
rect 17359 18581 17371 18584
rect 17313 18575 17371 18581
rect 17586 18572 17592 18584
rect 17644 18612 17650 18624
rect 18049 18615 18107 18621
rect 18049 18612 18061 18615
rect 17644 18584 18061 18612
rect 17644 18572 17650 18584
rect 18049 18581 18061 18584
rect 18095 18581 18107 18615
rect 18049 18575 18107 18581
rect 20530 18572 20536 18624
rect 20588 18612 20594 18624
rect 21269 18615 21327 18621
rect 21269 18612 21281 18615
rect 20588 18584 21281 18612
rect 20588 18572 20594 18584
rect 21269 18581 21281 18584
rect 21315 18581 21327 18615
rect 21269 18575 21327 18581
rect 22005 18615 22063 18621
rect 22005 18581 22017 18615
rect 22051 18612 22063 18615
rect 22094 18612 22100 18624
rect 22051 18584 22100 18612
rect 22051 18581 22063 18584
rect 22005 18575 22063 18581
rect 22094 18572 22100 18584
rect 22152 18572 22158 18624
rect 1104 18522 25852 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 25852 18522
rect 1104 18448 25852 18470
rect 9490 18368 9496 18420
rect 9548 18368 9554 18420
rect 9953 18411 10011 18417
rect 9953 18377 9965 18411
rect 9999 18377 10011 18411
rect 9953 18371 10011 18377
rect 10413 18411 10471 18417
rect 10413 18377 10425 18411
rect 10459 18408 10471 18411
rect 10502 18408 10508 18420
rect 10459 18380 10508 18408
rect 10459 18377 10471 18380
rect 10413 18371 10471 18377
rect 8294 18300 8300 18352
rect 8352 18340 8358 18352
rect 9968 18340 9996 18371
rect 10502 18368 10508 18380
rect 10560 18368 10566 18420
rect 10778 18368 10784 18420
rect 10836 18408 10842 18420
rect 12342 18408 12348 18420
rect 10836 18380 12348 18408
rect 10836 18368 10842 18380
rect 12342 18368 12348 18380
rect 12400 18368 12406 18420
rect 13814 18368 13820 18420
rect 13872 18408 13878 18420
rect 14277 18411 14335 18417
rect 14277 18408 14289 18411
rect 13872 18380 14289 18408
rect 13872 18368 13878 18380
rect 14277 18377 14289 18380
rect 14323 18377 14335 18411
rect 14277 18371 14335 18377
rect 14921 18411 14979 18417
rect 14921 18377 14933 18411
rect 14967 18408 14979 18411
rect 16666 18408 16672 18420
rect 14967 18380 16672 18408
rect 14967 18377 14979 18380
rect 14921 18371 14979 18377
rect 11790 18340 11796 18352
rect 8352 18312 8510 18340
rect 9968 18312 11796 18340
rect 8352 18300 8358 18312
rect 11790 18300 11796 18312
rect 11848 18300 11854 18352
rect 14185 18343 14243 18349
rect 14185 18309 14197 18343
rect 14231 18340 14243 18343
rect 14936 18340 14964 18371
rect 16666 18368 16672 18380
rect 16724 18368 16730 18420
rect 22646 18340 22652 18352
rect 14231 18312 14964 18340
rect 21284 18312 22652 18340
rect 14231 18309 14243 18312
rect 14185 18303 14243 18309
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18272 10379 18275
rect 10410 18272 10416 18284
rect 10367 18244 10416 18272
rect 10367 18241 10379 18244
rect 10321 18235 10379 18241
rect 10410 18232 10416 18244
rect 10468 18232 10474 18284
rect 11241 18275 11299 18281
rect 11241 18272 11253 18275
rect 10520 18244 11253 18272
rect 6638 18164 6644 18216
rect 6696 18204 6702 18216
rect 7745 18207 7803 18213
rect 7745 18204 7757 18207
rect 6696 18176 7757 18204
rect 6696 18164 6702 18176
rect 7745 18173 7757 18176
rect 7791 18173 7803 18207
rect 7745 18167 7803 18173
rect 8021 18207 8079 18213
rect 8021 18173 8033 18207
rect 8067 18204 8079 18207
rect 10520 18204 10548 18244
rect 11241 18241 11253 18244
rect 11287 18272 11299 18275
rect 11330 18272 11336 18284
rect 11287 18244 11336 18272
rect 11287 18241 11299 18244
rect 11241 18235 11299 18241
rect 11330 18232 11336 18244
rect 11388 18232 11394 18284
rect 12434 18232 12440 18284
rect 12492 18232 12498 18284
rect 16574 18232 16580 18284
rect 16632 18272 16638 18284
rect 21284 18281 21312 18312
rect 22646 18300 22652 18312
rect 22704 18300 22710 18352
rect 23293 18343 23351 18349
rect 23293 18309 23305 18343
rect 23339 18340 23351 18343
rect 24854 18340 24860 18352
rect 23339 18312 24860 18340
rect 23339 18309 23351 18312
rect 23293 18303 23351 18309
rect 24854 18300 24860 18312
rect 24912 18300 24918 18352
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16632 18244 16865 18272
rect 16632 18232 16638 18244
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 21269 18275 21327 18281
rect 18262 18244 19012 18272
rect 16853 18235 16911 18241
rect 8067 18176 10548 18204
rect 10597 18207 10655 18213
rect 8067 18173 8079 18176
rect 8021 18167 8079 18173
rect 10597 18173 10609 18207
rect 10643 18173 10655 18207
rect 10597 18167 10655 18173
rect 7760 18068 7788 18167
rect 9766 18136 9772 18148
rect 9048 18108 9772 18136
rect 9048 18068 9076 18108
rect 9766 18096 9772 18108
rect 9824 18096 9830 18148
rect 7760 18040 9076 18068
rect 9122 18028 9128 18080
rect 9180 18068 9186 18080
rect 10612 18068 10640 18167
rect 12802 18164 12808 18216
rect 12860 18204 12866 18216
rect 13173 18207 13231 18213
rect 13173 18204 13185 18207
rect 12860 18176 13185 18204
rect 12860 18164 12866 18176
rect 13173 18173 13185 18176
rect 13219 18173 13231 18207
rect 13173 18167 13231 18173
rect 14182 18164 14188 18216
rect 14240 18204 14246 18216
rect 14369 18207 14427 18213
rect 14369 18204 14381 18207
rect 14240 18176 14381 18204
rect 14240 18164 14246 18176
rect 14369 18173 14381 18176
rect 14415 18173 14427 18207
rect 14369 18167 14427 18173
rect 16666 18164 16672 18216
rect 16724 18204 16730 18216
rect 17129 18207 17187 18213
rect 17129 18204 17141 18207
rect 16724 18176 17141 18204
rect 16724 18164 16730 18176
rect 17129 18173 17141 18176
rect 17175 18204 17187 18207
rect 18690 18204 18696 18216
rect 17175 18176 18696 18204
rect 17175 18173 17187 18176
rect 17129 18167 17187 18173
rect 18690 18164 18696 18176
rect 18748 18164 18754 18216
rect 10870 18096 10876 18148
rect 10928 18136 10934 18148
rect 18984 18145 19012 18244
rect 21269 18241 21281 18275
rect 21315 18241 21327 18275
rect 21269 18235 21327 18241
rect 22094 18232 22100 18284
rect 22152 18232 22158 18284
rect 23474 18232 23480 18284
rect 23532 18272 23538 18284
rect 23937 18275 23995 18281
rect 23937 18272 23949 18275
rect 23532 18244 23949 18272
rect 23532 18232 23538 18244
rect 23937 18241 23949 18244
rect 23983 18241 23995 18275
rect 23937 18235 23995 18241
rect 24670 18164 24676 18216
rect 24728 18164 24734 18216
rect 13817 18139 13875 18145
rect 13817 18136 13829 18139
rect 10928 18108 13829 18136
rect 10928 18096 10934 18108
rect 13817 18105 13829 18108
rect 13863 18105 13875 18139
rect 13817 18099 13875 18105
rect 18969 18139 19027 18145
rect 18969 18105 18981 18139
rect 19015 18136 19027 18139
rect 20806 18136 20812 18148
rect 19015 18108 20812 18136
rect 19015 18105 19027 18108
rect 18969 18099 19027 18105
rect 20806 18096 20812 18108
rect 20864 18096 20870 18148
rect 9180 18040 10640 18068
rect 9180 18028 9186 18040
rect 11054 18028 11060 18080
rect 11112 18028 11118 18080
rect 18322 18028 18328 18080
rect 18380 18068 18386 18080
rect 18601 18071 18659 18077
rect 18601 18068 18613 18071
rect 18380 18040 18613 18068
rect 18380 18028 18386 18040
rect 18601 18037 18613 18040
rect 18647 18037 18659 18071
rect 18601 18031 18659 18037
rect 21082 18028 21088 18080
rect 21140 18028 21146 18080
rect 1104 17978 25852 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 25852 17978
rect 1104 17904 25852 17926
rect 7650 17824 7656 17876
rect 7708 17864 7714 17876
rect 7837 17867 7895 17873
rect 7837 17864 7849 17867
rect 7708 17836 7849 17864
rect 7708 17824 7714 17836
rect 7837 17833 7849 17836
rect 7883 17833 7895 17867
rect 7837 17827 7895 17833
rect 12253 17867 12311 17873
rect 12253 17833 12265 17867
rect 12299 17864 12311 17867
rect 15194 17864 15200 17876
rect 12299 17836 15200 17864
rect 12299 17833 12311 17836
rect 12253 17827 12311 17833
rect 15194 17824 15200 17836
rect 15252 17824 15258 17876
rect 20714 17824 20720 17876
rect 20772 17864 20778 17876
rect 24026 17864 24032 17876
rect 20772 17836 24032 17864
rect 20772 17824 20778 17836
rect 24026 17824 24032 17836
rect 24084 17824 24090 17876
rect 13814 17796 13820 17808
rect 12728 17768 13820 17796
rect 7834 17688 7840 17740
rect 7892 17728 7898 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 7892 17700 8401 17728
rect 7892 17688 7898 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 11698 17688 11704 17740
rect 11756 17728 11762 17740
rect 11793 17731 11851 17737
rect 11793 17728 11805 17731
rect 11756 17700 11805 17728
rect 11756 17688 11762 17700
rect 11793 17697 11805 17700
rect 11839 17697 11851 17731
rect 11793 17691 11851 17697
rect 11974 17688 11980 17740
rect 12032 17728 12038 17740
rect 12728 17737 12756 17768
rect 13814 17756 13820 17768
rect 13872 17756 13878 17808
rect 16298 17796 16304 17808
rect 16132 17768 16304 17796
rect 12713 17731 12771 17737
rect 12713 17728 12725 17731
rect 12032 17700 12725 17728
rect 12032 17688 12038 17700
rect 12713 17697 12725 17700
rect 12759 17697 12771 17731
rect 12713 17691 12771 17697
rect 12897 17731 12955 17737
rect 12897 17697 12909 17731
rect 12943 17728 12955 17731
rect 13354 17728 13360 17740
rect 12943 17700 13360 17728
rect 12943 17697 12955 17700
rect 12897 17691 12955 17697
rect 13354 17688 13360 17700
rect 13412 17688 13418 17740
rect 16132 17737 16160 17768
rect 16298 17756 16304 17768
rect 16356 17756 16362 17808
rect 17218 17756 17224 17808
rect 17276 17796 17282 17808
rect 17862 17796 17868 17808
rect 17276 17768 17868 17796
rect 17276 17756 17282 17768
rect 17862 17756 17868 17768
rect 17920 17756 17926 17808
rect 18322 17756 18328 17808
rect 18380 17796 18386 17808
rect 20625 17799 20683 17805
rect 18380 17768 20024 17796
rect 18380 17756 18386 17768
rect 16117 17731 16175 17737
rect 16117 17697 16129 17731
rect 16163 17697 16175 17731
rect 16117 17691 16175 17697
rect 17586 17688 17592 17740
rect 17644 17728 17650 17740
rect 17957 17731 18015 17737
rect 17957 17728 17969 17731
rect 17644 17700 17969 17728
rect 17644 17688 17650 17700
rect 17957 17697 17969 17700
rect 18003 17697 18015 17731
rect 17957 17691 18015 17697
rect 18874 17688 18880 17740
rect 18932 17728 18938 17740
rect 19996 17737 20024 17768
rect 20625 17765 20637 17799
rect 20671 17796 20683 17799
rect 21542 17796 21548 17808
rect 20671 17768 21548 17796
rect 20671 17765 20683 17768
rect 20625 17759 20683 17765
rect 21542 17756 21548 17768
rect 21600 17756 21606 17808
rect 25682 17796 25688 17808
rect 22066 17768 25688 17796
rect 19889 17731 19947 17737
rect 19889 17728 19901 17731
rect 18932 17700 19901 17728
rect 18932 17688 18938 17700
rect 19889 17697 19901 17700
rect 19935 17697 19947 17731
rect 19889 17691 19947 17697
rect 19981 17731 20039 17737
rect 19981 17697 19993 17731
rect 20027 17697 20039 17731
rect 19981 17691 20039 17697
rect 9766 17620 9772 17672
rect 9824 17620 9830 17672
rect 12621 17663 12679 17669
rect 12621 17629 12633 17663
rect 12667 17660 12679 17663
rect 14274 17660 14280 17672
rect 12667 17632 14280 17660
rect 12667 17629 12679 17632
rect 12621 17623 12679 17629
rect 14274 17620 14280 17632
rect 14332 17620 14338 17672
rect 15746 17620 15752 17672
rect 15804 17660 15810 17672
rect 16393 17663 16451 17669
rect 16393 17660 16405 17663
rect 15804 17632 16405 17660
rect 15804 17620 15810 17632
rect 16393 17629 16405 17632
rect 16439 17629 16451 17663
rect 16393 17623 16451 17629
rect 16942 17620 16948 17672
rect 17000 17660 17006 17672
rect 18417 17663 18475 17669
rect 18417 17660 18429 17663
rect 17000 17632 18429 17660
rect 17000 17620 17006 17632
rect 18417 17629 18429 17632
rect 18463 17629 18475 17663
rect 18417 17623 18475 17629
rect 19334 17620 19340 17672
rect 19392 17660 19398 17672
rect 20809 17663 20867 17669
rect 20809 17660 20821 17663
rect 19392 17632 20821 17660
rect 19392 17620 19398 17632
rect 20809 17629 20821 17632
rect 20855 17629 20867 17663
rect 20809 17623 20867 17629
rect 21450 17620 21456 17672
rect 21508 17620 21514 17672
rect 22066 17604 22094 17768
rect 25682 17756 25688 17768
rect 25740 17756 25746 17808
rect 23845 17731 23903 17737
rect 23845 17697 23857 17731
rect 23891 17728 23903 17731
rect 24854 17728 24860 17740
rect 23891 17700 24860 17728
rect 23891 17697 23903 17700
rect 23845 17691 23903 17697
rect 24854 17688 24860 17700
rect 24912 17688 24918 17740
rect 24946 17688 24952 17740
rect 25004 17728 25010 17740
rect 25041 17731 25099 17737
rect 25041 17728 25053 17731
rect 25004 17700 25053 17728
rect 25004 17688 25010 17700
rect 25041 17697 25053 17700
rect 25087 17697 25099 17731
rect 25041 17691 25099 17697
rect 25130 17688 25136 17740
rect 25188 17688 25194 17740
rect 22830 17620 22836 17672
rect 22888 17620 22894 17672
rect 8205 17595 8263 17601
rect 8205 17561 8217 17595
rect 8251 17592 8263 17595
rect 8846 17592 8852 17604
rect 8251 17564 8852 17592
rect 8251 17561 8263 17564
rect 8205 17555 8263 17561
rect 8846 17552 8852 17564
rect 8904 17552 8910 17604
rect 9950 17552 9956 17604
rect 10008 17592 10014 17604
rect 10045 17595 10103 17601
rect 10045 17592 10057 17595
rect 10008 17564 10057 17592
rect 10008 17552 10014 17564
rect 10045 17561 10057 17564
rect 10091 17561 10103 17595
rect 10045 17555 10103 17561
rect 11054 17552 11060 17604
rect 11112 17552 11118 17604
rect 13722 17552 13728 17604
rect 13780 17592 13786 17604
rect 14185 17595 14243 17601
rect 14185 17592 14197 17595
rect 13780 17564 14197 17592
rect 13780 17552 13786 17564
rect 14185 17561 14197 17564
rect 14231 17592 14243 17595
rect 16850 17592 16856 17604
rect 14231 17564 16856 17592
rect 14231 17561 14243 17564
rect 14185 17555 14243 17561
rect 16850 17552 16856 17564
rect 16908 17592 16914 17604
rect 17678 17592 17684 17604
rect 16908 17564 17684 17592
rect 16908 17552 16914 17564
rect 17678 17552 17684 17564
rect 17736 17552 17742 17604
rect 17770 17552 17776 17604
rect 17828 17592 17834 17604
rect 18785 17595 18843 17601
rect 18785 17592 18797 17595
rect 17828 17564 18797 17592
rect 17828 17552 17834 17564
rect 18785 17561 18797 17564
rect 18831 17561 18843 17595
rect 18785 17555 18843 17561
rect 19444 17564 20576 17592
rect 7190 17484 7196 17536
rect 7248 17484 7254 17536
rect 7650 17484 7656 17536
rect 7708 17524 7714 17536
rect 8297 17527 8355 17533
rect 8297 17524 8309 17527
rect 7708 17496 8309 17524
rect 7708 17484 7714 17496
rect 8297 17493 8309 17496
rect 8343 17493 8355 17527
rect 8297 17487 8355 17493
rect 9125 17527 9183 17533
rect 9125 17493 9137 17527
rect 9171 17524 9183 17527
rect 9398 17524 9404 17536
rect 9171 17496 9404 17524
rect 9171 17493 9183 17496
rect 9125 17487 9183 17493
rect 9398 17484 9404 17496
rect 9456 17484 9462 17536
rect 13170 17484 13176 17536
rect 13228 17524 13234 17536
rect 13449 17527 13507 17533
rect 13449 17524 13461 17527
rect 13228 17496 13461 17524
rect 13228 17484 13234 17496
rect 13449 17493 13461 17496
rect 13495 17493 13507 17527
rect 13449 17487 13507 17493
rect 15470 17484 15476 17536
rect 15528 17484 15534 17536
rect 17402 17484 17408 17536
rect 17460 17484 17466 17536
rect 17862 17484 17868 17536
rect 17920 17524 17926 17536
rect 18690 17524 18696 17536
rect 17920 17496 18696 17524
rect 17920 17484 17926 17496
rect 18690 17484 18696 17496
rect 18748 17484 18754 17536
rect 19444 17533 19472 17564
rect 19429 17527 19487 17533
rect 19429 17493 19441 17527
rect 19475 17493 19487 17527
rect 19429 17487 19487 17493
rect 19797 17527 19855 17533
rect 19797 17493 19809 17527
rect 19843 17524 19855 17527
rect 19886 17524 19892 17536
rect 19843 17496 19892 17524
rect 19843 17493 19855 17496
rect 19797 17487 19855 17493
rect 19886 17484 19892 17496
rect 19944 17484 19950 17536
rect 20548 17524 20576 17564
rect 22002 17552 22008 17604
rect 22060 17564 22094 17604
rect 22060 17552 22066 17564
rect 22186 17552 22192 17604
rect 22244 17552 22250 17604
rect 25038 17592 25044 17604
rect 23584 17564 25044 17592
rect 21082 17524 21088 17536
rect 20548 17496 21088 17524
rect 21082 17484 21088 17496
rect 21140 17484 21146 17536
rect 21269 17527 21327 17533
rect 21269 17493 21281 17527
rect 21315 17524 21327 17527
rect 23584 17524 23612 17564
rect 25038 17552 25044 17564
rect 25096 17552 25102 17604
rect 21315 17496 23612 17524
rect 21315 17493 21327 17496
rect 21269 17487 21327 17493
rect 23750 17484 23756 17536
rect 23808 17524 23814 17536
rect 24581 17527 24639 17533
rect 24581 17524 24593 17527
rect 23808 17496 24593 17524
rect 23808 17484 23814 17496
rect 24581 17493 24593 17496
rect 24627 17493 24639 17527
rect 24581 17487 24639 17493
rect 24670 17484 24676 17536
rect 24728 17524 24734 17536
rect 24949 17527 25007 17533
rect 24949 17524 24961 17527
rect 24728 17496 24961 17524
rect 24728 17484 24734 17496
rect 24949 17493 24961 17496
rect 24995 17493 25007 17527
rect 24949 17487 25007 17493
rect 1104 17434 25852 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 25852 17434
rect 1104 17360 25852 17382
rect 7190 17280 7196 17332
rect 7248 17320 7254 17332
rect 8021 17323 8079 17329
rect 8021 17320 8033 17323
rect 7248 17292 8033 17320
rect 7248 17280 7254 17292
rect 8021 17289 8033 17292
rect 8067 17289 8079 17323
rect 8021 17283 8079 17289
rect 9033 17323 9091 17329
rect 9033 17289 9045 17323
rect 9079 17320 9091 17323
rect 9214 17320 9220 17332
rect 9079 17292 9220 17320
rect 9079 17289 9091 17292
rect 9033 17283 9091 17289
rect 9214 17280 9220 17292
rect 9272 17280 9278 17332
rect 9398 17280 9404 17332
rect 9456 17280 9462 17332
rect 11514 17280 11520 17332
rect 11572 17320 11578 17332
rect 12434 17320 12440 17332
rect 11572 17292 12440 17320
rect 11572 17280 11578 17292
rect 12434 17280 12440 17292
rect 12492 17320 12498 17332
rect 13722 17320 13728 17332
rect 12492 17292 13728 17320
rect 12492 17280 12498 17292
rect 13722 17280 13728 17292
rect 13780 17280 13786 17332
rect 16390 17320 16396 17332
rect 14660 17292 16396 17320
rect 9766 17212 9772 17264
rect 9824 17252 9830 17264
rect 10965 17255 11023 17261
rect 10965 17252 10977 17255
rect 9824 17224 10977 17252
rect 9824 17212 9830 17224
rect 10965 17221 10977 17224
rect 11011 17221 11023 17255
rect 10965 17215 11023 17221
rect 13170 17212 13176 17264
rect 13228 17212 13234 17264
rect 14660 17252 14688 17292
rect 16390 17280 16396 17292
rect 16448 17320 16454 17332
rect 16574 17320 16580 17332
rect 16448 17292 16580 17320
rect 16448 17280 16454 17292
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 17497 17323 17555 17329
rect 17497 17289 17509 17323
rect 17543 17320 17555 17323
rect 17586 17320 17592 17332
rect 17543 17292 17592 17320
rect 17543 17289 17555 17292
rect 17497 17283 17555 17289
rect 17586 17280 17592 17292
rect 17644 17280 17650 17332
rect 20162 17280 20168 17332
rect 20220 17320 20226 17332
rect 20349 17323 20407 17329
rect 20349 17320 20361 17323
rect 20220 17292 20361 17320
rect 20220 17280 20226 17292
rect 20349 17289 20361 17292
rect 20395 17289 20407 17323
rect 20349 17283 20407 17289
rect 22002 17280 22008 17332
rect 22060 17280 22066 17332
rect 22741 17323 22799 17329
rect 22741 17289 22753 17323
rect 22787 17320 22799 17323
rect 24486 17320 24492 17332
rect 22787 17292 24492 17320
rect 22787 17289 22799 17292
rect 22741 17283 22799 17289
rect 24486 17280 24492 17292
rect 24544 17280 24550 17332
rect 14568 17224 14688 17252
rect 10229 17187 10287 17193
rect 10229 17153 10241 17187
rect 10275 17184 10287 17187
rect 11514 17184 11520 17196
rect 10275 17156 11520 17184
rect 10275 17153 10287 17156
rect 10229 17147 10287 17153
rect 11514 17144 11520 17156
rect 11572 17144 11578 17196
rect 14568 17193 14596 17224
rect 16942 17212 16948 17264
rect 17000 17212 17006 17264
rect 17957 17255 18015 17261
rect 17957 17221 17969 17255
rect 18003 17252 18015 17255
rect 18966 17252 18972 17264
rect 18003 17224 18972 17252
rect 18003 17221 18015 17224
rect 17957 17215 18015 17221
rect 18966 17212 18972 17224
rect 19024 17212 19030 17264
rect 20717 17255 20775 17261
rect 20717 17252 20729 17255
rect 20102 17224 20729 17252
rect 20717 17221 20729 17224
rect 20763 17252 20775 17255
rect 20806 17252 20812 17264
rect 20763 17224 20812 17252
rect 20763 17221 20775 17224
rect 20717 17215 20775 17221
rect 20806 17212 20812 17224
rect 20864 17252 20870 17264
rect 21818 17252 21824 17264
rect 20864 17224 21824 17252
rect 20864 17212 20870 17224
rect 21818 17212 21824 17224
rect 21876 17212 21882 17264
rect 23658 17212 23664 17264
rect 23716 17252 23722 17264
rect 23753 17255 23811 17261
rect 23753 17252 23765 17255
rect 23716 17224 23765 17252
rect 23716 17212 23722 17224
rect 23753 17221 23765 17224
rect 23799 17221 23811 17255
rect 23753 17215 23811 17221
rect 14553 17187 14611 17193
rect 14553 17153 14565 17187
rect 14599 17153 14611 17187
rect 21269 17187 21327 17193
rect 15962 17156 16988 17184
rect 14553 17147 14611 17153
rect 16960 17128 16988 17156
rect 21269 17153 21281 17187
rect 21315 17184 21327 17187
rect 22649 17187 22707 17193
rect 22649 17184 22661 17187
rect 21315 17156 22661 17184
rect 21315 17153 21327 17156
rect 21269 17147 21327 17153
rect 22649 17153 22661 17156
rect 22695 17153 22707 17187
rect 22649 17147 22707 17153
rect 23474 17144 23480 17196
rect 23532 17144 23538 17196
rect 24854 17144 24860 17196
rect 24912 17144 24918 17196
rect 8113 17119 8171 17125
rect 8113 17085 8125 17119
rect 8159 17085 8171 17119
rect 8113 17079 8171 17085
rect 8297 17119 8355 17125
rect 8297 17085 8309 17119
rect 8343 17116 8355 17119
rect 8570 17116 8576 17128
rect 8343 17088 8576 17116
rect 8343 17085 8355 17088
rect 8297 17079 8355 17085
rect 7558 17008 7564 17060
rect 7616 17048 7622 17060
rect 7653 17051 7711 17057
rect 7653 17048 7665 17051
rect 7616 17020 7665 17048
rect 7616 17008 7622 17020
rect 7653 17017 7665 17020
rect 7699 17017 7711 17051
rect 7653 17011 7711 17017
rect 3326 16940 3332 16992
rect 3384 16980 3390 16992
rect 7285 16983 7343 16989
rect 7285 16980 7297 16983
rect 3384 16952 7297 16980
rect 3384 16940 3390 16952
rect 7285 16949 7297 16952
rect 7331 16980 7343 16983
rect 8128 16980 8156 17079
rect 8570 17076 8576 17088
rect 8628 17076 8634 17128
rect 8757 17119 8815 17125
rect 8757 17085 8769 17119
rect 8803 17116 8815 17119
rect 9398 17116 9404 17128
rect 8803 17088 9404 17116
rect 8803 17085 8815 17088
rect 8757 17079 8815 17085
rect 9398 17076 9404 17088
rect 9456 17116 9462 17128
rect 9493 17119 9551 17125
rect 9493 17116 9505 17119
rect 9456 17088 9505 17116
rect 9456 17076 9462 17088
rect 9493 17085 9505 17088
rect 9539 17085 9551 17119
rect 9493 17079 9551 17085
rect 9582 17076 9588 17128
rect 9640 17076 9646 17128
rect 11054 17076 11060 17128
rect 11112 17116 11118 17128
rect 11885 17119 11943 17125
rect 11885 17116 11897 17119
rect 11112 17088 11897 17116
rect 11112 17076 11118 17088
rect 11885 17085 11897 17088
rect 11931 17116 11943 17119
rect 12529 17119 12587 17125
rect 11931 17088 12434 17116
rect 11931 17085 11943 17088
rect 11885 17079 11943 17085
rect 7331 16952 8156 16980
rect 7331 16949 7343 16952
rect 7285 16943 7343 16949
rect 11514 16940 11520 16992
rect 11572 16940 11578 16992
rect 11974 16940 11980 16992
rect 12032 16980 12038 16992
rect 12069 16983 12127 16989
rect 12069 16980 12081 16983
rect 12032 16952 12081 16980
rect 12032 16940 12038 16952
rect 12069 16949 12081 16952
rect 12115 16949 12127 16983
rect 12406 16980 12434 17088
rect 12529 17085 12541 17119
rect 12575 17116 12587 17119
rect 12710 17116 12716 17128
rect 12575 17088 12716 17116
rect 12575 17085 12587 17088
rect 12529 17079 12587 17085
rect 12710 17076 12716 17088
rect 12768 17116 12774 17128
rect 13265 17119 13323 17125
rect 13265 17116 13277 17119
rect 12768 17088 13277 17116
rect 12768 17076 12774 17088
rect 13265 17085 13277 17088
rect 13311 17085 13323 17119
rect 13265 17079 13323 17085
rect 13449 17119 13507 17125
rect 13449 17085 13461 17119
rect 13495 17116 13507 17119
rect 13538 17116 13544 17128
rect 13495 17088 13544 17116
rect 13495 17085 13507 17088
rect 13449 17079 13507 17085
rect 13538 17076 13544 17088
rect 13596 17076 13602 17128
rect 14829 17119 14887 17125
rect 14829 17085 14841 17119
rect 14875 17116 14887 17119
rect 15562 17116 15568 17128
rect 14875 17088 15568 17116
rect 14875 17085 14887 17088
rect 14829 17079 14887 17085
rect 15562 17076 15568 17088
rect 15620 17076 15626 17128
rect 16114 17116 16120 17128
rect 15948 17088 16120 17116
rect 15948 17060 15976 17088
rect 16114 17076 16120 17088
rect 16172 17116 16178 17128
rect 16301 17119 16359 17125
rect 16301 17116 16313 17119
rect 16172 17088 16313 17116
rect 16172 17076 16178 17088
rect 16301 17085 16313 17088
rect 16347 17085 16359 17119
rect 16301 17079 16359 17085
rect 16942 17076 16948 17128
rect 17000 17076 17006 17128
rect 17862 17076 17868 17128
rect 17920 17116 17926 17128
rect 18601 17119 18659 17125
rect 18601 17116 18613 17119
rect 17920 17088 18613 17116
rect 17920 17076 17926 17088
rect 18601 17085 18613 17088
rect 18647 17085 18659 17119
rect 18601 17079 18659 17085
rect 18874 17076 18880 17128
rect 18932 17076 18938 17128
rect 22554 17076 22560 17128
rect 22612 17116 22618 17128
rect 22833 17119 22891 17125
rect 22833 17116 22845 17119
rect 22612 17088 22845 17116
rect 22612 17076 22618 17088
rect 22833 17085 22845 17088
rect 22879 17116 22891 17119
rect 25225 17119 25283 17125
rect 25225 17116 25237 17119
rect 22879 17088 25237 17116
rect 22879 17085 22891 17088
rect 22833 17079 22891 17085
rect 25225 17085 25237 17088
rect 25271 17085 25283 17119
rect 25225 17079 25283 17085
rect 12805 17051 12863 17057
rect 12805 17017 12817 17051
rect 12851 17048 12863 17051
rect 13630 17048 13636 17060
rect 12851 17020 13636 17048
rect 12851 17017 12863 17020
rect 12805 17011 12863 17017
rect 13630 17008 13636 17020
rect 13688 17008 13694 17060
rect 15930 17008 15936 17060
rect 15988 17008 15994 17060
rect 16022 17008 16028 17060
rect 16080 17048 16086 17060
rect 18141 17051 18199 17057
rect 18141 17048 18153 17051
rect 16080 17020 18153 17048
rect 16080 17008 16086 17020
rect 18141 17017 18153 17020
rect 18187 17017 18199 17051
rect 18141 17011 18199 17017
rect 20898 17008 20904 17060
rect 20956 17048 20962 17060
rect 22281 17051 22339 17057
rect 22281 17048 22293 17051
rect 20956 17020 22293 17048
rect 20956 17008 20962 17020
rect 22281 17017 22293 17020
rect 22327 17017 22339 17051
rect 22281 17011 22339 17017
rect 13814 16980 13820 16992
rect 12406 16952 13820 16980
rect 12069 16943 12127 16949
rect 13814 16940 13820 16952
rect 13872 16940 13878 16992
rect 16666 16940 16672 16992
rect 16724 16980 16730 16992
rect 17037 16983 17095 16989
rect 17037 16980 17049 16983
rect 16724 16952 17049 16980
rect 16724 16940 16730 16952
rect 17037 16949 17049 16952
rect 17083 16949 17095 16983
rect 17037 16943 17095 16949
rect 18690 16940 18696 16992
rect 18748 16980 18754 16992
rect 18966 16980 18972 16992
rect 18748 16952 18972 16980
rect 18748 16940 18754 16952
rect 18966 16940 18972 16952
rect 19024 16940 19030 16992
rect 20346 16940 20352 16992
rect 20404 16980 20410 16992
rect 22094 16980 22100 16992
rect 20404 16952 22100 16980
rect 20404 16940 20410 16952
rect 22094 16940 22100 16952
rect 22152 16940 22158 16992
rect 1104 16890 25852 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 25852 16890
rect 1104 16816 25852 16838
rect 8570 16736 8576 16788
rect 8628 16736 8634 16788
rect 11330 16736 11336 16788
rect 11388 16776 11394 16788
rect 11882 16776 11888 16788
rect 11388 16748 11888 16776
rect 11388 16736 11394 16748
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 13909 16779 13967 16785
rect 13909 16745 13921 16779
rect 13955 16776 13967 16779
rect 14642 16776 14648 16788
rect 13955 16748 14648 16776
rect 13955 16745 13967 16748
rect 13909 16739 13967 16745
rect 11606 16708 11612 16720
rect 10704 16680 11612 16708
rect 10704 16649 10732 16680
rect 11606 16668 11612 16680
rect 11664 16668 11670 16720
rect 13814 16708 13820 16720
rect 13464 16680 13820 16708
rect 10689 16643 10747 16649
rect 10689 16609 10701 16643
rect 10735 16609 10747 16643
rect 10689 16603 10747 16609
rect 10873 16643 10931 16649
rect 10873 16609 10885 16643
rect 10919 16640 10931 16643
rect 11330 16640 11336 16652
rect 10919 16612 11336 16640
rect 10919 16609 10931 16612
rect 10873 16603 10931 16609
rect 11330 16600 11336 16612
rect 11388 16600 11394 16652
rect 11793 16643 11851 16649
rect 11793 16609 11805 16643
rect 11839 16640 11851 16643
rect 12802 16640 12808 16652
rect 11839 16612 12808 16640
rect 11839 16609 11851 16612
rect 11793 16603 11851 16609
rect 12802 16600 12808 16612
rect 12860 16600 12866 16652
rect 13464 16572 13492 16680
rect 13814 16668 13820 16680
rect 13872 16708 13878 16720
rect 13924 16708 13952 16739
rect 14642 16736 14648 16748
rect 14700 16776 14706 16788
rect 14700 16748 16896 16776
rect 14700 16736 14706 16748
rect 16482 16708 16488 16720
rect 13872 16680 13952 16708
rect 16316 16680 16488 16708
rect 13872 16668 13878 16680
rect 13538 16600 13544 16652
rect 13596 16640 13602 16652
rect 16316 16649 16344 16680
rect 16482 16668 16488 16680
rect 16540 16668 16546 16720
rect 16868 16717 16896 16748
rect 21818 16736 21824 16788
rect 21876 16776 21882 16788
rect 22281 16779 22339 16785
rect 22281 16776 22293 16779
rect 21876 16748 22293 16776
rect 21876 16736 21882 16748
rect 22281 16745 22293 16748
rect 22327 16745 22339 16779
rect 22281 16739 22339 16745
rect 16853 16711 16911 16717
rect 16853 16677 16865 16711
rect 16899 16708 16911 16711
rect 16942 16708 16948 16720
rect 16899 16680 16948 16708
rect 16899 16677 16911 16680
rect 16853 16671 16911 16677
rect 16942 16668 16948 16680
rect 17000 16668 17006 16720
rect 17770 16668 17776 16720
rect 17828 16708 17834 16720
rect 19794 16708 19800 16720
rect 17828 16680 19800 16708
rect 17828 16668 17834 16680
rect 19794 16668 19800 16680
rect 19852 16668 19858 16720
rect 15105 16643 15163 16649
rect 15105 16640 15117 16643
rect 13596 16612 15117 16640
rect 13596 16600 13602 16612
rect 15105 16609 15117 16612
rect 15151 16609 15163 16643
rect 16301 16643 16359 16649
rect 15105 16603 15163 16609
rect 15396 16612 16252 16640
rect 13630 16572 13636 16584
rect 13202 16544 13636 16572
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 15396 16572 15424 16612
rect 14568 16544 15424 16572
rect 10318 16504 10324 16516
rect 9876 16476 10324 16504
rect 9876 16448 9904 16476
rect 10318 16464 10324 16476
rect 10376 16504 10382 16516
rect 10597 16507 10655 16513
rect 10597 16504 10609 16507
rect 10376 16476 10609 16504
rect 10376 16464 10382 16476
rect 10597 16473 10609 16476
rect 10643 16473 10655 16507
rect 10597 16467 10655 16473
rect 12069 16507 12127 16513
rect 12069 16473 12081 16507
rect 12115 16473 12127 16507
rect 14366 16504 14372 16516
rect 12069 16467 12127 16473
rect 13464 16476 14372 16504
rect 9858 16396 9864 16448
rect 9916 16396 9922 16448
rect 10226 16396 10232 16448
rect 10284 16396 10290 16448
rect 12084 16436 12112 16467
rect 13464 16436 13492 16476
rect 14366 16464 14372 16476
rect 14424 16464 14430 16516
rect 12084 16408 13492 16436
rect 13538 16396 13544 16448
rect 13596 16396 13602 16448
rect 14274 16396 14280 16448
rect 14332 16396 14338 16448
rect 14568 16445 14596 16544
rect 15470 16532 15476 16584
rect 15528 16572 15534 16584
rect 16117 16575 16175 16581
rect 16117 16572 16129 16575
rect 15528 16544 16129 16572
rect 15528 16532 15534 16544
rect 16117 16541 16129 16544
rect 16163 16541 16175 16575
rect 16224 16572 16252 16612
rect 16301 16609 16313 16643
rect 16347 16609 16359 16643
rect 16301 16603 16359 16609
rect 16390 16600 16396 16652
rect 16448 16640 16454 16652
rect 17862 16640 17868 16652
rect 16448 16612 17868 16640
rect 16448 16600 16454 16612
rect 17862 16600 17868 16612
rect 17920 16640 17926 16652
rect 17957 16643 18015 16649
rect 17957 16640 17969 16643
rect 17920 16612 17969 16640
rect 17920 16600 17926 16612
rect 17957 16609 17969 16612
rect 18003 16609 18015 16643
rect 17957 16603 18015 16609
rect 20254 16600 20260 16652
rect 20312 16600 20318 16652
rect 22020 16612 22140 16640
rect 18877 16575 18935 16581
rect 18877 16572 18889 16575
rect 16224 16544 18889 16572
rect 16117 16535 16175 16541
rect 18877 16541 18889 16544
rect 18923 16541 18935 16575
rect 18877 16535 18935 16541
rect 19797 16575 19855 16581
rect 19797 16541 19809 16575
rect 19843 16541 19855 16575
rect 22020 16572 22048 16612
rect 19797 16535 19855 16541
rect 21928 16544 22048 16572
rect 22112 16572 22140 16612
rect 22370 16572 22376 16584
rect 22112 16544 22376 16572
rect 14921 16507 14979 16513
rect 14921 16473 14933 16507
rect 14967 16504 14979 16507
rect 15654 16504 15660 16516
rect 14967 16476 15660 16504
rect 14967 16473 14979 16476
rect 14921 16467 14979 16473
rect 15654 16464 15660 16476
rect 15712 16464 15718 16516
rect 16850 16464 16856 16516
rect 16908 16504 16914 16516
rect 17221 16507 17279 16513
rect 17221 16504 17233 16507
rect 16908 16476 17233 16504
rect 16908 16464 16914 16476
rect 17221 16473 17233 16476
rect 17267 16504 17279 16507
rect 17267 16476 19288 16504
rect 17267 16473 17279 16476
rect 17221 16467 17279 16473
rect 14553 16439 14611 16445
rect 14553 16405 14565 16439
rect 14599 16405 14611 16439
rect 14553 16399 14611 16405
rect 15010 16396 15016 16448
rect 15068 16396 15074 16448
rect 15749 16439 15807 16445
rect 15749 16405 15761 16439
rect 15795 16436 15807 16439
rect 15838 16436 15844 16448
rect 15795 16408 15844 16436
rect 15795 16405 15807 16408
rect 15749 16399 15807 16405
rect 15838 16396 15844 16408
rect 15896 16396 15902 16448
rect 16206 16396 16212 16448
rect 16264 16396 16270 16448
rect 18690 16396 18696 16448
rect 18748 16396 18754 16448
rect 19260 16445 19288 16476
rect 19245 16439 19303 16445
rect 19245 16405 19257 16439
rect 19291 16436 19303 16439
rect 19426 16436 19432 16448
rect 19291 16408 19432 16436
rect 19291 16405 19303 16408
rect 19245 16399 19303 16405
rect 19426 16396 19432 16408
rect 19484 16396 19490 16448
rect 19518 16396 19524 16448
rect 19576 16436 19582 16448
rect 19613 16439 19671 16445
rect 19613 16436 19625 16439
rect 19576 16408 19625 16436
rect 19576 16396 19582 16408
rect 19613 16405 19625 16408
rect 19659 16405 19671 16439
rect 19812 16436 19840 16535
rect 20438 16464 20444 16516
rect 20496 16504 20502 16516
rect 20533 16507 20591 16513
rect 20533 16504 20545 16507
rect 20496 16476 20545 16504
rect 20496 16464 20502 16476
rect 20533 16473 20545 16476
rect 20579 16473 20591 16507
rect 21818 16504 21824 16516
rect 21758 16476 21824 16504
rect 20533 16467 20591 16473
rect 21818 16464 21824 16476
rect 21876 16464 21882 16516
rect 21928 16436 21956 16544
rect 22370 16532 22376 16544
rect 22428 16532 22434 16584
rect 22646 16532 22652 16584
rect 22704 16532 22710 16584
rect 23382 16532 23388 16584
rect 23440 16572 23446 16584
rect 23569 16575 23627 16581
rect 23569 16572 23581 16575
rect 23440 16544 23581 16572
rect 23440 16532 23446 16544
rect 23569 16541 23581 16544
rect 23615 16541 23627 16575
rect 23569 16535 23627 16541
rect 24762 16532 24768 16584
rect 24820 16532 24826 16584
rect 22278 16464 22284 16516
rect 22336 16504 22342 16516
rect 23842 16504 23848 16516
rect 22336 16476 23848 16504
rect 22336 16464 22342 16476
rect 23842 16464 23848 16476
rect 23900 16464 23906 16516
rect 24210 16464 24216 16516
rect 24268 16504 24274 16516
rect 24854 16504 24860 16516
rect 24268 16476 24860 16504
rect 24268 16464 24274 16476
rect 24854 16464 24860 16476
rect 24912 16504 24918 16516
rect 25409 16507 25467 16513
rect 25409 16504 25421 16507
rect 24912 16476 25421 16504
rect 24912 16464 24918 16476
rect 25409 16473 25421 16476
rect 25455 16473 25467 16507
rect 25409 16467 25467 16473
rect 19812 16408 21956 16436
rect 22005 16439 22063 16445
rect 19613 16399 19671 16405
rect 22005 16405 22017 16439
rect 22051 16436 22063 16439
rect 22094 16436 22100 16448
rect 22051 16408 22100 16436
rect 22051 16405 22063 16408
rect 22005 16399 22063 16405
rect 22094 16396 22100 16408
rect 22152 16436 22158 16448
rect 22370 16436 22376 16448
rect 22152 16408 22376 16436
rect 22152 16396 22158 16408
rect 22370 16396 22376 16408
rect 22428 16396 22434 16448
rect 22830 16396 22836 16448
rect 22888 16436 22894 16448
rect 24581 16439 24639 16445
rect 24581 16436 24593 16439
rect 22888 16408 24593 16436
rect 22888 16396 22894 16408
rect 24581 16405 24593 16408
rect 24627 16405 24639 16439
rect 24581 16399 24639 16405
rect 1104 16346 25852 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 25852 16346
rect 1104 16272 25852 16294
rect 8294 16192 8300 16244
rect 8352 16232 8358 16244
rect 9306 16232 9312 16244
rect 8352 16204 9312 16232
rect 8352 16192 8358 16204
rect 9306 16192 9312 16204
rect 9364 16192 9370 16244
rect 11606 16192 11612 16244
rect 11664 16232 11670 16244
rect 13357 16235 13415 16241
rect 13357 16232 13369 16235
rect 11664 16204 13369 16232
rect 11664 16192 11670 16204
rect 13357 16201 13369 16204
rect 13403 16201 13415 16235
rect 13357 16195 13415 16201
rect 14553 16235 14611 16241
rect 14553 16201 14565 16235
rect 14599 16232 14611 16235
rect 15010 16232 15016 16244
rect 14599 16204 15016 16232
rect 14599 16201 14611 16204
rect 14553 16195 14611 16201
rect 15010 16192 15016 16204
rect 15068 16192 15074 16244
rect 15654 16192 15660 16244
rect 15712 16232 15718 16244
rect 15749 16235 15807 16241
rect 15749 16232 15761 16235
rect 15712 16204 15761 16232
rect 15712 16192 15718 16204
rect 15749 16201 15761 16204
rect 15795 16201 15807 16235
rect 15749 16195 15807 16201
rect 16206 16192 16212 16244
rect 16264 16192 16270 16244
rect 16850 16192 16856 16244
rect 16908 16192 16914 16244
rect 18690 16192 18696 16244
rect 18748 16232 18754 16244
rect 24762 16232 24768 16244
rect 18748 16204 24768 16232
rect 18748 16192 18754 16204
rect 24762 16192 24768 16204
rect 24820 16192 24826 16244
rect 8386 16164 8392 16176
rect 8050 16136 8392 16164
rect 8386 16124 8392 16136
rect 8444 16164 8450 16176
rect 8573 16167 8631 16173
rect 8573 16164 8585 16167
rect 8444 16136 8585 16164
rect 8444 16124 8450 16136
rect 8573 16133 8585 16136
rect 8619 16164 8631 16167
rect 8662 16164 8668 16176
rect 8619 16136 8668 16164
rect 8619 16133 8631 16136
rect 8573 16127 8631 16133
rect 8662 16124 8668 16136
rect 8720 16124 8726 16176
rect 11698 16124 11704 16176
rect 11756 16164 11762 16176
rect 11793 16167 11851 16173
rect 11793 16164 11805 16167
rect 11756 16136 11805 16164
rect 11756 16124 11762 16136
rect 11793 16133 11805 16136
rect 11839 16133 11851 16167
rect 11793 16127 11851 16133
rect 6546 16056 6552 16108
rect 6604 16056 6610 16108
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 8386 16028 8392 16040
rect 6871 16000 8392 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 8386 15988 8392 16000
rect 8444 16028 8450 16040
rect 9582 16028 9588 16040
rect 8444 16000 9588 16028
rect 8444 15988 8450 16000
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 11808 16028 11836 16127
rect 12710 16124 12716 16176
rect 12768 16164 12774 16176
rect 13817 16167 13875 16173
rect 13817 16164 13829 16167
rect 12768 16136 13829 16164
rect 12768 16124 12774 16136
rect 13817 16133 13829 16136
rect 13863 16133 13875 16167
rect 13817 16127 13875 16133
rect 14366 16124 14372 16176
rect 14424 16164 14430 16176
rect 14424 16136 15148 16164
rect 14424 16124 14430 16136
rect 12434 16056 12440 16108
rect 12492 16096 12498 16108
rect 12529 16099 12587 16105
rect 12529 16096 12541 16099
rect 12492 16068 12541 16096
rect 12492 16056 12498 16068
rect 12529 16065 12541 16068
rect 12575 16065 12587 16099
rect 12529 16059 12587 16065
rect 12621 16099 12679 16105
rect 12621 16065 12633 16099
rect 12667 16096 12679 16099
rect 13725 16099 13783 16105
rect 12667 16068 13308 16096
rect 12667 16065 12679 16068
rect 12621 16059 12679 16065
rect 12250 16028 12256 16040
rect 11808 16000 12256 16028
rect 12250 15988 12256 16000
rect 12308 16028 12314 16040
rect 12713 16031 12771 16037
rect 12308 16000 12434 16028
rect 12308 15988 12314 16000
rect 12066 15920 12072 15972
rect 12124 15960 12130 15972
rect 12161 15963 12219 15969
rect 12161 15960 12173 15963
rect 12124 15932 12173 15960
rect 12124 15920 12130 15932
rect 12161 15929 12173 15932
rect 12207 15929 12219 15963
rect 12406 15960 12434 16000
rect 12713 15997 12725 16031
rect 12759 15997 12771 16031
rect 12713 15991 12771 15997
rect 12728 15960 12756 15991
rect 12406 15932 12756 15960
rect 12161 15923 12219 15929
rect 5166 15852 5172 15904
rect 5224 15892 5230 15904
rect 11974 15892 11980 15904
rect 5224 15864 11980 15892
rect 5224 15852 5230 15864
rect 11974 15852 11980 15864
rect 12032 15852 12038 15904
rect 13280 15892 13308 16068
rect 13725 16065 13737 16099
rect 13771 16096 13783 16099
rect 14274 16096 14280 16108
rect 13771 16068 14280 16096
rect 13771 16065 13783 16068
rect 13725 16059 13783 16065
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 14734 16056 14740 16108
rect 14792 16096 14798 16108
rect 14921 16099 14979 16105
rect 14921 16096 14933 16099
rect 14792 16068 14933 16096
rect 14792 16056 14798 16068
rect 14921 16065 14933 16068
rect 14967 16065 14979 16099
rect 14921 16059 14979 16065
rect 14001 16031 14059 16037
rect 14001 15997 14013 16031
rect 14047 16028 14059 16031
rect 14366 16028 14372 16040
rect 14047 16000 14372 16028
rect 14047 15997 14059 16000
rect 14001 15991 14059 15997
rect 14366 15988 14372 16000
rect 14424 15988 14430 16040
rect 15010 15988 15016 16040
rect 15068 15988 15074 16040
rect 15120 16037 15148 16136
rect 17218 16124 17224 16176
rect 17276 16124 17282 16176
rect 19334 16164 19340 16176
rect 18708 16136 19340 16164
rect 18708 16105 18736 16136
rect 19334 16124 19340 16136
rect 19392 16124 19398 16176
rect 20073 16167 20131 16173
rect 20073 16133 20085 16167
rect 20119 16164 20131 16167
rect 20254 16164 20260 16176
rect 20119 16136 20260 16164
rect 20119 16133 20131 16136
rect 20073 16127 20131 16133
rect 20254 16124 20260 16136
rect 20312 16164 20318 16176
rect 20312 16136 21220 16164
rect 20312 16124 20318 16136
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16065 18107 16099
rect 18049 16059 18107 16065
rect 18693 16099 18751 16105
rect 18693 16065 18705 16099
rect 18739 16065 18751 16099
rect 18693 16059 18751 16065
rect 19245 16099 19303 16105
rect 19245 16065 19257 16099
rect 19291 16096 19303 16099
rect 19426 16096 19432 16108
rect 19291 16068 19432 16096
rect 19291 16065 19303 16068
rect 19245 16059 19303 16065
rect 15105 16031 15163 16037
rect 15105 15997 15117 16031
rect 15151 15997 15163 16031
rect 18064 16028 18092 16059
rect 19426 16056 19432 16068
rect 19484 16056 19490 16108
rect 19794 16056 19800 16108
rect 19852 16096 19858 16108
rect 21085 16099 21143 16105
rect 21085 16096 21097 16099
rect 19852 16068 21097 16096
rect 19852 16056 19858 16068
rect 21085 16065 21097 16068
rect 21131 16065 21143 16099
rect 21192 16096 21220 16136
rect 21818 16124 21824 16176
rect 21876 16164 21882 16176
rect 21876 16136 22770 16164
rect 21876 16124 21882 16136
rect 22005 16099 22063 16105
rect 22005 16096 22017 16099
rect 21192 16068 22017 16096
rect 21085 16059 21143 16065
rect 22005 16065 22017 16068
rect 22051 16065 22063 16099
rect 22005 16059 22063 16065
rect 18782 16028 18788 16040
rect 18064 16000 18788 16028
rect 15105 15991 15163 15997
rect 18782 15988 18788 16000
rect 18840 15988 18846 16040
rect 21174 15988 21180 16040
rect 21232 15988 21238 16040
rect 21358 15988 21364 16040
rect 21416 15988 21422 16040
rect 14274 15920 14280 15972
rect 14332 15960 14338 15972
rect 18690 15960 18696 15972
rect 14332 15932 18696 15960
rect 14332 15920 14338 15932
rect 18690 15920 18696 15932
rect 18748 15920 18754 15972
rect 19150 15920 19156 15972
rect 19208 15960 19214 15972
rect 20806 15960 20812 15972
rect 19208 15932 20812 15960
rect 19208 15920 19214 15932
rect 20806 15920 20812 15932
rect 20864 15920 20870 15972
rect 13998 15892 14004 15904
rect 13280 15864 14004 15892
rect 13998 15852 14004 15864
rect 14056 15852 14062 15904
rect 17310 15852 17316 15904
rect 17368 15852 17374 15904
rect 17678 15852 17684 15904
rect 17736 15892 17742 15904
rect 17865 15895 17923 15901
rect 17865 15892 17877 15895
rect 17736 15864 17877 15892
rect 17736 15852 17742 15864
rect 17865 15861 17877 15864
rect 17911 15861 17923 15895
rect 17865 15855 17923 15861
rect 18509 15895 18567 15901
rect 18509 15861 18521 15895
rect 18555 15892 18567 15895
rect 18598 15892 18604 15904
rect 18555 15864 18604 15892
rect 18555 15861 18567 15864
rect 18509 15855 18567 15861
rect 18598 15852 18604 15864
rect 18656 15852 18662 15904
rect 20717 15895 20775 15901
rect 20717 15861 20729 15895
rect 20763 15892 20775 15895
rect 21450 15892 21456 15904
rect 20763 15864 21456 15892
rect 20763 15861 20775 15864
rect 20717 15855 20775 15861
rect 21450 15852 21456 15864
rect 21508 15852 21514 15904
rect 22020 15892 22048 16059
rect 23566 16056 23572 16108
rect 23624 16096 23630 16108
rect 24765 16099 24823 16105
rect 24765 16096 24777 16099
rect 23624 16068 24777 16096
rect 23624 16056 23630 16068
rect 24765 16065 24777 16068
rect 24811 16065 24823 16099
rect 24765 16059 24823 16065
rect 22281 16031 22339 16037
rect 22281 15997 22293 16031
rect 22327 16028 22339 16031
rect 22370 16028 22376 16040
rect 22327 16000 22376 16028
rect 22327 15997 22339 16000
rect 22281 15991 22339 15997
rect 22370 15988 22376 16000
rect 22428 15988 22434 16040
rect 24489 16031 24547 16037
rect 24489 15997 24501 16031
rect 24535 16028 24547 16031
rect 24578 16028 24584 16040
rect 24535 16000 24584 16028
rect 24535 15997 24547 16000
rect 24489 15991 24547 15997
rect 24578 15988 24584 16000
rect 24636 15988 24642 16040
rect 22278 15892 22284 15904
rect 22020 15864 22284 15892
rect 22278 15852 22284 15864
rect 22336 15892 22342 15904
rect 23382 15892 23388 15904
rect 22336 15864 23388 15892
rect 22336 15852 22342 15864
rect 23382 15852 23388 15864
rect 23440 15852 23446 15904
rect 23750 15852 23756 15904
rect 23808 15852 23814 15904
rect 24121 15895 24179 15901
rect 24121 15861 24133 15895
rect 24167 15892 24179 15895
rect 24210 15892 24216 15904
rect 24167 15864 24216 15892
rect 24167 15861 24179 15864
rect 24121 15855 24179 15861
rect 24210 15852 24216 15864
rect 24268 15852 24274 15904
rect 1104 15802 25852 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 25852 15802
rect 1104 15728 25852 15750
rect 9030 15648 9036 15700
rect 9088 15688 9094 15700
rect 9125 15691 9183 15697
rect 9125 15688 9137 15691
rect 9088 15660 9137 15688
rect 9088 15648 9094 15660
rect 9125 15657 9137 15660
rect 9171 15657 9183 15691
rect 9125 15651 9183 15657
rect 11146 15648 11152 15700
rect 11204 15688 11210 15700
rect 11609 15691 11667 15697
rect 11609 15688 11621 15691
rect 11204 15660 11621 15688
rect 11204 15648 11210 15660
rect 11609 15657 11621 15660
rect 11655 15657 11667 15691
rect 11609 15651 11667 15657
rect 15010 15648 15016 15700
rect 15068 15688 15074 15700
rect 15473 15691 15531 15697
rect 15473 15688 15485 15691
rect 15068 15660 15485 15688
rect 15068 15648 15074 15660
rect 15473 15657 15485 15660
rect 15519 15688 15531 15691
rect 17126 15688 17132 15700
rect 15519 15660 17132 15688
rect 15519 15657 15531 15660
rect 15473 15651 15531 15657
rect 17126 15648 17132 15660
rect 17184 15688 17190 15700
rect 18230 15688 18236 15700
rect 17184 15660 18236 15688
rect 17184 15648 17190 15660
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 18509 15691 18567 15697
rect 18509 15657 18521 15691
rect 18555 15688 18567 15691
rect 19150 15688 19156 15700
rect 18555 15660 19156 15688
rect 18555 15657 18567 15660
rect 18509 15651 18567 15657
rect 5442 15580 5448 15632
rect 5500 15620 5506 15632
rect 12710 15620 12716 15632
rect 5500 15592 12716 15620
rect 5500 15580 5506 15592
rect 12710 15580 12716 15592
rect 12768 15620 12774 15632
rect 13173 15623 13231 15629
rect 13173 15620 13185 15623
rect 12768 15592 13185 15620
rect 12768 15580 12774 15592
rect 13173 15589 13185 15592
rect 13219 15589 13231 15623
rect 13173 15583 13231 15589
rect 9582 15512 9588 15564
rect 9640 15552 9646 15564
rect 9677 15555 9735 15561
rect 9677 15552 9689 15555
rect 9640 15524 9689 15552
rect 9640 15512 9646 15524
rect 9677 15521 9689 15524
rect 9723 15521 9735 15555
rect 9677 15515 9735 15521
rect 12250 15512 12256 15564
rect 12308 15552 12314 15564
rect 12621 15555 12679 15561
rect 12621 15552 12633 15555
rect 12308 15524 12633 15552
rect 12308 15512 12314 15524
rect 12621 15521 12633 15524
rect 12667 15521 12679 15555
rect 12621 15515 12679 15521
rect 16390 15512 16396 15564
rect 16448 15512 16454 15564
rect 16669 15555 16727 15561
rect 16669 15521 16681 15555
rect 16715 15552 16727 15555
rect 18322 15552 18328 15564
rect 16715 15524 18328 15552
rect 16715 15521 16727 15524
rect 16669 15515 16727 15521
rect 18322 15512 18328 15524
rect 18380 15512 18386 15564
rect 8662 15444 8668 15496
rect 8720 15484 8726 15496
rect 10137 15487 10195 15493
rect 10137 15484 10149 15487
rect 8720 15456 10149 15484
rect 8720 15444 8726 15456
rect 10137 15453 10149 15456
rect 10183 15453 10195 15487
rect 10137 15447 10195 15453
rect 12069 15487 12127 15493
rect 12069 15453 12081 15487
rect 12115 15484 12127 15487
rect 13354 15484 13360 15496
rect 12115 15456 13360 15484
rect 12115 15453 12127 15456
rect 12069 15447 12127 15453
rect 13354 15444 13360 15456
rect 13412 15444 13418 15496
rect 18524 15484 18552 15651
rect 19150 15648 19156 15660
rect 19208 15648 19214 15700
rect 20438 15648 20444 15700
rect 20496 15688 20502 15700
rect 21177 15691 21235 15697
rect 21177 15688 21189 15691
rect 20496 15660 21189 15688
rect 20496 15648 20502 15660
rect 21177 15657 21189 15660
rect 21223 15657 21235 15691
rect 21177 15651 21235 15657
rect 23014 15648 23020 15700
rect 23072 15688 23078 15700
rect 23072 15660 23888 15688
rect 23072 15648 23078 15660
rect 21358 15580 21364 15632
rect 21416 15620 21422 15632
rect 21416 15592 22416 15620
rect 21416 15580 21422 15592
rect 19429 15555 19487 15561
rect 19429 15521 19441 15555
rect 19475 15552 19487 15555
rect 20254 15552 20260 15564
rect 19475 15524 20260 15552
rect 19475 15521 19487 15524
rect 19429 15515 19487 15521
rect 20254 15512 20260 15524
rect 20312 15512 20318 15564
rect 22278 15512 22284 15564
rect 22336 15512 22342 15564
rect 22388 15552 22416 15592
rect 22557 15555 22615 15561
rect 22557 15552 22569 15555
rect 22388 15524 22569 15552
rect 22557 15521 22569 15524
rect 22603 15552 22615 15555
rect 23750 15552 23756 15564
rect 22603 15524 23756 15552
rect 22603 15521 22615 15524
rect 22557 15515 22615 15521
rect 23750 15512 23756 15524
rect 23808 15512 23814 15564
rect 17802 15456 18552 15484
rect 20806 15444 20812 15496
rect 20864 15484 20870 15496
rect 20864 15456 21036 15484
rect 20864 15444 20870 15456
rect 9214 15376 9220 15428
rect 9272 15416 9278 15428
rect 9585 15419 9643 15425
rect 9585 15416 9597 15419
rect 9272 15388 9597 15416
rect 9272 15376 9278 15388
rect 9585 15385 9597 15388
rect 9631 15385 9643 15419
rect 9585 15379 9643 15385
rect 11977 15419 12035 15425
rect 11977 15385 11989 15419
rect 12023 15416 12035 15419
rect 12526 15416 12532 15428
rect 12023 15388 12532 15416
rect 12023 15385 12035 15388
rect 11977 15379 12035 15385
rect 12526 15376 12532 15388
rect 12584 15376 12590 15428
rect 16390 15376 16396 15428
rect 16448 15416 16454 15428
rect 16942 15416 16948 15428
rect 16448 15388 16948 15416
rect 16448 15376 16454 15388
rect 16942 15376 16948 15388
rect 17000 15376 17006 15428
rect 19702 15376 19708 15428
rect 19760 15376 19766 15428
rect 21008 15416 21036 15456
rect 21082 15444 21088 15496
rect 21140 15484 21146 15496
rect 21821 15487 21879 15493
rect 21821 15484 21833 15487
rect 21140 15456 21833 15484
rect 21140 15444 21146 15456
rect 21821 15453 21833 15456
rect 21867 15453 21879 15487
rect 21821 15447 21879 15453
rect 21358 15416 21364 15428
rect 21008 15388 21364 15416
rect 21358 15376 21364 15388
rect 21416 15416 21422 15428
rect 23014 15416 23020 15428
rect 21416 15388 23020 15416
rect 21416 15376 21422 15388
rect 23014 15376 23020 15388
rect 23072 15376 23078 15428
rect 23860 15416 23888 15660
rect 23934 15512 23940 15564
rect 23992 15552 23998 15564
rect 24029 15555 24087 15561
rect 24029 15552 24041 15555
rect 23992 15524 24041 15552
rect 23992 15512 23998 15524
rect 24029 15521 24041 15524
rect 24075 15521 24087 15555
rect 24029 15515 24087 15521
rect 24581 15555 24639 15561
rect 24581 15521 24593 15555
rect 24627 15552 24639 15555
rect 24670 15552 24676 15564
rect 24627 15524 24676 15552
rect 24627 15521 24639 15524
rect 24581 15515 24639 15521
rect 24670 15512 24676 15524
rect 24728 15512 24734 15564
rect 23782 15388 24256 15416
rect 24228 15360 24256 15388
rect 9493 15351 9551 15357
rect 9493 15317 9505 15351
rect 9539 15348 9551 15351
rect 10042 15348 10048 15360
rect 9539 15320 10048 15348
rect 9539 15317 9551 15320
rect 9493 15311 9551 15317
rect 10042 15308 10048 15320
rect 10100 15308 10106 15360
rect 12434 15308 12440 15360
rect 12492 15348 12498 15360
rect 14182 15348 14188 15360
rect 12492 15320 14188 15348
rect 12492 15308 12498 15320
rect 14182 15308 14188 15320
rect 14240 15308 14246 15360
rect 14274 15308 14280 15360
rect 14332 15308 14338 15360
rect 14734 15308 14740 15360
rect 14792 15308 14798 15360
rect 15746 15308 15752 15360
rect 15804 15308 15810 15360
rect 16758 15308 16764 15360
rect 16816 15348 16822 15360
rect 17494 15348 17500 15360
rect 16816 15320 17500 15348
rect 16816 15308 16822 15320
rect 17494 15308 17500 15320
rect 17552 15348 17558 15360
rect 18141 15351 18199 15357
rect 18141 15348 18153 15351
rect 17552 15320 18153 15348
rect 17552 15308 17558 15320
rect 18141 15317 18153 15320
rect 18187 15317 18199 15351
rect 18141 15311 18199 15317
rect 19518 15308 19524 15360
rect 19576 15348 19582 15360
rect 20346 15348 20352 15360
rect 19576 15320 20352 15348
rect 19576 15308 19582 15320
rect 20346 15308 20352 15320
rect 20404 15308 20410 15360
rect 21637 15351 21695 15357
rect 21637 15317 21649 15351
rect 21683 15348 21695 15351
rect 23934 15348 23940 15360
rect 21683 15320 23940 15348
rect 21683 15317 21695 15320
rect 21637 15311 21695 15317
rect 23934 15308 23940 15320
rect 23992 15308 23998 15360
rect 24210 15308 24216 15360
rect 24268 15348 24274 15360
rect 25041 15351 25099 15357
rect 25041 15348 25053 15351
rect 24268 15320 25053 15348
rect 24268 15308 24274 15320
rect 25041 15317 25053 15320
rect 25087 15317 25099 15351
rect 25041 15311 25099 15317
rect 1104 15258 25852 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 25852 15258
rect 1104 15184 25852 15206
rect 10134 15104 10140 15156
rect 10192 15104 10198 15156
rect 13725 15147 13783 15153
rect 13725 15113 13737 15147
rect 13771 15113 13783 15147
rect 13725 15107 13783 15113
rect 14093 15147 14151 15153
rect 14093 15113 14105 15147
rect 14139 15144 14151 15147
rect 14274 15144 14280 15156
rect 14139 15116 14280 15144
rect 14139 15113 14151 15116
rect 14093 15107 14151 15113
rect 8662 15036 8668 15088
rect 8720 15036 8726 15088
rect 10505 15079 10563 15085
rect 10505 15045 10517 15079
rect 10551 15076 10563 15079
rect 11422 15076 11428 15088
rect 10551 15048 11428 15076
rect 10551 15045 10563 15048
rect 10505 15039 10563 15045
rect 11422 15036 11428 15048
rect 11480 15036 11486 15088
rect 13740 15076 13768 15107
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 15746 15104 15752 15156
rect 15804 15144 15810 15156
rect 15933 15147 15991 15153
rect 15933 15144 15945 15147
rect 15804 15116 15945 15144
rect 15804 15104 15810 15116
rect 15933 15113 15945 15116
rect 15979 15113 15991 15147
rect 15933 15107 15991 15113
rect 17218 15104 17224 15156
rect 17276 15144 17282 15156
rect 17497 15147 17555 15153
rect 17497 15144 17509 15147
rect 17276 15116 17509 15144
rect 17276 15104 17282 15116
rect 17497 15113 17509 15116
rect 17543 15113 17555 15147
rect 17497 15107 17555 15113
rect 19610 15104 19616 15156
rect 19668 15144 19674 15156
rect 20073 15147 20131 15153
rect 20073 15144 20085 15147
rect 19668 15116 20085 15144
rect 19668 15104 19674 15116
rect 20073 15113 20085 15116
rect 20119 15113 20131 15147
rect 20073 15107 20131 15113
rect 21082 15104 21088 15156
rect 21140 15144 21146 15156
rect 21910 15144 21916 15156
rect 21140 15116 21916 15144
rect 21140 15104 21146 15116
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 16114 15076 16120 15088
rect 13740 15048 16120 15076
rect 16114 15036 16120 15048
rect 16172 15036 16178 15088
rect 18693 15079 18751 15085
rect 18693 15045 18705 15079
rect 18739 15076 18751 15079
rect 19242 15076 19248 15088
rect 18739 15048 19248 15076
rect 18739 15045 18751 15048
rect 18693 15039 18751 15045
rect 19242 15036 19248 15048
rect 19300 15036 19306 15088
rect 23198 15076 23204 15088
rect 21008 15048 23204 15076
rect 9582 14968 9588 15020
rect 9640 15008 9646 15020
rect 15930 15008 15936 15020
rect 9640 14980 10732 15008
rect 9640 14968 9646 14980
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14940 7711 14943
rect 7929 14943 7987 14949
rect 7699 14912 7788 14940
rect 7699 14909 7711 14912
rect 7653 14903 7711 14909
rect 7760 14804 7788 14912
rect 7929 14909 7941 14943
rect 7975 14940 7987 14943
rect 8294 14940 8300 14952
rect 7975 14912 8300 14940
rect 7975 14909 7987 14912
rect 7929 14903 7987 14909
rect 8294 14900 8300 14912
rect 8352 14900 8358 14952
rect 10704 14949 10732 14980
rect 14384 14980 15936 15008
rect 9677 14943 9735 14949
rect 9677 14909 9689 14943
rect 9723 14909 9735 14943
rect 9677 14903 9735 14909
rect 10597 14943 10655 14949
rect 10597 14909 10609 14943
rect 10643 14909 10655 14943
rect 10597 14903 10655 14909
rect 10689 14943 10747 14949
rect 10689 14909 10701 14943
rect 10735 14909 10747 14943
rect 10689 14903 10747 14909
rect 9030 14832 9036 14884
rect 9088 14872 9094 14884
rect 9692 14872 9720 14903
rect 9088 14844 9720 14872
rect 10612 14872 10640 14903
rect 11238 14900 11244 14952
rect 11296 14940 11302 14952
rect 14384 14949 14412 14980
rect 15930 14968 15936 14980
rect 15988 14968 15994 15020
rect 19978 14968 19984 15020
rect 20036 14968 20042 15020
rect 21008 15017 21036 15048
rect 23198 15036 23204 15048
rect 23256 15036 23262 15088
rect 23290 15036 23296 15088
rect 23348 15036 23354 15088
rect 25130 15036 25136 15088
rect 25188 15036 25194 15088
rect 20993 15011 21051 15017
rect 20993 14977 21005 15011
rect 21039 14977 21051 15011
rect 20993 14971 21051 14977
rect 21358 14968 21364 15020
rect 21416 14968 21422 15020
rect 22002 14968 22008 15020
rect 22060 15008 22066 15020
rect 22097 15011 22155 15017
rect 22097 15008 22109 15011
rect 22060 14980 22109 15008
rect 22060 14968 22066 14980
rect 22097 14977 22109 14980
rect 22143 14977 22155 15011
rect 22097 14971 22155 14977
rect 24118 14968 24124 15020
rect 24176 14968 24182 15020
rect 13449 14943 13507 14949
rect 13449 14940 13461 14943
rect 11296 14912 13461 14940
rect 11296 14900 11302 14912
rect 13449 14909 13461 14912
rect 13495 14940 13507 14943
rect 14185 14943 14243 14949
rect 14185 14940 14197 14943
rect 13495 14912 14197 14940
rect 13495 14909 13507 14912
rect 13449 14903 13507 14909
rect 14185 14909 14197 14912
rect 14231 14909 14243 14943
rect 14185 14903 14243 14909
rect 14369 14943 14427 14949
rect 14369 14909 14381 14943
rect 14415 14909 14427 14943
rect 16025 14943 16083 14949
rect 16025 14940 16037 14943
rect 14369 14903 14427 14909
rect 15488 14912 16037 14940
rect 11606 14872 11612 14884
rect 10612 14844 11612 14872
rect 9088 14832 9094 14844
rect 11606 14832 11612 14844
rect 11664 14832 11670 14884
rect 11974 14832 11980 14884
rect 12032 14872 12038 14884
rect 12161 14875 12219 14881
rect 12161 14872 12173 14875
rect 12032 14844 12173 14872
rect 12032 14832 12038 14844
rect 12161 14841 12173 14844
rect 12207 14872 12219 14875
rect 13630 14872 13636 14884
rect 12207 14844 13636 14872
rect 12207 14841 12219 14844
rect 12161 14835 12219 14841
rect 13630 14832 13636 14844
rect 13688 14832 13694 14884
rect 15488 14816 15516 14912
rect 16025 14909 16037 14912
rect 16071 14909 16083 14943
rect 16025 14903 16083 14909
rect 16209 14943 16267 14949
rect 16209 14909 16221 14943
rect 16255 14940 16267 14943
rect 16574 14940 16580 14952
rect 16255 14912 16580 14940
rect 16255 14909 16267 14912
rect 16209 14903 16267 14909
rect 16574 14900 16580 14912
rect 16632 14900 16638 14952
rect 19886 14940 19892 14952
rect 17696 14912 19892 14940
rect 15565 14875 15623 14881
rect 15565 14841 15577 14875
rect 15611 14872 15623 14875
rect 17696 14872 17724 14912
rect 19886 14900 19892 14912
rect 19944 14900 19950 14952
rect 20257 14943 20315 14949
rect 20257 14909 20269 14943
rect 20303 14940 20315 14943
rect 20438 14940 20444 14952
rect 20303 14912 20444 14940
rect 20303 14909 20315 14912
rect 20257 14903 20315 14909
rect 20438 14900 20444 14912
rect 20496 14900 20502 14952
rect 22738 14940 22744 14952
rect 20732 14912 22744 14940
rect 15611 14844 17724 14872
rect 19613 14875 19671 14881
rect 15611 14841 15623 14844
rect 15565 14835 15623 14841
rect 19613 14841 19625 14875
rect 19659 14872 19671 14875
rect 20732 14872 20760 14912
rect 22738 14900 22744 14912
rect 22796 14900 22802 14952
rect 19659 14844 20760 14872
rect 20809 14875 20867 14881
rect 19659 14841 19671 14844
rect 19613 14835 19671 14841
rect 20809 14841 20821 14875
rect 20855 14872 20867 14875
rect 20855 14844 21496 14872
rect 20855 14841 20867 14844
rect 20809 14835 20867 14841
rect 8294 14804 8300 14816
rect 7760 14776 8300 14804
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 11333 14807 11391 14813
rect 11333 14773 11345 14807
rect 11379 14804 11391 14807
rect 11514 14804 11520 14816
rect 11379 14776 11520 14804
rect 11379 14773 11391 14776
rect 11333 14767 11391 14773
rect 11514 14764 11520 14776
rect 11572 14804 11578 14816
rect 12342 14804 12348 14816
rect 11572 14776 12348 14804
rect 11572 14764 11578 14776
rect 12342 14764 12348 14776
rect 12400 14764 12406 14816
rect 12529 14807 12587 14813
rect 12529 14773 12541 14807
rect 12575 14804 12587 14807
rect 12802 14804 12808 14816
rect 12575 14776 12808 14804
rect 12575 14773 12587 14776
rect 12529 14767 12587 14773
rect 12802 14764 12808 14776
rect 12860 14764 12866 14816
rect 15289 14807 15347 14813
rect 15289 14773 15301 14807
rect 15335 14804 15347 14807
rect 15470 14804 15476 14816
rect 15335 14776 15476 14804
rect 15335 14773 15347 14776
rect 15289 14767 15347 14773
rect 15470 14764 15476 14776
rect 15528 14764 15534 14816
rect 15838 14764 15844 14816
rect 15896 14804 15902 14816
rect 18785 14807 18843 14813
rect 18785 14804 18797 14807
rect 15896 14776 18797 14804
rect 15896 14764 15902 14776
rect 18785 14773 18797 14776
rect 18831 14773 18843 14807
rect 21468 14804 21496 14844
rect 22278 14804 22284 14816
rect 21468 14776 22284 14804
rect 18785 14767 18843 14773
rect 22278 14764 22284 14776
rect 22336 14764 22342 14816
rect 1104 14714 25852 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 25852 14714
rect 1104 14640 25852 14662
rect 7834 14560 7840 14612
rect 7892 14600 7898 14612
rect 8205 14603 8263 14609
rect 8205 14600 8217 14603
rect 7892 14572 8217 14600
rect 7892 14560 7898 14572
rect 8205 14569 8217 14572
rect 8251 14569 8263 14603
rect 8205 14563 8263 14569
rect 8573 14603 8631 14609
rect 8573 14569 8585 14603
rect 8619 14600 8631 14603
rect 8662 14600 8668 14612
rect 8619 14572 8668 14600
rect 8619 14569 8631 14572
rect 8573 14563 8631 14569
rect 8588 14532 8616 14563
rect 8662 14560 8668 14572
rect 8720 14560 8726 14612
rect 9030 14560 9036 14612
rect 9088 14600 9094 14612
rect 12437 14603 12495 14609
rect 9088 14572 11284 14600
rect 9088 14560 9094 14572
rect 9585 14535 9643 14541
rect 9585 14532 9597 14535
rect 8588 14504 9597 14532
rect 6454 14424 6460 14476
rect 6512 14464 6518 14476
rect 8294 14464 8300 14476
rect 6512 14436 8300 14464
rect 6512 14424 6518 14436
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 8588 14396 8616 14504
rect 7866 14368 8616 14396
rect 6733 14331 6791 14337
rect 6733 14297 6745 14331
rect 6779 14297 6791 14331
rect 9306 14328 9312 14340
rect 6733 14291 6791 14297
rect 8404 14300 9312 14328
rect 6748 14260 6776 14291
rect 8404 14260 8432 14300
rect 9306 14288 9312 14300
rect 9364 14288 9370 14340
rect 9508 14328 9536 14504
rect 9585 14501 9597 14504
rect 9631 14501 9643 14535
rect 11256 14532 11284 14572
rect 12437 14569 12449 14603
rect 12483 14600 12495 14603
rect 12618 14600 12624 14612
rect 12483 14572 12624 14600
rect 12483 14569 12495 14572
rect 12437 14563 12495 14569
rect 12618 14560 12624 14572
rect 12676 14560 12682 14612
rect 14642 14560 14648 14612
rect 14700 14600 14706 14612
rect 15381 14603 15439 14609
rect 15381 14600 15393 14603
rect 14700 14572 15393 14600
rect 14700 14560 14706 14572
rect 15381 14569 15393 14572
rect 15427 14600 15439 14603
rect 20162 14600 20168 14612
rect 15427 14572 20168 14600
rect 15427 14569 15439 14572
rect 15381 14563 15439 14569
rect 20162 14560 20168 14572
rect 20220 14560 20226 14612
rect 21453 14603 21511 14609
rect 21453 14569 21465 14603
rect 21499 14600 21511 14603
rect 24026 14600 24032 14612
rect 21499 14572 24032 14600
rect 21499 14569 21511 14572
rect 21453 14563 21511 14569
rect 24026 14560 24032 14572
rect 24084 14560 24090 14612
rect 11256 14504 14964 14532
rect 9585 14495 9643 14501
rect 10226 14424 10232 14476
rect 10284 14424 10290 14476
rect 11882 14424 11888 14476
rect 11940 14464 11946 14476
rect 11977 14467 12035 14473
rect 11977 14464 11989 14467
rect 11940 14436 11989 14464
rect 11940 14424 11946 14436
rect 11977 14433 11989 14436
rect 12023 14464 12035 14467
rect 12250 14464 12256 14476
rect 12023 14436 12256 14464
rect 12023 14433 12035 14436
rect 11977 14427 12035 14433
rect 12250 14424 12256 14436
rect 12308 14464 12314 14476
rect 14936 14473 14964 14504
rect 16850 14492 16856 14544
rect 16908 14532 16914 14544
rect 16908 14504 16988 14532
rect 16908 14492 16914 14504
rect 12989 14467 13047 14473
rect 12989 14464 13001 14467
rect 12308 14436 13001 14464
rect 12308 14424 12314 14436
rect 12989 14433 13001 14436
rect 13035 14433 13047 14467
rect 12989 14427 13047 14433
rect 14921 14467 14979 14473
rect 14921 14433 14933 14467
rect 14967 14464 14979 14467
rect 15378 14464 15384 14476
rect 14967 14436 15384 14464
rect 14967 14433 14979 14436
rect 14921 14427 14979 14433
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 16960 14473 16988 14504
rect 19518 14492 19524 14544
rect 19576 14532 19582 14544
rect 22462 14532 22468 14544
rect 19576 14504 22468 14532
rect 19576 14492 19582 14504
rect 22462 14492 22468 14504
rect 22520 14492 22526 14544
rect 16945 14467 17003 14473
rect 16945 14433 16957 14467
rect 16991 14433 17003 14467
rect 16945 14427 17003 14433
rect 17126 14424 17132 14476
rect 17184 14424 17190 14476
rect 20622 14424 20628 14476
rect 20680 14464 20686 14476
rect 21913 14467 21971 14473
rect 21913 14464 21925 14467
rect 20680 14436 21925 14464
rect 20680 14424 20686 14436
rect 21913 14433 21925 14436
rect 21959 14433 21971 14467
rect 21913 14427 21971 14433
rect 22097 14467 22155 14473
rect 22097 14433 22109 14467
rect 22143 14464 22155 14467
rect 23290 14464 23296 14476
rect 22143 14436 23296 14464
rect 22143 14433 22155 14436
rect 22097 14427 22155 14433
rect 23290 14424 23296 14436
rect 23348 14424 23354 14476
rect 23845 14467 23903 14473
rect 23845 14433 23857 14467
rect 23891 14464 23903 14467
rect 24854 14464 24860 14476
rect 23891 14436 24860 14464
rect 23891 14433 23903 14436
rect 23845 14427 23903 14433
rect 24854 14424 24860 14436
rect 24912 14424 24918 14476
rect 9582 14356 9588 14408
rect 9640 14396 9646 14408
rect 9953 14399 10011 14405
rect 9953 14396 9965 14399
rect 9640 14368 9965 14396
rect 9640 14356 9646 14368
rect 9953 14365 9965 14368
rect 9999 14365 10011 14399
rect 9953 14359 10011 14365
rect 13078 14356 13084 14408
rect 13136 14396 13142 14408
rect 13449 14399 13507 14405
rect 13449 14396 13461 14399
rect 13136 14368 13461 14396
rect 13136 14356 13142 14368
rect 13449 14365 13461 14368
rect 13495 14396 13507 14399
rect 13495 14368 14872 14396
rect 13495 14365 13507 14368
rect 13449 14359 13507 14365
rect 12897 14331 12955 14337
rect 9508 14300 10718 14328
rect 12897 14297 12909 14331
rect 12943 14328 12955 14331
rect 13630 14328 13636 14340
rect 12943 14300 13636 14328
rect 12943 14297 12955 14300
rect 12897 14291 12955 14297
rect 13630 14288 13636 14300
rect 13688 14288 13694 14340
rect 14734 14328 14740 14340
rect 13924 14300 14740 14328
rect 13924 14272 13952 14300
rect 14734 14288 14740 14300
rect 14792 14288 14798 14340
rect 14844 14328 14872 14368
rect 16114 14356 16120 14408
rect 16172 14396 16178 14408
rect 19610 14396 19616 14408
rect 16172 14368 19616 14396
rect 16172 14356 16178 14368
rect 19610 14356 19616 14368
rect 19668 14356 19674 14408
rect 20441 14399 20499 14405
rect 20441 14365 20453 14399
rect 20487 14396 20499 14399
rect 21634 14396 21640 14408
rect 20487 14368 21640 14396
rect 20487 14365 20499 14368
rect 20441 14359 20499 14365
rect 21634 14356 21640 14368
rect 21692 14356 21698 14408
rect 22833 14399 22891 14405
rect 22833 14365 22845 14399
rect 22879 14396 22891 14399
rect 24486 14396 24492 14408
rect 22879 14368 24492 14396
rect 22879 14365 22891 14368
rect 22833 14359 22891 14365
rect 24486 14356 24492 14368
rect 24544 14356 24550 14408
rect 25038 14356 25044 14408
rect 25096 14356 25102 14408
rect 16853 14331 16911 14337
rect 14844 14300 16620 14328
rect 6748 14232 8432 14260
rect 12710 14220 12716 14272
rect 12768 14260 12774 14272
rect 12805 14263 12863 14269
rect 12805 14260 12817 14263
rect 12768 14232 12817 14260
rect 12768 14220 12774 14232
rect 12805 14229 12817 14232
rect 12851 14229 12863 14263
rect 12805 14223 12863 14229
rect 13906 14220 13912 14272
rect 13964 14220 13970 14272
rect 14274 14220 14280 14272
rect 14332 14220 14338 14272
rect 14642 14220 14648 14272
rect 14700 14220 14706 14272
rect 16482 14220 16488 14272
rect 16540 14220 16546 14272
rect 16592 14260 16620 14300
rect 16853 14297 16865 14331
rect 16899 14328 16911 14331
rect 17681 14331 17739 14337
rect 17681 14328 17693 14331
rect 16899 14300 17693 14328
rect 16899 14297 16911 14300
rect 16853 14291 16911 14297
rect 17681 14297 17693 14300
rect 17727 14297 17739 14331
rect 21266 14328 21272 14340
rect 17681 14291 17739 14297
rect 19306 14300 21272 14328
rect 19306 14272 19334 14300
rect 21266 14288 21272 14300
rect 21324 14288 21330 14340
rect 19306 14260 19340 14272
rect 16592 14232 19340 14260
rect 19334 14220 19340 14232
rect 19392 14220 19398 14272
rect 19886 14220 19892 14272
rect 19944 14260 19950 14272
rect 20257 14263 20315 14269
rect 20257 14260 20269 14263
rect 19944 14232 20269 14260
rect 19944 14220 19950 14232
rect 20257 14229 20269 14232
rect 20303 14229 20315 14263
rect 20257 14223 20315 14229
rect 21818 14220 21824 14272
rect 21876 14220 21882 14272
rect 24854 14220 24860 14272
rect 24912 14220 24918 14272
rect 1104 14170 25852 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 25852 14170
rect 1104 14096 25852 14118
rect 8294 14056 8300 14068
rect 7852 14028 8300 14056
rect 7852 13988 7880 14028
rect 8294 14016 8300 14028
rect 8352 14056 8358 14068
rect 9582 14056 9588 14068
rect 8352 14028 9588 14056
rect 8352 14016 8358 14028
rect 9582 14016 9588 14028
rect 9640 14016 9646 14068
rect 12250 14016 12256 14068
rect 12308 14016 12314 14068
rect 12989 14059 13047 14065
rect 12989 14025 13001 14059
rect 13035 14056 13047 14059
rect 13078 14056 13084 14068
rect 13035 14028 13084 14056
rect 13035 14025 13047 14028
rect 12989 14019 13047 14025
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 15562 14016 15568 14068
rect 15620 14016 15626 14068
rect 16482 14016 16488 14068
rect 16540 14056 16546 14068
rect 23382 14056 23388 14068
rect 16540 14028 20392 14056
rect 16540 14016 16546 14028
rect 7760 13960 7880 13988
rect 7760 13929 7788 13960
rect 7926 13948 7932 14000
rect 7984 13988 7990 14000
rect 8021 13991 8079 13997
rect 8021 13988 8033 13991
rect 7984 13960 8033 13988
rect 7984 13948 7990 13960
rect 8021 13957 8033 13960
rect 8067 13957 8079 13991
rect 8021 13951 8079 13957
rect 8662 13948 8668 14000
rect 8720 13948 8726 14000
rect 10229 13991 10287 13997
rect 10229 13957 10241 13991
rect 10275 13988 10287 13991
rect 12342 13988 12348 14000
rect 10275 13960 12348 13988
rect 10275 13957 10287 13960
rect 10229 13951 10287 13957
rect 12342 13948 12348 13960
rect 12400 13948 12406 14000
rect 15580 13988 15608 14016
rect 17126 13988 17132 14000
rect 15580 13960 17132 13988
rect 17126 13948 17132 13960
rect 17184 13948 17190 14000
rect 19150 13988 19156 14000
rect 18354 13960 19156 13988
rect 19150 13948 19156 13960
rect 19208 13948 19214 14000
rect 19518 13948 19524 14000
rect 19576 13948 19582 14000
rect 19610 13948 19616 14000
rect 19668 13988 19674 14000
rect 19705 13991 19763 13997
rect 19705 13988 19717 13991
rect 19668 13960 19717 13988
rect 19668 13948 19674 13960
rect 19705 13957 19717 13960
rect 19751 13957 19763 13991
rect 19705 13951 19763 13957
rect 7745 13923 7803 13929
rect 7745 13889 7757 13923
rect 7791 13889 7803 13923
rect 7745 13883 7803 13889
rect 9582 13880 9588 13932
rect 9640 13920 9646 13932
rect 20364 13929 20392 14028
rect 21192 14028 23388 14056
rect 10965 13923 11023 13929
rect 10965 13920 10977 13923
rect 9640 13892 10977 13920
rect 9640 13880 9646 13892
rect 10965 13889 10977 13892
rect 11011 13889 11023 13923
rect 18969 13923 19027 13929
rect 18969 13920 18981 13923
rect 10965 13883 11023 13889
rect 9769 13855 9827 13861
rect 9769 13821 9781 13855
rect 9815 13852 9827 13855
rect 10226 13852 10232 13864
rect 9815 13824 10232 13852
rect 9815 13821 9827 13824
rect 9769 13815 9827 13821
rect 10226 13812 10232 13824
rect 10284 13812 10290 13864
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 11112 13824 11713 13852
rect 11112 13812 11118 13824
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 11701 13815 11759 13821
rect 12250 13812 12256 13864
rect 12308 13852 12314 13864
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 12308 13824 13093 13852
rect 12308 13812 12314 13824
rect 13081 13821 13093 13824
rect 13127 13821 13139 13855
rect 13081 13815 13139 13821
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13821 13231 13855
rect 13173 13815 13231 13821
rect 12802 13744 12808 13796
rect 12860 13784 12866 13796
rect 13188 13784 13216 13815
rect 13814 13812 13820 13864
rect 13872 13812 13878 13864
rect 15212 13852 15240 13906
rect 18340 13892 18981 13920
rect 15933 13855 15991 13861
rect 15933 13852 15945 13855
rect 13924 13824 15148 13852
rect 15212 13824 15945 13852
rect 13924 13784 13952 13824
rect 12860 13756 13952 13784
rect 15120 13784 15148 13824
rect 15933 13821 15945 13824
rect 15979 13852 15991 13855
rect 16482 13852 16488 13864
rect 15979 13824 16488 13852
rect 15979 13821 15991 13824
rect 15933 13815 15991 13821
rect 16482 13812 16488 13824
rect 16540 13812 16546 13864
rect 16850 13812 16856 13864
rect 16908 13812 16914 13864
rect 17129 13855 17187 13861
rect 17129 13821 17141 13855
rect 17175 13852 17187 13855
rect 17586 13852 17592 13864
rect 17175 13824 17592 13852
rect 17175 13821 17187 13824
rect 17129 13815 17187 13821
rect 17586 13812 17592 13824
rect 17644 13852 17650 13864
rect 17862 13852 17868 13864
rect 17644 13824 17868 13852
rect 17644 13812 17650 13824
rect 17862 13812 17868 13824
rect 17920 13852 17926 13864
rect 18340 13852 18368 13892
rect 18969 13889 18981 13892
rect 19015 13889 19027 13923
rect 18969 13883 19027 13889
rect 20349 13923 20407 13929
rect 20349 13889 20361 13923
rect 20395 13889 20407 13923
rect 20349 13883 20407 13889
rect 21082 13880 21088 13932
rect 21140 13880 21146 13932
rect 17920 13824 18368 13852
rect 18601 13855 18659 13861
rect 17920 13812 17926 13824
rect 18601 13821 18613 13855
rect 18647 13852 18659 13855
rect 18874 13852 18880 13864
rect 18647 13824 18880 13852
rect 18647 13821 18659 13824
rect 18601 13815 18659 13821
rect 18874 13812 18880 13824
rect 18932 13812 18938 13864
rect 21192 13852 21220 14028
rect 23382 14016 23388 14028
rect 23440 14016 23446 14068
rect 23492 14028 25268 14056
rect 21542 13948 21548 14000
rect 21600 13988 21606 14000
rect 23492 13988 23520 14028
rect 21600 13960 23520 13988
rect 21600 13948 21606 13960
rect 21266 13880 21272 13932
rect 21324 13920 21330 13932
rect 22189 13923 22247 13929
rect 22189 13920 22201 13923
rect 21324 13892 22201 13920
rect 21324 13880 21330 13892
rect 22189 13889 22201 13892
rect 22235 13889 22247 13923
rect 22189 13883 22247 13889
rect 24210 13880 24216 13932
rect 24268 13880 24274 13932
rect 25240 13929 25268 14028
rect 25225 13923 25283 13929
rect 25225 13889 25237 13923
rect 25271 13889 25283 13923
rect 25225 13883 25283 13889
rect 22646 13852 22652 13864
rect 20180 13824 21220 13852
rect 22020 13824 22652 13852
rect 15562 13784 15568 13796
rect 15120 13756 15568 13784
rect 12860 13744 12866 13756
rect 15562 13744 15568 13756
rect 15620 13744 15626 13796
rect 20180 13793 20208 13824
rect 22020 13793 22048 13824
rect 22646 13812 22652 13824
rect 22704 13812 22710 13864
rect 22830 13812 22836 13864
rect 22888 13812 22894 13864
rect 23109 13855 23167 13861
rect 23109 13852 23121 13855
rect 22940 13824 23121 13852
rect 20165 13787 20223 13793
rect 20165 13753 20177 13787
rect 20211 13753 20223 13787
rect 20165 13747 20223 13753
rect 22005 13787 22063 13793
rect 22005 13753 22017 13787
rect 22051 13753 22063 13787
rect 22005 13747 22063 13753
rect 12618 13676 12624 13728
rect 12676 13676 12682 13728
rect 14090 13725 14096 13728
rect 14080 13719 14096 13725
rect 14080 13685 14092 13719
rect 14080 13679 14096 13685
rect 14090 13676 14096 13679
rect 14148 13676 14154 13728
rect 18322 13676 18328 13728
rect 18380 13716 18386 13728
rect 20622 13716 20628 13728
rect 18380 13688 20628 13716
rect 18380 13676 18386 13688
rect 20622 13676 20628 13688
rect 20680 13676 20686 13728
rect 20898 13676 20904 13728
rect 20956 13676 20962 13728
rect 20990 13676 20996 13728
rect 21048 13716 21054 13728
rect 22940 13716 22968 13824
rect 23109 13821 23121 13824
rect 23155 13821 23167 13855
rect 23109 13815 23167 13821
rect 23198 13812 23204 13864
rect 23256 13852 23262 13864
rect 24581 13855 24639 13861
rect 24581 13852 24593 13855
rect 23256 13824 24593 13852
rect 23256 13812 23262 13824
rect 24581 13821 24593 13824
rect 24627 13821 24639 13855
rect 24581 13815 24639 13821
rect 23842 13716 23848 13728
rect 21048 13688 23848 13716
rect 21048 13676 21054 13688
rect 23842 13676 23848 13688
rect 23900 13676 23906 13728
rect 25038 13676 25044 13728
rect 25096 13676 25102 13728
rect 1104 13626 25852 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 25852 13626
rect 1104 13552 25852 13574
rect 8297 13515 8355 13521
rect 8297 13481 8309 13515
rect 8343 13512 8355 13515
rect 8386 13512 8392 13524
rect 8343 13484 8392 13512
rect 8343 13481 8355 13484
rect 8297 13475 8355 13481
rect 8386 13472 8392 13484
rect 8444 13472 8450 13524
rect 8662 13472 8668 13524
rect 8720 13472 8726 13524
rect 8846 13472 8852 13524
rect 8904 13512 8910 13524
rect 9217 13515 9275 13521
rect 9217 13512 9229 13515
rect 8904 13484 9229 13512
rect 8904 13472 8910 13484
rect 9217 13481 9229 13484
rect 9263 13481 9275 13515
rect 9217 13475 9275 13481
rect 10676 13515 10734 13521
rect 10676 13481 10688 13515
rect 10722 13512 10734 13515
rect 13538 13512 13544 13524
rect 10722 13484 13544 13512
rect 10722 13481 10734 13484
rect 10676 13475 10734 13481
rect 13538 13472 13544 13484
rect 13596 13472 13602 13524
rect 14734 13472 14740 13524
rect 14792 13512 14798 13524
rect 21082 13512 21088 13524
rect 14792 13484 21088 13512
rect 14792 13472 14798 13484
rect 21082 13472 21088 13484
rect 21140 13472 21146 13524
rect 24486 13472 24492 13524
rect 24544 13512 24550 13524
rect 24581 13515 24639 13521
rect 24581 13512 24593 13515
rect 24544 13484 24593 13512
rect 24544 13472 24550 13484
rect 24581 13481 24593 13484
rect 24627 13481 24639 13515
rect 24581 13475 24639 13481
rect 9306 13404 9312 13456
rect 9364 13444 9370 13456
rect 9364 13416 9812 13444
rect 9364 13404 9370 13416
rect 6454 13336 6460 13388
rect 6512 13376 6518 13388
rect 6549 13379 6607 13385
rect 6549 13376 6561 13379
rect 6512 13348 6561 13376
rect 6512 13336 6518 13348
rect 6549 13345 6561 13348
rect 6595 13345 6607 13379
rect 6549 13339 6607 13345
rect 6825 13379 6883 13385
rect 6825 13345 6837 13379
rect 6871 13376 6883 13379
rect 9674 13376 9680 13388
rect 6871 13348 9680 13376
rect 6871 13345 6883 13348
rect 6825 13339 6883 13345
rect 9674 13336 9680 13348
rect 9732 13336 9738 13388
rect 9784 13385 9812 13416
rect 11790 13404 11796 13456
rect 11848 13444 11854 13456
rect 14550 13444 14556 13456
rect 11848 13416 14556 13444
rect 11848 13404 11854 13416
rect 14550 13404 14556 13416
rect 14608 13404 14614 13456
rect 17126 13404 17132 13456
rect 17184 13444 17190 13456
rect 24210 13444 24216 13456
rect 17184 13416 24216 13444
rect 17184 13404 17190 13416
rect 24210 13404 24216 13416
rect 24268 13404 24274 13456
rect 9769 13379 9827 13385
rect 9769 13345 9781 13379
rect 9815 13345 9827 13379
rect 9769 13339 9827 13345
rect 10413 13379 10471 13385
rect 10413 13345 10425 13379
rect 10459 13376 10471 13379
rect 11698 13376 11704 13388
rect 10459 13348 11704 13376
rect 10459 13345 10471 13348
rect 10413 13339 10471 13345
rect 11698 13336 11704 13348
rect 11756 13376 11762 13388
rect 13449 13379 13507 13385
rect 13449 13376 13461 13379
rect 11756 13348 13461 13376
rect 11756 13336 11762 13348
rect 13449 13345 13461 13348
rect 13495 13376 13507 13379
rect 13814 13376 13820 13388
rect 13495 13348 13820 13376
rect 13495 13345 13507 13348
rect 13449 13339 13507 13345
rect 13814 13336 13820 13348
rect 13872 13336 13878 13388
rect 15378 13336 15384 13388
rect 15436 13376 15442 13388
rect 15746 13376 15752 13388
rect 15436 13348 15752 13376
rect 15436 13336 15442 13348
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 16301 13379 16359 13385
rect 16301 13345 16313 13379
rect 16347 13376 16359 13379
rect 20070 13376 20076 13388
rect 16347 13348 20076 13376
rect 16347 13345 16359 13348
rect 16301 13339 16359 13345
rect 12434 13268 12440 13320
rect 12492 13308 12498 13320
rect 12621 13311 12679 13317
rect 12621 13308 12633 13311
rect 12492 13280 12633 13308
rect 12492 13268 12498 13280
rect 12621 13277 12633 13280
rect 12667 13308 12679 13311
rect 12667 13280 12848 13308
rect 12667 13277 12679 13280
rect 12621 13271 12679 13277
rect 8662 13240 8668 13252
rect 8050 13212 8668 13240
rect 8662 13200 8668 13212
rect 8720 13200 8726 13252
rect 9585 13243 9643 13249
rect 9585 13209 9597 13243
rect 9631 13240 9643 13243
rect 11974 13240 11980 13252
rect 9631 13212 11100 13240
rect 11914 13212 11980 13240
rect 9631 13209 9643 13212
rect 9585 13203 9643 13209
rect 9674 13132 9680 13184
rect 9732 13132 9738 13184
rect 11072 13172 11100 13212
rect 11974 13200 11980 13212
rect 12032 13200 12038 13252
rect 12066 13172 12072 13184
rect 11072 13144 12072 13172
rect 12066 13132 12072 13144
rect 12124 13132 12130 13184
rect 12158 13132 12164 13184
rect 12216 13132 12222 13184
rect 12820 13172 12848 13280
rect 12986 13268 12992 13320
rect 13044 13308 13050 13320
rect 13354 13308 13360 13320
rect 13044 13280 13360 13308
rect 13044 13268 13050 13280
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 14366 13268 14372 13320
rect 14424 13308 14430 13320
rect 14550 13308 14556 13320
rect 14424 13280 14556 13308
rect 14424 13268 14430 13280
rect 14550 13268 14556 13280
rect 14608 13268 14614 13320
rect 14918 13268 14924 13320
rect 14976 13308 14982 13320
rect 15657 13311 15715 13317
rect 15657 13308 15669 13311
rect 14976 13280 15669 13308
rect 14976 13268 14982 13280
rect 15657 13277 15669 13280
rect 15703 13308 15715 13311
rect 16206 13308 16212 13320
rect 15703 13280 16212 13308
rect 15703 13277 15715 13280
rect 15657 13271 15715 13277
rect 16206 13268 16212 13280
rect 16264 13268 16270 13320
rect 15565 13243 15623 13249
rect 15565 13209 15577 13243
rect 15611 13240 15623 13243
rect 16316 13240 16344 13339
rect 20070 13336 20076 13348
rect 20128 13336 20134 13388
rect 20257 13379 20315 13385
rect 20257 13345 20269 13379
rect 20303 13376 20315 13379
rect 20438 13376 20444 13388
rect 20303 13348 20444 13376
rect 20303 13345 20315 13348
rect 20257 13339 20315 13345
rect 20438 13336 20444 13348
rect 20496 13376 20502 13388
rect 22830 13376 22836 13388
rect 20496 13348 22836 13376
rect 20496 13336 20502 13348
rect 22830 13336 22836 13348
rect 22888 13336 22894 13388
rect 23750 13336 23756 13388
rect 23808 13336 23814 13388
rect 25038 13376 25044 13388
rect 23860 13348 25044 13376
rect 17494 13268 17500 13320
rect 17552 13308 17558 13320
rect 17865 13311 17923 13317
rect 17865 13308 17877 13311
rect 17552 13280 17877 13308
rect 17552 13268 17558 13280
rect 17865 13277 17877 13280
rect 17911 13277 17923 13311
rect 17865 13271 17923 13277
rect 18601 13311 18659 13317
rect 18601 13277 18613 13311
rect 18647 13308 18659 13311
rect 18690 13308 18696 13320
rect 18647 13280 18696 13308
rect 18647 13277 18659 13280
rect 18601 13271 18659 13277
rect 18690 13268 18696 13280
rect 18748 13308 18754 13320
rect 18748 13280 19380 13308
rect 18748 13268 18754 13280
rect 15611 13212 16344 13240
rect 18049 13243 18107 13249
rect 15611 13209 15623 13212
rect 15565 13203 15623 13209
rect 18049 13209 18061 13243
rect 18095 13240 18107 13243
rect 18322 13240 18328 13252
rect 18095 13212 18328 13240
rect 18095 13209 18107 13212
rect 18049 13203 18107 13209
rect 18322 13200 18328 13212
rect 18380 13200 18386 13252
rect 18414 13200 18420 13252
rect 18472 13240 18478 13252
rect 18785 13243 18843 13249
rect 18785 13240 18797 13243
rect 18472 13212 18797 13240
rect 18472 13200 18478 13212
rect 18785 13209 18797 13212
rect 18831 13209 18843 13243
rect 19352 13240 19380 13280
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 20809 13311 20867 13317
rect 20809 13308 20821 13311
rect 19484 13280 20821 13308
rect 19484 13268 19490 13280
rect 20809 13277 20821 13280
rect 20855 13277 20867 13311
rect 20809 13271 20867 13277
rect 21361 13311 21419 13317
rect 21361 13277 21373 13311
rect 21407 13277 21419 13311
rect 21361 13271 21419 13277
rect 20714 13240 20720 13252
rect 19352 13212 20720 13240
rect 18785 13203 18843 13209
rect 20714 13200 20720 13212
rect 20772 13200 20778 13252
rect 13906 13172 13912 13184
rect 12820 13144 13912 13172
rect 13906 13132 13912 13144
rect 13964 13132 13970 13184
rect 14642 13132 14648 13184
rect 14700 13132 14706 13184
rect 15197 13175 15255 13181
rect 15197 13141 15209 13175
rect 15243 13172 15255 13175
rect 15286 13172 15292 13184
rect 15243 13144 15292 13172
rect 15243 13141 15255 13144
rect 15197 13135 15255 13141
rect 15286 13132 15292 13144
rect 15344 13132 15350 13184
rect 15378 13132 15384 13184
rect 15436 13172 15442 13184
rect 15838 13172 15844 13184
rect 15436 13144 15844 13172
rect 15436 13132 15442 13144
rect 15838 13132 15844 13144
rect 15896 13132 15902 13184
rect 21376 13172 21404 13271
rect 21542 13268 21548 13320
rect 21600 13308 21606 13320
rect 21637 13311 21695 13317
rect 21637 13308 21649 13311
rect 21600 13280 21649 13308
rect 21600 13268 21606 13280
rect 21637 13277 21649 13280
rect 21683 13277 21695 13311
rect 21637 13271 21695 13277
rect 22741 13311 22799 13317
rect 22741 13277 22753 13311
rect 22787 13308 22799 13311
rect 23860 13308 23888 13348
rect 25038 13336 25044 13348
rect 25096 13336 25102 13388
rect 22787 13280 23888 13308
rect 24765 13311 24823 13317
rect 22787 13277 22799 13280
rect 22741 13271 22799 13277
rect 24765 13277 24777 13311
rect 24811 13277 24823 13311
rect 24765 13271 24823 13277
rect 23382 13200 23388 13252
rect 23440 13240 23446 13252
rect 24780 13240 24808 13271
rect 23440 13212 24808 13240
rect 23440 13200 23446 13212
rect 21634 13172 21640 13184
rect 21376 13144 21640 13172
rect 21634 13132 21640 13144
rect 21692 13132 21698 13184
rect 24302 13132 24308 13184
rect 24360 13172 24366 13184
rect 25041 13175 25099 13181
rect 25041 13172 25053 13175
rect 24360 13144 25053 13172
rect 24360 13132 24366 13144
rect 25041 13141 25053 13144
rect 25087 13141 25099 13175
rect 25041 13135 25099 13141
rect 1104 13082 25852 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 25852 13082
rect 1104 13008 25852 13030
rect 7742 12928 7748 12980
rect 7800 12968 7806 12980
rect 7837 12971 7895 12977
rect 7837 12968 7849 12971
rect 7800 12940 7849 12968
rect 7800 12928 7806 12940
rect 7837 12937 7849 12940
rect 7883 12937 7895 12971
rect 7837 12931 7895 12937
rect 9033 12971 9091 12977
rect 9033 12937 9045 12971
rect 9079 12968 9091 12971
rect 9214 12968 9220 12980
rect 9079 12940 9220 12968
rect 9079 12937 9091 12940
rect 9033 12931 9091 12937
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 9398 12928 9404 12980
rect 9456 12928 9462 12980
rect 10042 12928 10048 12980
rect 10100 12968 10106 12980
rect 10413 12971 10471 12977
rect 10413 12968 10425 12971
rect 10100 12940 10425 12968
rect 10100 12928 10106 12940
rect 10413 12937 10425 12940
rect 10459 12937 10471 12971
rect 10413 12931 10471 12937
rect 10781 12971 10839 12977
rect 10781 12937 10793 12971
rect 10827 12968 10839 12971
rect 11054 12968 11060 12980
rect 10827 12940 11060 12968
rect 10827 12937 10839 12940
rect 10781 12931 10839 12937
rect 11054 12928 11060 12940
rect 11112 12928 11118 12980
rect 11609 12971 11667 12977
rect 11609 12937 11621 12971
rect 11655 12968 11667 12971
rect 11790 12968 11796 12980
rect 11655 12940 11796 12968
rect 11655 12937 11667 12940
rect 11609 12931 11667 12937
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 11882 12928 11888 12980
rect 11940 12928 11946 12980
rect 11974 12928 11980 12980
rect 12032 12968 12038 12980
rect 12069 12971 12127 12977
rect 12069 12968 12081 12971
rect 12032 12940 12081 12968
rect 12032 12928 12038 12940
rect 12069 12937 12081 12940
rect 12115 12937 12127 12971
rect 12069 12931 12127 12937
rect 12250 12928 12256 12980
rect 12308 12928 12314 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12492 12940 14320 12968
rect 12492 12928 12498 12940
rect 9493 12903 9551 12909
rect 9493 12869 9505 12903
rect 9539 12900 9551 12903
rect 12618 12900 12624 12912
rect 9539 12872 12624 12900
rect 9539 12869 9551 12872
rect 9493 12863 9551 12869
rect 12618 12860 12624 12872
rect 12676 12860 12682 12912
rect 13078 12860 13084 12912
rect 13136 12860 13142 12912
rect 13446 12860 13452 12912
rect 13504 12900 13510 12912
rect 14185 12903 14243 12909
rect 14185 12900 14197 12903
rect 13504 12872 14197 12900
rect 13504 12860 13510 12872
rect 14185 12869 14197 12872
rect 14231 12869 14243 12903
rect 14292 12900 14320 12940
rect 14366 12928 14372 12980
rect 14424 12968 14430 12980
rect 16942 12968 16948 12980
rect 14424 12940 16948 12968
rect 14424 12928 14430 12940
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 17313 12971 17371 12977
rect 17313 12937 17325 12971
rect 17359 12968 17371 12971
rect 17402 12968 17408 12980
rect 17359 12940 17408 12968
rect 17359 12937 17371 12940
rect 17313 12931 17371 12937
rect 17402 12928 17408 12940
rect 17460 12928 17466 12980
rect 18049 12971 18107 12977
rect 18049 12937 18061 12971
rect 18095 12968 18107 12971
rect 18785 12971 18843 12977
rect 18095 12940 18736 12968
rect 18095 12937 18107 12940
rect 18049 12931 18107 12937
rect 18708 12900 18736 12940
rect 18785 12937 18797 12971
rect 18831 12968 18843 12971
rect 19426 12968 19432 12980
rect 18831 12940 19432 12968
rect 18831 12937 18843 12940
rect 18785 12931 18843 12937
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 21266 12968 21272 12980
rect 20088 12940 21272 12968
rect 20088 12900 20116 12940
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 22465 12971 22523 12977
rect 22465 12968 22477 12971
rect 21468 12940 22477 12968
rect 14292 12872 18276 12900
rect 18708 12872 20116 12900
rect 14185 12863 14243 12869
rect 7006 12792 7012 12844
rect 7064 12792 7070 12844
rect 7101 12835 7159 12841
rect 7101 12801 7113 12835
rect 7147 12832 7159 12835
rect 7282 12832 7288 12844
rect 7147 12804 7288 12832
rect 7147 12801 7159 12804
rect 7101 12795 7159 12801
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 8202 12792 8208 12844
rect 8260 12792 8266 12844
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12832 10931 12835
rect 11790 12832 11796 12844
rect 10919 12804 11796 12832
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 11790 12792 11796 12804
rect 11848 12792 11854 12844
rect 12802 12832 12808 12844
rect 11900 12804 12808 12832
rect 6914 12724 6920 12776
rect 6972 12764 6978 12776
rect 7193 12767 7251 12773
rect 7193 12764 7205 12767
rect 6972 12736 7205 12764
rect 6972 12724 6978 12736
rect 7193 12733 7205 12736
rect 7239 12733 7251 12767
rect 7193 12727 7251 12733
rect 7834 12724 7840 12776
rect 7892 12764 7898 12776
rect 8297 12767 8355 12773
rect 8297 12764 8309 12767
rect 7892 12736 8309 12764
rect 7892 12724 7898 12736
rect 8297 12733 8309 12736
rect 8343 12733 8355 12767
rect 8297 12727 8355 12733
rect 8478 12724 8484 12776
rect 8536 12724 8542 12776
rect 9677 12767 9735 12773
rect 9677 12733 9689 12767
rect 9723 12764 9735 12767
rect 9766 12764 9772 12776
rect 9723 12736 9772 12764
rect 9723 12733 9735 12736
rect 9677 12727 9735 12733
rect 9766 12724 9772 12736
rect 9824 12764 9830 12776
rect 9950 12764 9956 12776
rect 9824 12736 9956 12764
rect 9824 12724 9830 12736
rect 9950 12724 9956 12736
rect 10008 12764 10014 12776
rect 10962 12764 10968 12776
rect 10008 12736 10968 12764
rect 10008 12724 10014 12736
rect 10962 12724 10968 12736
rect 11020 12724 11026 12776
rect 11900 12764 11928 12804
rect 12802 12792 12808 12804
rect 12860 12792 12866 12844
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12832 13047 12835
rect 14277 12835 14335 12841
rect 13035 12804 13308 12832
rect 13035 12801 13047 12804
rect 12989 12795 13047 12801
rect 13173 12767 13231 12773
rect 13173 12764 13185 12767
rect 11716 12736 11928 12764
rect 12406 12736 13185 12764
rect 6641 12699 6699 12705
rect 6641 12665 6653 12699
rect 6687 12696 6699 12699
rect 10410 12696 10416 12708
rect 6687 12668 10416 12696
rect 6687 12665 6699 12668
rect 6641 12659 6699 12665
rect 10410 12656 10416 12668
rect 10468 12656 10474 12708
rect 8846 12588 8852 12640
rect 8904 12628 8910 12640
rect 11716 12637 11744 12736
rect 11882 12656 11888 12708
rect 11940 12696 11946 12708
rect 12406 12696 12434 12736
rect 13173 12733 13185 12736
rect 13219 12733 13231 12767
rect 13173 12727 13231 12733
rect 11940 12668 12434 12696
rect 11940 12656 11946 12668
rect 11701 12631 11759 12637
rect 11701 12628 11713 12631
rect 8904 12600 11713 12628
rect 8904 12588 8910 12600
rect 11701 12597 11713 12600
rect 11747 12597 11759 12631
rect 11701 12591 11759 12597
rect 12621 12631 12679 12637
rect 12621 12597 12633 12631
rect 12667 12628 12679 12631
rect 12986 12628 12992 12640
rect 12667 12600 12992 12628
rect 12667 12597 12679 12600
rect 12621 12591 12679 12597
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 13280 12628 13308 12804
rect 14277 12801 14289 12835
rect 14323 12832 14335 12835
rect 15102 12832 15108 12844
rect 14323 12804 15108 12832
rect 14323 12801 14335 12804
rect 14277 12795 14335 12801
rect 15102 12792 15108 12804
rect 15160 12792 15166 12844
rect 15381 12835 15439 12841
rect 15381 12801 15393 12835
rect 15427 12801 15439 12835
rect 15381 12795 15439 12801
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 14090 12764 14096 12776
rect 13872 12736 14096 12764
rect 13872 12724 13878 12736
rect 14090 12724 14096 12736
rect 14148 12764 14154 12776
rect 14369 12767 14427 12773
rect 14369 12764 14381 12767
rect 14148 12736 14381 12764
rect 14148 12724 14154 12736
rect 14369 12733 14381 12736
rect 14415 12733 14427 12767
rect 14369 12727 14427 12733
rect 13538 12628 13544 12640
rect 13280 12600 13544 12628
rect 13538 12588 13544 12600
rect 13596 12588 13602 12640
rect 13817 12631 13875 12637
rect 13817 12597 13829 12631
rect 13863 12628 13875 12631
rect 14366 12628 14372 12640
rect 13863 12600 14372 12628
rect 13863 12597 13875 12600
rect 13817 12591 13875 12597
rect 14366 12588 14372 12600
rect 14424 12588 14430 12640
rect 15010 12588 15016 12640
rect 15068 12588 15074 12640
rect 15396 12628 15424 12795
rect 15470 12792 15476 12844
rect 15528 12792 15534 12844
rect 17218 12792 17224 12844
rect 17276 12792 17282 12844
rect 18248 12841 18276 12872
rect 20622 12860 20628 12912
rect 20680 12900 20686 12912
rect 21177 12903 21235 12909
rect 21177 12900 21189 12903
rect 20680 12872 21189 12900
rect 20680 12860 20686 12872
rect 21177 12869 21189 12872
rect 21223 12900 21235 12903
rect 21468 12900 21496 12940
rect 22465 12937 22477 12940
rect 22511 12937 22523 12971
rect 24302 12968 24308 12980
rect 22465 12931 22523 12937
rect 23216 12940 24308 12968
rect 23216 12900 23244 12940
rect 21223 12872 21496 12900
rect 22480 12872 23244 12900
rect 21223 12869 21235 12872
rect 21177 12863 21235 12869
rect 22480 12844 22508 12872
rect 23290 12860 23296 12912
rect 23348 12900 23354 12912
rect 23385 12903 23443 12909
rect 23385 12900 23397 12903
rect 23348 12872 23397 12900
rect 23348 12860 23354 12872
rect 23385 12869 23397 12872
rect 23431 12869 23443 12903
rect 23768 12900 23796 12940
rect 24302 12928 24308 12940
rect 24360 12968 24366 12980
rect 25133 12971 25191 12977
rect 25133 12968 25145 12971
rect 24360 12940 25145 12968
rect 24360 12928 24366 12940
rect 25133 12937 25145 12940
rect 25179 12937 25191 12971
rect 25133 12931 25191 12937
rect 23768 12872 23874 12900
rect 23385 12863 23443 12869
rect 18233 12835 18291 12841
rect 18233 12801 18245 12835
rect 18279 12801 18291 12835
rect 18233 12795 18291 12801
rect 18782 12792 18788 12844
rect 18840 12832 18846 12844
rect 19153 12836 19211 12841
rect 19076 12835 19211 12836
rect 19076 12832 19165 12835
rect 18840 12808 19165 12832
rect 18840 12804 19104 12808
rect 18840 12792 18846 12804
rect 19153 12801 19165 12808
rect 19199 12801 19211 12835
rect 19153 12795 19211 12801
rect 20165 12835 20223 12841
rect 20165 12801 20177 12835
rect 20211 12832 20223 12835
rect 20806 12832 20812 12844
rect 20211 12804 20812 12832
rect 20211 12801 20223 12804
rect 20165 12795 20223 12801
rect 20806 12792 20812 12804
rect 20864 12792 20870 12844
rect 21082 12792 21088 12844
rect 21140 12792 21146 12844
rect 22094 12832 22100 12844
rect 21284 12804 22100 12832
rect 15562 12724 15568 12776
rect 15620 12764 15626 12776
rect 15838 12764 15844 12776
rect 15620 12736 15844 12764
rect 15620 12724 15626 12736
rect 15838 12724 15844 12736
rect 15896 12724 15902 12776
rect 17497 12767 17555 12773
rect 17497 12733 17509 12767
rect 17543 12764 17555 12767
rect 18874 12764 18880 12776
rect 17543 12736 18880 12764
rect 17543 12733 17555 12736
rect 17497 12727 17555 12733
rect 18874 12724 18880 12736
rect 18932 12724 18938 12776
rect 19242 12724 19248 12776
rect 19300 12724 19306 12776
rect 19429 12767 19487 12773
rect 19429 12733 19441 12767
rect 19475 12764 19487 12767
rect 21284 12764 21312 12804
rect 22094 12792 22100 12804
rect 22152 12792 22158 12844
rect 22186 12792 22192 12844
rect 22244 12792 22250 12844
rect 22462 12792 22468 12844
rect 22520 12792 22526 12844
rect 22830 12792 22836 12844
rect 22888 12832 22894 12844
rect 23109 12835 23167 12841
rect 23109 12832 23121 12835
rect 22888 12804 23121 12832
rect 22888 12792 22894 12804
rect 23109 12801 23121 12804
rect 23155 12801 23167 12835
rect 23109 12795 23167 12801
rect 19475 12736 21312 12764
rect 21361 12767 21419 12773
rect 19475 12733 19487 12736
rect 19429 12727 19487 12733
rect 21361 12733 21373 12767
rect 21407 12764 21419 12767
rect 21407 12736 23244 12764
rect 21407 12733 21419 12736
rect 21361 12727 21419 12733
rect 16853 12699 16911 12705
rect 16853 12665 16865 12699
rect 16899 12696 16911 12699
rect 17126 12696 17132 12708
rect 16899 12668 17132 12696
rect 16899 12665 16911 12668
rect 16853 12659 16911 12665
rect 17126 12656 17132 12668
rect 17184 12656 17190 12708
rect 21174 12696 21180 12708
rect 19306 12668 21180 12696
rect 16117 12631 16175 12637
rect 16117 12628 16129 12631
rect 15396 12600 16129 12628
rect 16117 12597 16129 12600
rect 16163 12628 16175 12631
rect 19306 12628 19334 12668
rect 21174 12656 21180 12668
rect 21232 12656 21238 12708
rect 22002 12656 22008 12708
rect 22060 12656 22066 12708
rect 22554 12656 22560 12708
rect 22612 12696 22618 12708
rect 22612 12668 22876 12696
rect 22612 12656 22618 12668
rect 22848 12640 22876 12668
rect 16163 12600 19334 12628
rect 16163 12597 16175 12600
rect 16117 12591 16175 12597
rect 19426 12588 19432 12640
rect 19484 12628 19490 12640
rect 19981 12631 20039 12637
rect 19981 12628 19993 12631
rect 19484 12600 19993 12628
rect 19484 12588 19490 12600
rect 19981 12597 19993 12600
rect 20027 12597 20039 12631
rect 19981 12591 20039 12597
rect 20717 12631 20775 12637
rect 20717 12597 20729 12631
rect 20763 12628 20775 12631
rect 21910 12628 21916 12640
rect 20763 12600 21916 12628
rect 20763 12597 20775 12600
rect 20717 12591 20775 12597
rect 21910 12588 21916 12600
rect 21968 12588 21974 12640
rect 22094 12588 22100 12640
rect 22152 12628 22158 12640
rect 22462 12628 22468 12640
rect 22152 12600 22468 12628
rect 22152 12588 22158 12600
rect 22462 12588 22468 12600
rect 22520 12628 22526 12640
rect 22649 12631 22707 12637
rect 22649 12628 22661 12631
rect 22520 12600 22661 12628
rect 22520 12588 22526 12600
rect 22649 12597 22661 12600
rect 22695 12597 22707 12631
rect 22649 12591 22707 12597
rect 22830 12588 22836 12640
rect 22888 12588 22894 12640
rect 23216 12628 23244 12736
rect 23382 12628 23388 12640
rect 23216 12600 23388 12628
rect 23382 12588 23388 12600
rect 23440 12628 23446 12640
rect 24857 12631 24915 12637
rect 24857 12628 24869 12631
rect 23440 12600 24869 12628
rect 23440 12588 23446 12600
rect 24857 12597 24869 12600
rect 24903 12597 24915 12631
rect 24857 12591 24915 12597
rect 1104 12538 25852 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 25852 12538
rect 1104 12464 25852 12486
rect 7558 12384 7564 12436
rect 7616 12424 7622 12436
rect 10229 12427 10287 12433
rect 10229 12424 10241 12427
rect 7616 12396 10241 12424
rect 7616 12384 7622 12396
rect 10229 12393 10241 12396
rect 10275 12393 10287 12427
rect 10229 12387 10287 12393
rect 11422 12384 11428 12436
rect 11480 12384 11486 12436
rect 12526 12384 12532 12436
rect 12584 12424 12590 12436
rect 12621 12427 12679 12433
rect 12621 12424 12633 12427
rect 12584 12396 12633 12424
rect 12584 12384 12590 12396
rect 12621 12393 12633 12396
rect 12667 12393 12679 12427
rect 12621 12387 12679 12393
rect 13906 12384 13912 12436
rect 13964 12424 13970 12436
rect 16301 12427 16359 12433
rect 16301 12424 16313 12427
rect 13964 12396 16313 12424
rect 13964 12384 13970 12396
rect 16301 12393 16313 12396
rect 16347 12424 16359 12427
rect 17310 12424 17316 12436
rect 16347 12396 17316 12424
rect 16347 12393 16359 12396
rect 16301 12387 16359 12393
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 18506 12384 18512 12436
rect 18564 12424 18570 12436
rect 18874 12424 18880 12436
rect 18564 12396 18880 12424
rect 18564 12384 18570 12396
rect 18874 12384 18880 12396
rect 18932 12384 18938 12436
rect 21726 12384 21732 12436
rect 21784 12424 21790 12436
rect 22189 12427 22247 12433
rect 22189 12424 22201 12427
rect 21784 12396 22201 12424
rect 21784 12384 21790 12396
rect 22189 12393 22201 12396
rect 22235 12393 22247 12427
rect 22189 12387 22247 12393
rect 24118 12384 24124 12436
rect 24176 12424 24182 12436
rect 24581 12427 24639 12433
rect 24581 12424 24593 12427
rect 24176 12396 24593 12424
rect 24176 12384 24182 12396
rect 24581 12393 24593 12396
rect 24627 12393 24639 12427
rect 24581 12387 24639 12393
rect 12434 12316 12440 12368
rect 12492 12356 12498 12368
rect 14090 12356 14096 12368
rect 12492 12328 14096 12356
rect 12492 12316 12498 12328
rect 14090 12316 14096 12328
rect 14148 12316 14154 12368
rect 14182 12316 14188 12368
rect 14240 12356 14246 12368
rect 14277 12359 14335 12365
rect 14277 12356 14289 12359
rect 14240 12328 14289 12356
rect 14240 12316 14246 12328
rect 14277 12325 14289 12328
rect 14323 12325 14335 12359
rect 14277 12319 14335 12325
rect 15194 12316 15200 12368
rect 15252 12356 15258 12368
rect 15289 12359 15347 12365
rect 15289 12356 15301 12359
rect 15252 12328 15301 12356
rect 15252 12316 15258 12328
rect 15289 12325 15301 12328
rect 15335 12356 15347 12359
rect 18598 12356 18604 12368
rect 15335 12328 18604 12356
rect 15335 12325 15347 12328
rect 15289 12319 15347 12325
rect 18598 12316 18604 12328
rect 18656 12356 18662 12368
rect 18966 12356 18972 12368
rect 18656 12328 18972 12356
rect 18656 12316 18662 12328
rect 18966 12316 18972 12328
rect 19024 12316 19030 12368
rect 22462 12316 22468 12368
rect 22520 12356 22526 12368
rect 22830 12356 22836 12368
rect 22520 12328 22836 12356
rect 22520 12316 22526 12328
rect 22830 12316 22836 12328
rect 22888 12316 22894 12368
rect 7006 12248 7012 12300
rect 7064 12288 7070 12300
rect 7377 12291 7435 12297
rect 7377 12288 7389 12291
rect 7064 12260 7389 12288
rect 7064 12248 7070 12260
rect 7377 12257 7389 12260
rect 7423 12257 7435 12291
rect 7377 12251 7435 12257
rect 8202 12248 8208 12300
rect 8260 12248 8266 12300
rect 9306 12248 9312 12300
rect 9364 12288 9370 12300
rect 10781 12291 10839 12297
rect 10781 12288 10793 12291
rect 9364 12260 10793 12288
rect 9364 12248 9370 12260
rect 10781 12257 10793 12260
rect 10827 12257 10839 12291
rect 10781 12251 10839 12257
rect 11054 12248 11060 12300
rect 11112 12288 11118 12300
rect 11974 12288 11980 12300
rect 11112 12260 11980 12288
rect 11112 12248 11118 12260
rect 11974 12248 11980 12260
rect 12032 12248 12038 12300
rect 13265 12291 13323 12297
rect 12406 12260 12756 12288
rect 11793 12223 11851 12229
rect 11793 12189 11805 12223
rect 11839 12220 11851 12223
rect 12406 12220 12434 12260
rect 11839 12192 12434 12220
rect 11839 12189 11851 12192
rect 11793 12183 11851 12189
rect 10689 12155 10747 12161
rect 10689 12121 10701 12155
rect 10735 12152 10747 12155
rect 12526 12152 12532 12164
rect 10735 12124 12532 12152
rect 10735 12121 10747 12124
rect 10689 12115 10747 12121
rect 12526 12112 12532 12124
rect 12584 12112 12590 12164
rect 12728 12152 12756 12260
rect 13265 12257 13277 12291
rect 13311 12288 13323 12291
rect 13722 12288 13728 12300
rect 13311 12260 13728 12288
rect 13311 12257 13323 12260
rect 13265 12251 13323 12257
rect 13722 12248 13728 12260
rect 13780 12288 13786 12300
rect 14829 12291 14887 12297
rect 14829 12288 14841 12291
rect 13780 12260 14841 12288
rect 13780 12248 13786 12260
rect 14829 12257 14841 12260
rect 14875 12257 14887 12291
rect 14829 12251 14887 12257
rect 15565 12291 15623 12297
rect 15565 12257 15577 12291
rect 15611 12288 15623 12291
rect 15838 12288 15844 12300
rect 15611 12260 15844 12288
rect 15611 12257 15623 12260
rect 15565 12251 15623 12257
rect 15838 12248 15844 12260
rect 15896 12248 15902 12300
rect 16850 12248 16856 12300
rect 16908 12288 16914 12300
rect 18693 12291 18751 12297
rect 16908 12260 17448 12288
rect 16908 12248 16914 12260
rect 12802 12180 12808 12232
rect 12860 12220 12866 12232
rect 13081 12223 13139 12229
rect 13081 12220 13093 12223
rect 12860 12192 13093 12220
rect 12860 12180 12866 12192
rect 13081 12189 13093 12192
rect 13127 12220 13139 12223
rect 13446 12220 13452 12232
rect 13127 12192 13452 12220
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 13446 12180 13452 12192
rect 13504 12220 13510 12232
rect 13633 12223 13691 12229
rect 13633 12220 13645 12223
rect 13504 12192 13645 12220
rect 13504 12180 13510 12192
rect 13633 12189 13645 12192
rect 13679 12189 13691 12223
rect 13633 12183 13691 12189
rect 13909 12223 13967 12229
rect 13909 12189 13921 12223
rect 13955 12220 13967 12223
rect 14642 12220 14648 12232
rect 13955 12192 14648 12220
rect 13955 12189 13967 12192
rect 13909 12183 13967 12189
rect 14642 12180 14648 12192
rect 14700 12220 14706 12232
rect 14737 12223 14795 12229
rect 14737 12220 14749 12223
rect 14700 12192 14749 12220
rect 14700 12180 14706 12192
rect 14737 12189 14749 12192
rect 14783 12189 14795 12223
rect 14737 12183 14795 12189
rect 17310 12180 17316 12232
rect 17368 12180 17374 12232
rect 17420 12220 17448 12260
rect 18693 12257 18705 12291
rect 18739 12288 18751 12291
rect 18782 12288 18788 12300
rect 18739 12260 18788 12288
rect 18739 12257 18751 12260
rect 18693 12251 18751 12257
rect 18782 12248 18788 12260
rect 18840 12248 18846 12300
rect 19981 12291 20039 12297
rect 19981 12288 19993 12291
rect 19260 12260 19993 12288
rect 19260 12232 19288 12260
rect 19981 12257 19993 12260
rect 20027 12257 20039 12291
rect 19981 12251 20039 12257
rect 20438 12248 20444 12300
rect 20496 12248 20502 12300
rect 20717 12291 20775 12297
rect 20717 12257 20729 12291
rect 20763 12288 20775 12291
rect 21266 12288 21272 12300
rect 20763 12260 21272 12288
rect 20763 12257 20775 12260
rect 20717 12251 20775 12257
rect 21266 12248 21272 12260
rect 21324 12248 21330 12300
rect 19242 12220 19248 12232
rect 17420 12192 19248 12220
rect 19242 12180 19248 12192
rect 19300 12180 19306 12232
rect 19521 12223 19579 12229
rect 19521 12189 19533 12223
rect 19567 12220 19579 12223
rect 20162 12220 20168 12232
rect 19567 12192 20168 12220
rect 19567 12189 19579 12192
rect 19521 12183 19579 12189
rect 20162 12180 20168 12192
rect 20220 12180 20226 12232
rect 22833 12223 22891 12229
rect 22833 12189 22845 12223
rect 22879 12189 22891 12223
rect 22833 12183 22891 12189
rect 15010 12152 15016 12164
rect 12728 12124 13676 12152
rect 8478 12044 8484 12096
rect 8536 12084 8542 12096
rect 8941 12087 8999 12093
rect 8941 12084 8953 12087
rect 8536 12056 8953 12084
rect 8536 12044 8542 12056
rect 8941 12053 8953 12056
rect 8987 12084 8999 12087
rect 9398 12084 9404 12096
rect 8987 12056 9404 12084
rect 8987 12053 8999 12056
rect 8941 12047 8999 12053
rect 9398 12044 9404 12056
rect 9456 12044 9462 12096
rect 10594 12044 10600 12096
rect 10652 12044 10658 12096
rect 11885 12087 11943 12093
rect 11885 12053 11897 12087
rect 11931 12084 11943 12087
rect 12434 12084 12440 12096
rect 11931 12056 12440 12084
rect 11931 12053 11943 12056
rect 11885 12047 11943 12053
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 12989 12087 13047 12093
rect 12989 12053 13001 12087
rect 13035 12084 13047 12087
rect 13262 12084 13268 12096
rect 13035 12056 13268 12084
rect 13035 12053 13047 12056
rect 12989 12047 13047 12053
rect 13262 12044 13268 12056
rect 13320 12044 13326 12096
rect 13648 12084 13676 12124
rect 13924 12124 15016 12152
rect 13924 12084 13952 12124
rect 15010 12112 15016 12124
rect 15068 12112 15074 12164
rect 16942 12112 16948 12164
rect 17000 12152 17006 12164
rect 18049 12155 18107 12161
rect 18049 12152 18061 12155
rect 17000 12124 18061 12152
rect 17000 12112 17006 12124
rect 18049 12121 18061 12124
rect 18095 12121 18107 12155
rect 18049 12115 18107 12121
rect 19702 12112 19708 12164
rect 19760 12152 19766 12164
rect 22002 12152 22008 12164
rect 19760 12124 21128 12152
rect 21942 12124 22008 12152
rect 19760 12112 19766 12124
rect 13648 12056 13952 12084
rect 14645 12087 14703 12093
rect 14645 12053 14657 12087
rect 14691 12084 14703 12087
rect 15562 12084 15568 12096
rect 14691 12056 15568 12084
rect 14691 12053 14703 12056
rect 14645 12047 14703 12053
rect 15562 12044 15568 12056
rect 15620 12084 15626 12096
rect 15657 12087 15715 12093
rect 15657 12084 15669 12087
rect 15620 12056 15669 12084
rect 15620 12044 15626 12056
rect 15657 12053 15669 12056
rect 15703 12084 15715 12087
rect 16022 12084 16028 12096
rect 15703 12056 16028 12084
rect 15703 12053 15715 12056
rect 15657 12047 15715 12053
rect 16022 12044 16028 12056
rect 16080 12044 16086 12096
rect 16669 12087 16727 12093
rect 16669 12053 16681 12087
rect 16715 12084 16727 12087
rect 18414 12084 18420 12096
rect 16715 12056 18420 12084
rect 16715 12053 16727 12056
rect 16669 12047 16727 12053
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 18966 12044 18972 12096
rect 19024 12084 19030 12096
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 19024 12056 19625 12084
rect 19024 12044 19030 12056
rect 19613 12053 19625 12056
rect 19659 12053 19671 12087
rect 21100 12084 21128 12124
rect 22002 12112 22008 12124
rect 22060 12112 22066 12164
rect 22848 12152 22876 12183
rect 24486 12180 24492 12232
rect 24544 12220 24550 12232
rect 24765 12223 24823 12229
rect 24765 12220 24777 12223
rect 24544 12192 24777 12220
rect 24544 12180 24550 12192
rect 24765 12189 24777 12192
rect 24811 12189 24823 12223
rect 24765 12183 24823 12189
rect 23566 12152 23572 12164
rect 22848 12124 23572 12152
rect 23566 12112 23572 12124
rect 23624 12112 23630 12164
rect 23845 12155 23903 12161
rect 23845 12121 23857 12155
rect 23891 12152 23903 12155
rect 24946 12152 24952 12164
rect 23891 12124 24952 12152
rect 23891 12121 23903 12124
rect 23845 12115 23903 12121
rect 24946 12112 24952 12124
rect 25004 12112 25010 12164
rect 21726 12084 21732 12096
rect 21100 12056 21732 12084
rect 19613 12047 19671 12053
rect 21726 12044 21732 12056
rect 21784 12044 21790 12096
rect 1104 11994 25852 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 25852 11994
rect 1104 11920 25852 11942
rect 3694 11840 3700 11892
rect 3752 11880 3758 11892
rect 9033 11883 9091 11889
rect 3752 11852 8984 11880
rect 3752 11840 3758 11852
rect 8956 11812 8984 11852
rect 9033 11849 9045 11883
rect 9079 11880 9091 11883
rect 9306 11880 9312 11892
rect 9079 11852 9312 11880
rect 9079 11849 9091 11852
rect 9033 11843 9091 11849
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 9861 11883 9919 11889
rect 9861 11880 9873 11883
rect 9732 11852 9873 11880
rect 9732 11840 9738 11852
rect 9861 11849 9873 11852
rect 9907 11849 9919 11883
rect 9861 11843 9919 11849
rect 10229 11883 10287 11889
rect 10229 11849 10241 11883
rect 10275 11880 10287 11883
rect 10870 11880 10876 11892
rect 10275 11852 10876 11880
rect 10275 11849 10287 11852
rect 10229 11843 10287 11849
rect 9585 11815 9643 11821
rect 9585 11812 9597 11815
rect 8956 11784 9597 11812
rect 9585 11781 9597 11784
rect 9631 11812 9643 11815
rect 10244 11812 10272 11843
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 11885 11883 11943 11889
rect 11885 11849 11897 11883
rect 11931 11880 11943 11883
rect 12710 11880 12716 11892
rect 11931 11852 12716 11880
rect 11931 11849 11943 11852
rect 11885 11843 11943 11849
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 13081 11883 13139 11889
rect 13081 11849 13093 11883
rect 13127 11880 13139 11883
rect 13354 11880 13360 11892
rect 13127 11852 13360 11880
rect 13127 11849 13139 11852
rect 13081 11843 13139 11849
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 13446 11840 13452 11892
rect 13504 11840 13510 11892
rect 13541 11883 13599 11889
rect 13541 11849 13553 11883
rect 13587 11880 13599 11883
rect 13906 11880 13912 11892
rect 13587 11852 13912 11880
rect 13587 11849 13599 11852
rect 13541 11843 13599 11849
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 13998 11840 14004 11892
rect 14056 11880 14062 11892
rect 14277 11883 14335 11889
rect 14277 11880 14289 11883
rect 14056 11852 14289 11880
rect 14056 11840 14062 11852
rect 14277 11849 14289 11852
rect 14323 11849 14335 11883
rect 14277 11843 14335 11849
rect 14737 11883 14795 11889
rect 14737 11849 14749 11883
rect 14783 11880 14795 11883
rect 14826 11880 14832 11892
rect 14783 11852 14832 11880
rect 14783 11849 14795 11852
rect 14737 11843 14795 11849
rect 14826 11840 14832 11852
rect 14884 11840 14890 11892
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 16758 11880 16764 11892
rect 15252 11852 16764 11880
rect 15252 11840 15258 11852
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 17034 11840 17040 11892
rect 17092 11880 17098 11892
rect 17313 11883 17371 11889
rect 17313 11880 17325 11883
rect 17092 11852 17325 11880
rect 17092 11840 17098 11852
rect 17313 11849 17325 11852
rect 17359 11849 17371 11883
rect 17313 11843 17371 11849
rect 18049 11883 18107 11889
rect 18049 11849 18061 11883
rect 18095 11849 18107 11883
rect 18049 11843 18107 11849
rect 9631 11784 10272 11812
rect 10321 11815 10379 11821
rect 9631 11781 9643 11784
rect 9585 11775 9643 11781
rect 10321 11781 10333 11815
rect 10367 11812 10379 11815
rect 14182 11812 14188 11824
rect 10367 11784 14188 11812
rect 10367 11781 10379 11784
rect 10321 11775 10379 11781
rect 14182 11772 14188 11784
rect 14240 11772 14246 11824
rect 15010 11772 15016 11824
rect 15068 11812 15074 11824
rect 18064 11812 18092 11843
rect 18414 11840 18420 11892
rect 18472 11840 18478 11892
rect 19518 11840 19524 11892
rect 19576 11880 19582 11892
rect 19576 11852 20116 11880
rect 19576 11840 19582 11852
rect 19978 11812 19984 11824
rect 15068 11784 17908 11812
rect 18064 11784 19984 11812
rect 15068 11772 15074 11784
rect 8662 11704 8668 11756
rect 8720 11744 8726 11756
rect 9398 11744 9404 11756
rect 8720 11716 9404 11744
rect 8720 11704 8726 11716
rect 9398 11704 9404 11716
rect 9456 11704 9462 11756
rect 9490 11704 9496 11756
rect 9548 11744 9554 11756
rect 11238 11744 11244 11756
rect 9548 11716 11244 11744
rect 9548 11704 9554 11716
rect 11238 11704 11244 11716
rect 11296 11704 11302 11756
rect 11609 11747 11667 11753
rect 11609 11713 11621 11747
rect 11655 11744 11667 11747
rect 12253 11747 12311 11753
rect 12253 11744 12265 11747
rect 11655 11716 12265 11744
rect 11655 11713 11667 11716
rect 11609 11707 11667 11713
rect 12253 11713 12265 11716
rect 12299 11744 12311 11747
rect 13998 11744 14004 11756
rect 12299 11716 14004 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 13998 11704 14004 11716
rect 14056 11704 14062 11756
rect 14645 11747 14703 11753
rect 14645 11713 14657 11747
rect 14691 11744 14703 11747
rect 15102 11744 15108 11756
rect 14691 11716 15108 11744
rect 14691 11713 14703 11716
rect 14645 11707 14703 11713
rect 15102 11704 15108 11716
rect 15160 11744 15166 11756
rect 15378 11744 15384 11756
rect 15160 11716 15384 11744
rect 15160 11704 15166 11716
rect 15378 11704 15384 11716
rect 15436 11704 15442 11756
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11744 15623 11747
rect 15654 11744 15660 11756
rect 15611 11716 15660 11744
rect 15611 11713 15623 11716
rect 15565 11707 15623 11713
rect 15654 11704 15660 11716
rect 15712 11744 15718 11756
rect 16114 11744 16120 11756
rect 15712 11716 16120 11744
rect 15712 11704 15718 11716
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 16574 11704 16580 11756
rect 16632 11744 16638 11756
rect 17221 11747 17279 11753
rect 17221 11744 17233 11747
rect 16632 11716 17233 11744
rect 16632 11704 16638 11716
rect 17221 11713 17233 11716
rect 17267 11713 17279 11747
rect 17221 11707 17279 11713
rect 7285 11679 7343 11685
rect 7285 11645 7297 11679
rect 7331 11645 7343 11679
rect 7285 11639 7343 11645
rect 7561 11679 7619 11685
rect 7561 11645 7573 11679
rect 7607 11676 7619 11679
rect 10413 11679 10471 11685
rect 7607 11648 10272 11676
rect 7607 11645 7619 11648
rect 7561 11639 7619 11645
rect 7300 11540 7328 11639
rect 10244 11608 10272 11648
rect 10413 11645 10425 11679
rect 10459 11645 10471 11679
rect 11256 11676 11284 11704
rect 17880 11688 17908 11784
rect 19978 11772 19984 11784
rect 20036 11772 20042 11824
rect 20088 11812 20116 11852
rect 20162 11840 20168 11892
rect 20220 11880 20226 11892
rect 21177 11883 21235 11889
rect 21177 11880 21189 11883
rect 20220 11852 21189 11880
rect 20220 11840 20226 11852
rect 21177 11849 21189 11852
rect 21223 11880 21235 11883
rect 24394 11880 24400 11892
rect 21223 11852 24400 11880
rect 21223 11849 21235 11852
rect 21177 11843 21235 11849
rect 24394 11840 24400 11852
rect 24452 11840 24458 11892
rect 21361 11815 21419 11821
rect 21361 11812 21373 11815
rect 20088 11784 21373 11812
rect 21361 11781 21373 11784
rect 21407 11781 21419 11815
rect 21361 11775 21419 11781
rect 23293 11815 23351 11821
rect 23293 11781 23305 11815
rect 23339 11812 23351 11815
rect 24854 11812 24860 11824
rect 23339 11784 24860 11812
rect 23339 11781 23351 11784
rect 23293 11775 23351 11781
rect 24854 11772 24860 11784
rect 24912 11772 24918 11824
rect 19337 11747 19395 11753
rect 19337 11713 19349 11747
rect 19383 11744 19395 11747
rect 19518 11744 19524 11756
rect 19383 11716 19524 11744
rect 19383 11713 19395 11716
rect 19337 11707 19395 11713
rect 19518 11704 19524 11716
rect 19576 11704 19582 11756
rect 20070 11704 20076 11756
rect 20128 11744 20134 11756
rect 22281 11747 22339 11753
rect 20128 11716 21496 11744
rect 20128 11704 20134 11716
rect 12345 11679 12403 11685
rect 12345 11676 12357 11679
rect 11256 11648 12357 11676
rect 10413 11639 10471 11645
rect 12345 11645 12357 11648
rect 12391 11645 12403 11679
rect 12345 11639 12403 11645
rect 10428 11608 10456 11639
rect 12434 11636 12440 11688
rect 12492 11636 12498 11688
rect 13722 11636 13728 11688
rect 13780 11676 13786 11688
rect 14829 11679 14887 11685
rect 14829 11676 14841 11679
rect 13780 11648 14841 11676
rect 13780 11636 13786 11648
rect 14829 11645 14841 11648
rect 14875 11645 14887 11679
rect 14829 11639 14887 11645
rect 16666 11636 16672 11688
rect 16724 11676 16730 11688
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 16724 11648 17417 11676
rect 16724 11636 16730 11648
rect 17405 11645 17417 11648
rect 17451 11645 17463 11679
rect 17405 11639 17463 11645
rect 17862 11636 17868 11688
rect 17920 11676 17926 11688
rect 18509 11679 18567 11685
rect 18509 11676 18521 11679
rect 17920 11648 18521 11676
rect 17920 11636 17926 11648
rect 18509 11645 18521 11648
rect 18555 11645 18567 11679
rect 18509 11639 18567 11645
rect 18693 11679 18751 11685
rect 18693 11645 18705 11679
rect 18739 11676 18751 11679
rect 19702 11676 19708 11688
rect 18739 11648 19708 11676
rect 18739 11645 18751 11648
rect 18693 11639 18751 11645
rect 19702 11636 19708 11648
rect 19760 11636 19766 11688
rect 19978 11636 19984 11688
rect 20036 11676 20042 11688
rect 20717 11679 20775 11685
rect 20717 11676 20729 11679
rect 20036 11648 20729 11676
rect 20036 11636 20042 11648
rect 20717 11645 20729 11648
rect 20763 11645 20775 11679
rect 21468 11676 21496 11716
rect 22281 11713 22293 11747
rect 22327 11744 22339 11747
rect 23750 11744 23756 11756
rect 22327 11716 23756 11744
rect 22327 11713 22339 11716
rect 22281 11707 22339 11713
rect 23750 11704 23756 11716
rect 23808 11704 23814 11756
rect 24121 11747 24179 11753
rect 24121 11713 24133 11747
rect 24167 11744 24179 11747
rect 24946 11744 24952 11756
rect 24167 11716 24952 11744
rect 24167 11713 24179 11716
rect 24121 11707 24179 11713
rect 24946 11704 24952 11716
rect 25004 11704 25010 11756
rect 21637 11679 21695 11685
rect 21637 11676 21649 11679
rect 21468 11648 21649 11676
rect 20717 11639 20775 11645
rect 21637 11645 21649 11648
rect 21683 11676 21695 11679
rect 21683 11648 21864 11676
rect 21683 11645 21695 11648
rect 21637 11639 21695 11645
rect 11054 11608 11060 11620
rect 10244 11580 11060 11608
rect 11054 11568 11060 11580
rect 11112 11568 11118 11620
rect 16853 11611 16911 11617
rect 14936 11580 15608 11608
rect 8294 11540 8300 11552
rect 7300 11512 8300 11540
rect 8294 11500 8300 11512
rect 8352 11540 8358 11552
rect 8938 11540 8944 11552
rect 8352 11512 8944 11540
rect 8352 11500 8358 11512
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 9398 11500 9404 11552
rect 9456 11540 9462 11552
rect 10410 11540 10416 11552
rect 9456 11512 10416 11540
rect 9456 11500 9462 11512
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 11790 11500 11796 11552
rect 11848 11540 11854 11552
rect 14936 11540 14964 11580
rect 11848 11512 14964 11540
rect 15580 11540 15608 11580
rect 16853 11577 16865 11611
rect 16899 11608 16911 11611
rect 21726 11608 21732 11620
rect 16899 11580 21732 11608
rect 16899 11577 16911 11580
rect 16853 11571 16911 11577
rect 21726 11568 21732 11580
rect 21784 11568 21790 11620
rect 21836 11608 21864 11648
rect 24762 11636 24768 11688
rect 24820 11636 24826 11688
rect 25774 11608 25780 11620
rect 21836 11580 25780 11608
rect 25774 11568 25780 11580
rect 25832 11568 25838 11620
rect 17218 11540 17224 11552
rect 15580 11512 17224 11540
rect 11848 11500 11854 11512
rect 17218 11500 17224 11512
rect 17276 11500 17282 11552
rect 18506 11500 18512 11552
rect 18564 11540 18570 11552
rect 19150 11540 19156 11552
rect 18564 11512 19156 11540
rect 18564 11500 18570 11512
rect 19150 11500 19156 11512
rect 19208 11500 19214 11552
rect 19426 11500 19432 11552
rect 19484 11500 19490 11552
rect 20165 11543 20223 11549
rect 20165 11509 20177 11543
rect 20211 11540 20223 11543
rect 21358 11540 21364 11552
rect 20211 11512 21364 11540
rect 20211 11509 20223 11512
rect 20165 11503 20223 11509
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 22278 11500 22284 11552
rect 22336 11540 22342 11552
rect 23290 11540 23296 11552
rect 22336 11512 23296 11540
rect 22336 11500 22342 11512
rect 23290 11500 23296 11512
rect 23348 11500 23354 11552
rect 1104 11450 25852 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 25852 11450
rect 1104 11376 25852 11398
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 12621 11339 12679 11345
rect 12621 11336 12633 11339
rect 10652 11308 12633 11336
rect 10652 11296 10658 11308
rect 12621 11305 12633 11308
rect 12667 11305 12679 11339
rect 15286 11336 15292 11348
rect 12621 11299 12679 11305
rect 13004 11308 15292 11336
rect 11425 11271 11483 11277
rect 11425 11237 11437 11271
rect 11471 11268 11483 11271
rect 12802 11268 12808 11280
rect 11471 11240 12808 11268
rect 11471 11237 11483 11240
rect 11425 11231 11483 11237
rect 12802 11228 12808 11240
rect 12860 11228 12866 11280
rect 12894 11228 12900 11280
rect 12952 11228 12958 11280
rect 9401 11203 9459 11209
rect 9401 11169 9413 11203
rect 9447 11200 9459 11203
rect 12069 11203 12127 11209
rect 12069 11200 12081 11203
rect 9447 11172 12081 11200
rect 9447 11169 9459 11172
rect 9401 11163 9459 11169
rect 12069 11169 12081 11172
rect 12115 11200 12127 11203
rect 12158 11200 12164 11212
rect 12115 11172 12164 11200
rect 12115 11169 12127 11172
rect 12069 11163 12127 11169
rect 12158 11160 12164 11172
rect 12216 11160 12222 11212
rect 12912 11200 12940 11228
rect 12268 11172 12940 11200
rect 9030 11092 9036 11144
rect 9088 11132 9094 11144
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 9088 11104 9137 11132
rect 9088 11092 9094 11104
rect 9125 11101 9137 11104
rect 9171 11101 9183 11135
rect 9125 11095 9183 11101
rect 11054 11092 11060 11144
rect 11112 11132 11118 11144
rect 12268 11132 12296 11172
rect 11112 11104 12296 11132
rect 11112 11092 11118 11104
rect 12526 11092 12532 11144
rect 12584 11132 12590 11144
rect 12894 11132 12900 11144
rect 12584 11104 12900 11132
rect 12584 11092 12590 11104
rect 12894 11092 12900 11104
rect 12952 11092 12958 11144
rect 13004 11141 13032 11308
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 15378 11296 15384 11348
rect 15436 11336 15442 11348
rect 16298 11336 16304 11348
rect 15436 11308 16304 11336
rect 15436 11296 15442 11308
rect 16298 11296 16304 11308
rect 16356 11296 16362 11348
rect 17218 11296 17224 11348
rect 17276 11336 17282 11348
rect 21818 11336 21824 11348
rect 17276 11308 21824 11336
rect 17276 11296 17282 11308
rect 21818 11296 21824 11308
rect 21876 11296 21882 11348
rect 22097 11339 22155 11345
rect 22097 11305 22109 11339
rect 22143 11336 22155 11339
rect 22143 11308 22692 11336
rect 22143 11305 22155 11308
rect 22097 11299 22155 11305
rect 13078 11228 13084 11280
rect 13136 11228 13142 11280
rect 13354 11228 13360 11280
rect 13412 11268 13418 11280
rect 13412 11240 13676 11268
rect 13412 11228 13418 11240
rect 13096 11200 13124 11228
rect 13265 11203 13323 11209
rect 13265 11200 13277 11203
rect 13096 11172 13277 11200
rect 13265 11169 13277 11172
rect 13311 11200 13323 11203
rect 13538 11200 13544 11212
rect 13311 11172 13544 11200
rect 13311 11169 13323 11172
rect 13265 11163 13323 11169
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 13648 11141 13676 11240
rect 13998 11228 14004 11280
rect 14056 11268 14062 11280
rect 14182 11268 14188 11280
rect 14056 11240 14188 11268
rect 14056 11228 14062 11240
rect 14182 11228 14188 11240
rect 14240 11268 14246 11280
rect 14734 11268 14740 11280
rect 14240 11240 14740 11268
rect 14240 11228 14246 11240
rect 14734 11228 14740 11240
rect 14792 11228 14798 11280
rect 16666 11228 16672 11280
rect 16724 11228 16730 11280
rect 17862 11228 17868 11280
rect 17920 11228 17926 11280
rect 18141 11271 18199 11277
rect 18141 11237 18153 11271
rect 18187 11268 18199 11271
rect 20622 11268 20628 11280
rect 18187 11240 20628 11268
rect 18187 11237 18199 11240
rect 18141 11231 18199 11237
rect 20622 11228 20628 11240
rect 20680 11228 20686 11280
rect 21545 11271 21603 11277
rect 21545 11237 21557 11271
rect 21591 11268 21603 11271
rect 22554 11268 22560 11280
rect 21591 11240 22560 11268
rect 21591 11237 21603 11240
rect 21545 11231 21603 11237
rect 22554 11228 22560 11240
rect 22612 11228 22618 11280
rect 22664 11268 22692 11308
rect 23566 11296 23572 11348
rect 23624 11336 23630 11348
rect 25041 11339 25099 11345
rect 25041 11336 25053 11339
rect 23624 11308 25053 11336
rect 23624 11296 23630 11308
rect 25041 11305 25053 11308
rect 25087 11305 25099 11339
rect 25041 11299 25099 11305
rect 25498 11268 25504 11280
rect 22664 11240 25504 11268
rect 14921 11203 14979 11209
rect 14921 11169 14933 11203
rect 14967 11200 14979 11203
rect 16942 11200 16948 11212
rect 14967 11172 16948 11200
rect 14967 11169 14979 11172
rect 14921 11163 14979 11169
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 18598 11160 18604 11212
rect 18656 11160 18662 11212
rect 18785 11203 18843 11209
rect 18785 11169 18797 11203
rect 18831 11200 18843 11203
rect 20257 11203 20315 11209
rect 18831 11172 20208 11200
rect 18831 11169 18843 11172
rect 18785 11163 18843 11169
rect 12989 11135 13047 11141
rect 12989 11101 13001 11135
rect 13035 11101 13047 11135
rect 12989 11095 13047 11101
rect 13633 11135 13691 11141
rect 13633 11101 13645 11135
rect 13679 11132 13691 11135
rect 13679 11104 14964 11132
rect 13679 11101 13691 11104
rect 13633 11095 13691 11101
rect 10410 11024 10416 11076
rect 10468 11024 10474 11076
rect 12250 11064 12256 11076
rect 11808 11036 12256 11064
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 10870 10996 10876 11008
rect 9732 10968 10876 10996
rect 9732 10956 9738 10968
rect 10870 10956 10876 10968
rect 10928 10956 10934 11008
rect 11238 10956 11244 11008
rect 11296 10996 11302 11008
rect 11808 11005 11836 11036
rect 12250 11024 12256 11036
rect 12308 11024 12314 11076
rect 13081 11067 13139 11073
rect 12360 11036 13032 11064
rect 11793 10999 11851 11005
rect 11793 10996 11805 10999
rect 11296 10968 11805 10996
rect 11296 10956 11302 10968
rect 11793 10965 11805 10968
rect 11839 10965 11851 10999
rect 11793 10959 11851 10965
rect 11885 10999 11943 11005
rect 11885 10965 11897 10999
rect 11931 10996 11943 10999
rect 12360 10996 12388 11036
rect 11931 10968 12388 10996
rect 13004 10996 13032 11036
rect 13081 11033 13093 11067
rect 13127 11064 13139 11067
rect 13722 11064 13728 11076
rect 13127 11036 13728 11064
rect 13127 11033 13139 11036
rect 13081 11027 13139 11033
rect 13722 11024 13728 11036
rect 13780 11024 13786 11076
rect 13909 11067 13967 11073
rect 13909 11064 13921 11067
rect 13832 11036 13921 11064
rect 13832 10996 13860 11036
rect 13909 11033 13921 11036
rect 13955 11064 13967 11067
rect 13998 11064 14004 11076
rect 13955 11036 14004 11064
rect 13955 11033 13967 11036
rect 13909 11027 13967 11033
rect 13998 11024 14004 11036
rect 14056 11024 14062 11076
rect 14936 11064 14964 11104
rect 16206 11092 16212 11144
rect 16264 11132 16270 11144
rect 17037 11135 17095 11141
rect 17037 11132 17049 11135
rect 16264 11104 17049 11132
rect 16264 11092 16270 11104
rect 17037 11101 17049 11104
rect 17083 11132 17095 11135
rect 17494 11132 17500 11144
rect 17083 11104 17500 11132
rect 17083 11101 17095 11104
rect 17037 11095 17095 11101
rect 17494 11092 17500 11104
rect 17552 11092 17558 11144
rect 18616 11132 18644 11160
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 18616 11104 19257 11132
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 19978 11092 19984 11144
rect 20036 11092 20042 11144
rect 20180 11132 20208 11172
rect 20257 11169 20269 11203
rect 20303 11200 20315 11203
rect 20990 11200 20996 11212
rect 20303 11172 20996 11200
rect 20303 11169 20315 11172
rect 20257 11163 20315 11169
rect 20990 11160 20996 11172
rect 21048 11160 21054 11212
rect 22664 11200 22692 11240
rect 25498 11228 25504 11240
rect 25556 11228 25562 11280
rect 21652 11172 22692 11200
rect 20714 11132 20720 11144
rect 20180 11104 20720 11132
rect 20714 11092 20720 11104
rect 20772 11092 20778 11144
rect 20901 11135 20959 11141
rect 20901 11101 20913 11135
rect 20947 11132 20959 11135
rect 21174 11132 21180 11144
rect 20947 11104 21180 11132
rect 20947 11101 20959 11104
rect 20901 11095 20959 11101
rect 21174 11092 21180 11104
rect 21232 11132 21238 11144
rect 21652 11132 21680 11172
rect 23290 11160 23296 11212
rect 23348 11160 23354 11212
rect 21232 11104 21680 11132
rect 21232 11092 21238 11104
rect 21726 11092 21732 11144
rect 21784 11092 21790 11144
rect 21818 11092 21824 11144
rect 21876 11132 21882 11144
rect 22278 11132 22284 11144
rect 21876 11104 22284 11132
rect 21876 11092 21882 11104
rect 22278 11092 22284 11104
rect 22336 11092 22342 11144
rect 22833 11135 22891 11141
rect 22833 11101 22845 11135
rect 22879 11101 22891 11135
rect 22833 11095 22891 11101
rect 14936 11036 15148 11064
rect 13004 10968 13860 10996
rect 11931 10965 11943 10968
rect 11885 10959 11943 10965
rect 14274 10956 14280 11008
rect 14332 10956 14338 11008
rect 15120 10996 15148 11036
rect 15194 11024 15200 11076
rect 15252 11024 15258 11076
rect 15286 11024 15292 11076
rect 15344 11024 15350 11076
rect 16868 11036 17080 11064
rect 15304 10996 15332 11024
rect 15120 10968 15332 10996
rect 15470 10956 15476 11008
rect 15528 10996 15534 11008
rect 16868 10996 16896 11036
rect 15528 10968 16896 10996
rect 17052 10996 17080 11036
rect 17402 11024 17408 11076
rect 17460 11064 17466 11076
rect 17589 11067 17647 11073
rect 17589 11064 17601 11067
rect 17460 11036 17601 11064
rect 17460 11024 17466 11036
rect 17589 11033 17601 11036
rect 17635 11064 17647 11067
rect 18509 11067 18567 11073
rect 18509 11064 18521 11067
rect 17635 11036 18521 11064
rect 17635 11033 17647 11036
rect 17589 11027 17647 11033
rect 18509 11033 18521 11036
rect 18555 11033 18567 11067
rect 20806 11064 20812 11076
rect 18509 11027 18567 11033
rect 19628 11036 20812 11064
rect 19334 10996 19340 11008
rect 17052 10968 19340 10996
rect 15528 10956 15534 10968
rect 19334 10956 19340 10968
rect 19392 10956 19398 11008
rect 19628 11005 19656 11036
rect 20806 11024 20812 11036
rect 20864 11024 20870 11076
rect 20990 11024 20996 11076
rect 21048 11064 21054 11076
rect 21085 11067 21143 11073
rect 21085 11064 21097 11067
rect 21048 11036 21097 11064
rect 21048 11024 21054 11036
rect 21085 11033 21097 11036
rect 21131 11033 21143 11067
rect 22848 11064 22876 11095
rect 23934 11092 23940 11144
rect 23992 11132 23998 11144
rect 25225 11135 25283 11141
rect 25225 11132 25237 11135
rect 23992 11104 25237 11132
rect 23992 11092 23998 11104
rect 25225 11101 25237 11104
rect 25271 11101 25283 11135
rect 25225 11095 25283 11101
rect 25038 11064 25044 11076
rect 22848 11036 25044 11064
rect 21085 11027 21143 11033
rect 25038 11024 25044 11036
rect 25096 11024 25102 11076
rect 19613 10999 19671 11005
rect 19613 10965 19625 10999
rect 19659 10965 19671 10999
rect 19613 10959 19671 10965
rect 19794 10956 19800 11008
rect 19852 10996 19858 11008
rect 20073 10999 20131 11005
rect 20073 10996 20085 10999
rect 19852 10968 20085 10996
rect 19852 10956 19858 10968
rect 20073 10965 20085 10968
rect 20119 10965 20131 10999
rect 20073 10959 20131 10965
rect 20162 10956 20168 11008
rect 20220 10996 20226 11008
rect 24486 10996 24492 11008
rect 20220 10968 24492 10996
rect 20220 10956 20226 10968
rect 24486 10956 24492 10968
rect 24544 10956 24550 11008
rect 1104 10906 25852 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 25852 10906
rect 1104 10832 25852 10854
rect 9950 10752 9956 10804
rect 10008 10752 10014 10804
rect 12342 10752 12348 10804
rect 12400 10752 12406 10804
rect 12710 10752 12716 10804
rect 12768 10752 12774 10804
rect 14185 10795 14243 10801
rect 14185 10761 14197 10795
rect 14231 10792 14243 10795
rect 15933 10795 15991 10801
rect 14231 10764 15884 10792
rect 14231 10761 14243 10764
rect 14185 10755 14243 10761
rect 8481 10727 8539 10733
rect 8481 10724 8493 10727
rect 7852 10696 8493 10724
rect 7098 10412 7104 10464
rect 7156 10452 7162 10464
rect 7852 10461 7880 10696
rect 8481 10693 8493 10696
rect 8527 10693 8539 10727
rect 10410 10724 10416 10736
rect 9706 10696 10416 10724
rect 8481 10687 8539 10693
rect 10410 10684 10416 10696
rect 10468 10684 10474 10736
rect 12406 10696 12940 10724
rect 10870 10616 10876 10668
rect 10928 10656 10934 10668
rect 12406 10656 12434 10696
rect 10928 10628 12434 10656
rect 10928 10616 10934 10628
rect 12802 10616 12808 10668
rect 12860 10616 12866 10668
rect 8205 10591 8263 10597
rect 8205 10557 8217 10591
rect 8251 10557 8263 10591
rect 8205 10551 8263 10557
rect 11701 10591 11759 10597
rect 11701 10557 11713 10591
rect 11747 10588 11759 10591
rect 12710 10588 12716 10600
rect 11747 10560 12716 10588
rect 11747 10557 11759 10560
rect 11701 10551 11759 10557
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 7156 10424 7849 10452
rect 7156 10412 7162 10424
rect 7837 10421 7849 10424
rect 7883 10421 7895 10455
rect 8220 10452 8248 10551
rect 12710 10548 12716 10560
rect 12768 10548 12774 10600
rect 12912 10597 12940 10696
rect 13446 10684 13452 10736
rect 13504 10724 13510 10736
rect 15378 10724 15384 10736
rect 13504 10696 15384 10724
rect 13504 10684 13510 10696
rect 15378 10684 15384 10696
rect 15436 10684 15442 10736
rect 15856 10724 15884 10764
rect 15933 10761 15945 10795
rect 15979 10792 15991 10795
rect 17218 10792 17224 10804
rect 15979 10764 17224 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 17218 10752 17224 10764
rect 17276 10752 17282 10804
rect 17678 10792 17684 10804
rect 17328 10764 17684 10792
rect 17328 10724 17356 10764
rect 17678 10752 17684 10764
rect 17736 10752 17742 10804
rect 18414 10752 18420 10804
rect 18472 10792 18478 10804
rect 18874 10792 18880 10804
rect 18472 10764 18880 10792
rect 18472 10752 18478 10764
rect 18874 10752 18880 10764
rect 18932 10752 18938 10804
rect 19889 10795 19947 10801
rect 19889 10761 19901 10795
rect 19935 10792 19947 10795
rect 20162 10792 20168 10804
rect 19935 10764 20168 10792
rect 19935 10761 19947 10764
rect 19889 10755 19947 10761
rect 20162 10752 20168 10764
rect 20220 10752 20226 10804
rect 20717 10795 20775 10801
rect 20717 10761 20729 10795
rect 20763 10761 20775 10795
rect 20717 10755 20775 10761
rect 15856 10696 17356 10724
rect 17589 10727 17647 10733
rect 17589 10693 17601 10727
rect 17635 10724 17647 10727
rect 17770 10724 17776 10736
rect 17635 10696 17776 10724
rect 17635 10693 17647 10696
rect 17589 10687 17647 10693
rect 17770 10684 17776 10696
rect 17828 10684 17834 10736
rect 18322 10684 18328 10736
rect 18380 10724 18386 10736
rect 18598 10724 18604 10736
rect 18380 10696 18604 10724
rect 18380 10684 18386 10696
rect 18598 10684 18604 10696
rect 18656 10684 18662 10736
rect 20732 10724 20760 10755
rect 21266 10752 21272 10804
rect 21324 10792 21330 10804
rect 22002 10792 22008 10804
rect 21324 10764 22008 10792
rect 21324 10752 21330 10764
rect 22002 10752 22008 10764
rect 22060 10752 22066 10804
rect 23658 10792 23664 10804
rect 22572 10764 23664 10792
rect 22465 10727 22523 10733
rect 22465 10724 22477 10727
rect 19076 10696 20760 10724
rect 20824 10696 22477 10724
rect 16850 10656 16856 10668
rect 13004 10628 15332 10656
rect 12897 10591 12955 10597
rect 12897 10557 12909 10591
rect 12943 10557 12955 10591
rect 12897 10551 12955 10557
rect 10410 10480 10416 10532
rect 10468 10520 10474 10532
rect 11057 10523 11115 10529
rect 11057 10520 11069 10523
rect 10468 10492 11069 10520
rect 10468 10480 10474 10492
rect 11057 10489 11069 10492
rect 11103 10520 11115 10523
rect 11103 10492 11376 10520
rect 11103 10489 11115 10492
rect 11057 10483 11115 10489
rect 9030 10452 9036 10464
rect 8220 10424 9036 10452
rect 7837 10415 7895 10421
rect 9030 10412 9036 10424
rect 9088 10412 9094 10464
rect 11238 10412 11244 10464
rect 11296 10412 11302 10464
rect 11348 10452 11376 10492
rect 12250 10480 12256 10532
rect 12308 10520 12314 10532
rect 13004 10520 13032 10628
rect 13998 10548 14004 10600
rect 14056 10588 14062 10600
rect 14277 10591 14335 10597
rect 14277 10588 14289 10591
rect 14056 10560 14289 10588
rect 14056 10548 14062 10560
rect 14277 10557 14289 10560
rect 14323 10557 14335 10591
rect 14277 10551 14335 10557
rect 14458 10548 14464 10600
rect 14516 10548 14522 10600
rect 15304 10597 15332 10628
rect 16132 10628 16856 10656
rect 15289 10591 15347 10597
rect 15289 10557 15301 10591
rect 15335 10588 15347 10591
rect 16025 10591 16083 10597
rect 16025 10588 16037 10591
rect 15335 10560 16037 10588
rect 15335 10557 15347 10560
rect 15289 10551 15347 10557
rect 16025 10557 16037 10560
rect 16071 10588 16083 10591
rect 16132 10588 16160 10628
rect 16850 10616 16856 10628
rect 16908 10616 16914 10668
rect 17034 10616 17040 10668
rect 17092 10616 17098 10668
rect 18417 10659 18475 10665
rect 18417 10625 18429 10659
rect 18463 10656 18475 10659
rect 18782 10656 18788 10668
rect 18463 10628 18788 10656
rect 18463 10625 18475 10628
rect 18417 10619 18475 10625
rect 18782 10616 18788 10628
rect 18840 10616 18846 10668
rect 19076 10665 19104 10696
rect 19061 10659 19119 10665
rect 19061 10625 19073 10659
rect 19107 10625 19119 10659
rect 19061 10619 19119 10625
rect 19978 10616 19984 10668
rect 20036 10656 20042 10668
rect 20824 10656 20852 10696
rect 22465 10693 22477 10696
rect 22511 10693 22523 10727
rect 22465 10687 22523 10693
rect 20036 10628 20852 10656
rect 20036 10616 20042 10628
rect 21082 10616 21088 10668
rect 21140 10616 21146 10668
rect 22189 10659 22247 10665
rect 21376 10628 22094 10656
rect 16071 10560 16160 10588
rect 16209 10591 16267 10597
rect 16071 10557 16083 10560
rect 16025 10551 16083 10557
rect 16209 10557 16221 10591
rect 16255 10588 16267 10591
rect 16482 10588 16488 10600
rect 16255 10560 16488 10588
rect 16255 10557 16267 10560
rect 16209 10551 16267 10557
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 20070 10588 20076 10600
rect 16868 10560 20076 10588
rect 12308 10492 13032 10520
rect 12308 10480 12314 10492
rect 13630 10480 13636 10532
rect 13688 10520 13694 10532
rect 13817 10523 13875 10529
rect 13817 10520 13829 10523
rect 13688 10492 13829 10520
rect 13688 10480 13694 10492
rect 13817 10489 13829 10492
rect 13863 10489 13875 10523
rect 13817 10483 13875 10489
rect 15378 10480 15384 10532
rect 15436 10520 15442 10532
rect 16868 10529 16896 10560
rect 20070 10548 20076 10560
rect 20128 10548 20134 10600
rect 20165 10591 20223 10597
rect 20165 10557 20177 10591
rect 20211 10557 20223 10591
rect 20165 10551 20223 10557
rect 15565 10523 15623 10529
rect 15565 10520 15577 10523
rect 15436 10492 15577 10520
rect 15436 10480 15442 10492
rect 15565 10489 15577 10492
rect 15611 10489 15623 10523
rect 15565 10483 15623 10489
rect 16853 10523 16911 10529
rect 16853 10489 16865 10523
rect 16899 10489 16911 10523
rect 16853 10483 16911 10489
rect 18233 10523 18291 10529
rect 18233 10489 18245 10523
rect 18279 10520 18291 10523
rect 20180 10520 20208 10551
rect 20622 10548 20628 10600
rect 20680 10588 20686 10600
rect 21177 10591 21235 10597
rect 21177 10588 21189 10591
rect 20680 10560 21189 10588
rect 20680 10548 20686 10560
rect 21177 10557 21189 10560
rect 21223 10557 21235 10591
rect 21177 10551 21235 10557
rect 21266 10548 21272 10600
rect 21324 10548 21330 10600
rect 21376 10520 21404 10628
rect 22066 10588 22094 10628
rect 22189 10625 22201 10659
rect 22235 10656 22247 10659
rect 22572 10656 22600 10764
rect 23658 10752 23664 10764
rect 23716 10752 23722 10804
rect 23382 10684 23388 10736
rect 23440 10684 23446 10736
rect 22235 10628 22600 10656
rect 22235 10625 22247 10628
rect 22189 10619 22247 10625
rect 22646 10616 22652 10668
rect 22704 10656 22710 10668
rect 23109 10659 23167 10665
rect 23109 10656 23121 10659
rect 22704 10628 23121 10656
rect 22704 10616 22710 10628
rect 23109 10625 23121 10628
rect 23155 10625 23167 10659
rect 23109 10619 23167 10625
rect 22462 10588 22468 10600
rect 22066 10560 22468 10588
rect 22462 10548 22468 10560
rect 22520 10548 22526 10600
rect 22186 10520 22192 10532
rect 18279 10492 20116 10520
rect 20180 10492 21404 10520
rect 21468 10492 22192 10520
rect 18279 10489 18291 10492
rect 18233 10483 18291 10489
rect 11882 10452 11888 10464
rect 11348 10424 11888 10452
rect 11882 10412 11888 10424
rect 11940 10452 11946 10464
rect 13449 10455 13507 10461
rect 13449 10452 13461 10455
rect 11940 10424 13461 10452
rect 11940 10412 11946 10424
rect 13449 10421 13461 10424
rect 13495 10421 13507 10455
rect 13449 10415 13507 10421
rect 17678 10412 17684 10464
rect 17736 10412 17742 10464
rect 18046 10412 18052 10464
rect 18104 10452 18110 10464
rect 18877 10455 18935 10461
rect 18877 10452 18889 10455
rect 18104 10424 18889 10452
rect 18104 10412 18110 10424
rect 18877 10421 18889 10424
rect 18923 10421 18935 10455
rect 18877 10415 18935 10421
rect 19518 10412 19524 10464
rect 19576 10412 19582 10464
rect 20088 10452 20116 10492
rect 21468 10452 21496 10492
rect 22186 10480 22192 10492
rect 22244 10480 22250 10532
rect 24394 10480 24400 10532
rect 24452 10520 24458 10532
rect 24504 10520 24532 10642
rect 25133 10523 25191 10529
rect 25133 10520 25145 10523
rect 24452 10492 25145 10520
rect 24452 10480 24458 10492
rect 25133 10489 25145 10492
rect 25179 10489 25191 10523
rect 25133 10483 25191 10489
rect 20088 10424 21496 10452
rect 21818 10412 21824 10464
rect 21876 10452 21882 10464
rect 22005 10455 22063 10461
rect 22005 10452 22017 10455
rect 21876 10424 22017 10452
rect 21876 10412 21882 10424
rect 22005 10421 22017 10424
rect 22051 10421 22063 10455
rect 22005 10415 22063 10421
rect 22094 10412 22100 10464
rect 22152 10452 22158 10464
rect 22649 10455 22707 10461
rect 22649 10452 22661 10455
rect 22152 10424 22661 10452
rect 22152 10412 22158 10424
rect 22649 10421 22661 10424
rect 22695 10421 22707 10455
rect 22649 10415 22707 10421
rect 23382 10412 23388 10464
rect 23440 10452 23446 10464
rect 24857 10455 24915 10461
rect 24857 10452 24869 10455
rect 23440 10424 24869 10452
rect 23440 10412 23446 10424
rect 24857 10421 24869 10424
rect 24903 10421 24915 10455
rect 24857 10415 24915 10421
rect 1104 10362 25852 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 25852 10362
rect 1104 10288 25852 10310
rect 11054 10208 11060 10260
rect 11112 10208 11118 10260
rect 11606 10208 11612 10260
rect 11664 10208 11670 10260
rect 12066 10208 12072 10260
rect 12124 10248 12130 10260
rect 12805 10251 12863 10257
rect 12805 10248 12817 10251
rect 12124 10220 12817 10248
rect 12124 10208 12130 10220
rect 12805 10217 12817 10220
rect 12851 10217 12863 10251
rect 12805 10211 12863 10217
rect 13630 10208 13636 10260
rect 13688 10248 13694 10260
rect 13906 10248 13912 10260
rect 13688 10220 13912 10248
rect 13688 10208 13694 10220
rect 13906 10208 13912 10220
rect 13964 10208 13970 10260
rect 14090 10208 14096 10260
rect 14148 10248 14154 10260
rect 14553 10251 14611 10257
rect 14553 10248 14565 10251
rect 14148 10220 14565 10248
rect 14148 10208 14154 10220
rect 14553 10217 14565 10220
rect 14599 10217 14611 10251
rect 14553 10211 14611 10217
rect 15654 10208 15660 10260
rect 15712 10248 15718 10260
rect 19334 10248 19340 10260
rect 15712 10220 19340 10248
rect 15712 10208 15718 10220
rect 19334 10208 19340 10220
rect 19392 10208 19398 10260
rect 19518 10208 19524 10260
rect 19576 10248 19582 10260
rect 19576 10220 21864 10248
rect 19576 10208 19582 10220
rect 12526 10180 12532 10192
rect 11900 10152 12532 10180
rect 9122 10072 9128 10124
rect 9180 10112 9186 10124
rect 9585 10115 9643 10121
rect 9585 10112 9597 10115
rect 9180 10084 9597 10112
rect 9180 10072 9186 10084
rect 9585 10081 9597 10084
rect 9631 10081 9643 10115
rect 9585 10075 9643 10081
rect 9950 10072 9956 10124
rect 10008 10112 10014 10124
rect 11900 10112 11928 10152
rect 12526 10140 12532 10152
rect 12584 10140 12590 10192
rect 14826 10140 14832 10192
rect 14884 10180 14890 10192
rect 17586 10180 17592 10192
rect 14884 10152 17592 10180
rect 14884 10140 14890 10152
rect 17586 10140 17592 10152
rect 17644 10140 17650 10192
rect 17957 10183 18015 10189
rect 17957 10149 17969 10183
rect 18003 10180 18015 10183
rect 18322 10180 18328 10192
rect 18003 10152 18328 10180
rect 18003 10149 18015 10152
rect 17957 10143 18015 10149
rect 18322 10140 18328 10152
rect 18380 10140 18386 10192
rect 20346 10180 20352 10192
rect 18524 10152 20352 10180
rect 10008 10084 11928 10112
rect 10008 10072 10014 10084
rect 11974 10072 11980 10124
rect 12032 10112 12038 10124
rect 12161 10115 12219 10121
rect 12161 10112 12173 10115
rect 12032 10084 12173 10112
rect 12032 10072 12038 10084
rect 12161 10081 12173 10084
rect 12207 10081 12219 10115
rect 12161 10075 12219 10081
rect 13449 10115 13507 10121
rect 13449 10081 13461 10115
rect 13495 10112 13507 10115
rect 13538 10112 13544 10124
rect 13495 10084 13544 10112
rect 13495 10081 13507 10084
rect 13449 10075 13507 10081
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 13909 10115 13967 10121
rect 13909 10081 13921 10115
rect 13955 10112 13967 10115
rect 15010 10112 15016 10124
rect 13955 10084 15016 10112
rect 13955 10081 13967 10084
rect 13909 10075 13967 10081
rect 9030 10004 9036 10056
rect 9088 10044 9094 10056
rect 9309 10047 9367 10053
rect 9309 10044 9321 10047
rect 9088 10016 9321 10044
rect 9088 10004 9094 10016
rect 9309 10013 9321 10016
rect 9355 10013 9367 10047
rect 9309 10007 9367 10013
rect 12710 10004 12716 10056
rect 12768 10044 12774 10056
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 12768 10016 13185 10044
rect 12768 10004 12774 10016
rect 13173 10013 13185 10016
rect 13219 10013 13231 10047
rect 13173 10007 13231 10013
rect 10318 9936 10324 9988
rect 10376 9936 10382 9988
rect 11977 9979 12035 9985
rect 11977 9945 11989 9979
rect 12023 9976 12035 9979
rect 12342 9976 12348 9988
rect 12023 9948 12348 9976
rect 12023 9945 12035 9948
rect 11977 9939 12035 9945
rect 12342 9936 12348 9948
rect 12400 9936 12406 9988
rect 12526 9936 12532 9988
rect 12584 9976 12590 9988
rect 13924 9976 13952 10075
rect 15010 10072 15016 10084
rect 15068 10072 15074 10124
rect 15105 10115 15163 10121
rect 15105 10081 15117 10115
rect 15151 10112 15163 10115
rect 15838 10112 15844 10124
rect 15151 10084 15844 10112
rect 15151 10081 15163 10084
rect 15105 10075 15163 10081
rect 14277 10047 14335 10053
rect 14277 10013 14289 10047
rect 14323 10044 14335 10047
rect 14550 10044 14556 10056
rect 14323 10016 14556 10044
rect 14323 10013 14335 10016
rect 14277 10007 14335 10013
rect 14550 10004 14556 10016
rect 14608 10044 14614 10056
rect 15120 10044 15148 10075
rect 15838 10072 15844 10084
rect 15896 10072 15902 10124
rect 18524 10112 18552 10152
rect 20346 10140 20352 10152
rect 20404 10140 20410 10192
rect 21836 10180 21864 10220
rect 22002 10208 22008 10260
rect 22060 10248 22066 10260
rect 22281 10251 22339 10257
rect 22281 10248 22293 10251
rect 22060 10220 22293 10248
rect 22060 10208 22066 10220
rect 22281 10217 22293 10220
rect 22327 10217 22339 10251
rect 22281 10211 22339 10217
rect 24578 10208 24584 10260
rect 24636 10208 24642 10260
rect 24486 10180 24492 10192
rect 21836 10152 24492 10180
rect 24486 10140 24492 10152
rect 24544 10140 24550 10192
rect 16132 10084 18552 10112
rect 18601 10115 18659 10121
rect 14608 10016 15148 10044
rect 14608 10004 14614 10016
rect 12584 9948 13952 9976
rect 14921 9979 14979 9985
rect 12584 9936 12590 9948
rect 14921 9945 14933 9979
rect 14967 9976 14979 9979
rect 15654 9976 15660 9988
rect 14967 9948 15660 9976
rect 14967 9945 14979 9948
rect 14921 9939 14979 9945
rect 15654 9936 15660 9948
rect 15712 9936 15718 9988
rect 7098 9868 7104 9920
rect 7156 9908 7162 9920
rect 11882 9908 11888 9920
rect 7156 9880 11888 9908
rect 7156 9868 7162 9880
rect 11882 9868 11888 9880
rect 11940 9868 11946 9920
rect 12069 9911 12127 9917
rect 12069 9877 12081 9911
rect 12115 9908 12127 9911
rect 12802 9908 12808 9920
rect 12115 9880 12808 9908
rect 12115 9877 12127 9880
rect 12069 9871 12127 9877
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 13265 9911 13323 9917
rect 13265 9877 13277 9911
rect 13311 9908 13323 9911
rect 14734 9908 14740 9920
rect 13311 9880 14740 9908
rect 13311 9877 13323 9880
rect 13265 9871 13323 9877
rect 14734 9868 14740 9880
rect 14792 9908 14798 9920
rect 15470 9908 15476 9920
rect 14792 9880 15476 9908
rect 14792 9868 14798 9880
rect 15470 9868 15476 9880
rect 15528 9868 15534 9920
rect 15838 9868 15844 9920
rect 15896 9868 15902 9920
rect 16132 9917 16160 10084
rect 18601 10081 18613 10115
rect 18647 10112 18659 10115
rect 19242 10112 19248 10124
rect 18647 10084 19248 10112
rect 18647 10081 18659 10084
rect 18601 10075 18659 10081
rect 19242 10072 19248 10084
rect 19300 10072 19306 10124
rect 19334 10072 19340 10124
rect 19392 10112 19398 10124
rect 20254 10112 20260 10124
rect 19392 10084 20260 10112
rect 19392 10072 19398 10084
rect 20254 10072 20260 10084
rect 20312 10072 20318 10124
rect 22002 10072 22008 10124
rect 22060 10112 22066 10124
rect 23293 10115 23351 10121
rect 23293 10112 23305 10115
rect 22060 10084 23305 10112
rect 22060 10072 22066 10084
rect 23293 10081 23305 10084
rect 23339 10081 23351 10115
rect 23293 10075 23351 10081
rect 23382 10072 23388 10124
rect 23440 10072 23446 10124
rect 16942 10004 16948 10056
rect 17000 10044 17006 10056
rect 20533 10047 20591 10053
rect 20533 10044 20545 10047
rect 17000 10016 20545 10044
rect 17000 10004 17006 10016
rect 20533 10013 20545 10016
rect 20579 10013 20591 10047
rect 22094 10044 22100 10056
rect 21942 10016 22100 10044
rect 20533 10007 20591 10013
rect 22094 10004 22100 10016
rect 22152 10004 22158 10056
rect 22738 10004 22744 10056
rect 22796 10044 22802 10056
rect 24765 10047 24823 10053
rect 24765 10044 24777 10047
rect 22796 10016 24777 10044
rect 22796 10004 22802 10016
rect 24765 10013 24777 10016
rect 24811 10013 24823 10047
rect 24765 10007 24823 10013
rect 16853 9979 16911 9985
rect 16853 9945 16865 9979
rect 16899 9976 16911 9979
rect 19058 9976 19064 9988
rect 16899 9948 19064 9976
rect 16899 9945 16911 9948
rect 16853 9939 16911 9945
rect 19058 9936 19064 9948
rect 19116 9936 19122 9988
rect 19521 9979 19579 9985
rect 19521 9945 19533 9979
rect 19567 9976 19579 9979
rect 20438 9976 20444 9988
rect 19567 9948 20444 9976
rect 19567 9945 19579 9948
rect 19521 9939 19579 9945
rect 20438 9936 20444 9948
rect 20496 9936 20502 9988
rect 20714 9936 20720 9988
rect 20772 9976 20778 9988
rect 20809 9979 20867 9985
rect 20809 9976 20821 9979
rect 20772 9948 20821 9976
rect 20772 9936 20778 9948
rect 20809 9945 20821 9948
rect 20855 9976 20867 9979
rect 20898 9976 20904 9988
rect 20855 9948 20904 9976
rect 20855 9945 20867 9948
rect 20809 9939 20867 9945
rect 20898 9936 20904 9948
rect 20956 9936 20962 9988
rect 22204 9948 22876 9976
rect 16025 9911 16083 9917
rect 16025 9877 16037 9911
rect 16071 9908 16083 9911
rect 16117 9911 16175 9917
rect 16117 9908 16129 9911
rect 16071 9880 16129 9908
rect 16071 9877 16083 9880
rect 16025 9871 16083 9877
rect 16117 9877 16129 9880
rect 16163 9877 16175 9911
rect 16117 9871 16175 9877
rect 16758 9868 16764 9920
rect 16816 9908 16822 9920
rect 16945 9911 17003 9917
rect 16945 9908 16957 9911
rect 16816 9880 16957 9908
rect 16816 9868 16822 9880
rect 16945 9877 16957 9880
rect 16991 9877 17003 9911
rect 16945 9871 17003 9877
rect 17586 9868 17592 9920
rect 17644 9908 17650 9920
rect 18325 9911 18383 9917
rect 18325 9908 18337 9911
rect 17644 9880 18337 9908
rect 17644 9868 17650 9880
rect 18325 9877 18337 9880
rect 18371 9877 18383 9911
rect 18325 9871 18383 9877
rect 18417 9911 18475 9917
rect 18417 9877 18429 9911
rect 18463 9908 18475 9911
rect 18506 9908 18512 9920
rect 18463 9880 18512 9908
rect 18463 9877 18475 9880
rect 18417 9871 18475 9877
rect 18506 9868 18512 9880
rect 18564 9908 18570 9920
rect 18969 9911 19027 9917
rect 18969 9908 18981 9911
rect 18564 9880 18981 9908
rect 18564 9868 18570 9880
rect 18969 9877 18981 9880
rect 19015 9877 19027 9911
rect 18969 9871 19027 9877
rect 19613 9911 19671 9917
rect 19613 9877 19625 9911
rect 19659 9908 19671 9911
rect 19702 9908 19708 9920
rect 19659 9880 19708 9908
rect 19659 9877 19671 9880
rect 19613 9871 19671 9877
rect 19702 9868 19708 9880
rect 19760 9868 19766 9920
rect 19794 9868 19800 9920
rect 19852 9908 19858 9920
rect 19981 9911 20039 9917
rect 19981 9908 19993 9911
rect 19852 9880 19993 9908
rect 19852 9868 19858 9880
rect 19981 9877 19993 9880
rect 20027 9877 20039 9911
rect 19981 9871 20039 9877
rect 20162 9868 20168 9920
rect 20220 9868 20226 9920
rect 20622 9868 20628 9920
rect 20680 9908 20686 9920
rect 22204 9908 22232 9948
rect 22848 9917 22876 9948
rect 20680 9880 22232 9908
rect 22833 9911 22891 9917
rect 20680 9868 20686 9880
rect 22833 9877 22845 9911
rect 22879 9877 22891 9911
rect 22833 9871 22891 9877
rect 23201 9911 23259 9917
rect 23201 9877 23213 9911
rect 23247 9908 23259 9911
rect 24670 9908 24676 9920
rect 23247 9880 24676 9908
rect 23247 9877 23259 9880
rect 23201 9871 23259 9877
rect 24670 9868 24676 9880
rect 24728 9868 24734 9920
rect 1104 9818 25852 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 25852 9818
rect 1104 9744 25852 9766
rect 10962 9664 10968 9716
rect 11020 9704 11026 9716
rect 11333 9707 11391 9713
rect 11333 9704 11345 9707
rect 11020 9676 11345 9704
rect 11020 9664 11026 9676
rect 11333 9673 11345 9676
rect 11379 9704 11391 9707
rect 11379 9676 12434 9704
rect 11379 9673 11391 9676
rect 11333 9667 11391 9673
rect 12406 9648 12434 9676
rect 12710 9664 12716 9716
rect 12768 9704 12774 9716
rect 14550 9704 14556 9716
rect 12768 9676 14556 9704
rect 12768 9664 12774 9676
rect 14550 9664 14556 9676
rect 14608 9664 14614 9716
rect 15838 9664 15844 9716
rect 15896 9704 15902 9716
rect 20162 9704 20168 9716
rect 15896 9676 20168 9704
rect 15896 9664 15902 9676
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 20254 9664 20260 9716
rect 20312 9704 20318 9716
rect 20312 9676 21036 9704
rect 20312 9664 20318 9676
rect 10502 9596 10508 9648
rect 10560 9636 10566 9648
rect 12250 9636 12256 9648
rect 10560 9608 12256 9636
rect 10560 9596 10566 9608
rect 12250 9596 12256 9608
rect 12308 9596 12314 9648
rect 12406 9608 12440 9648
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 15473 9639 15531 9645
rect 15473 9605 15485 9639
rect 15519 9636 15531 9639
rect 15519 9608 16436 9636
rect 15519 9605 15531 9608
rect 15473 9599 15531 9605
rect 11698 9528 11704 9580
rect 11756 9528 11762 9580
rect 14277 9571 14335 9577
rect 14277 9537 14289 9571
rect 14323 9568 14335 9571
rect 15378 9568 15384 9580
rect 14323 9540 15384 9568
rect 14323 9537 14335 9540
rect 14277 9531 14335 9537
rect 15378 9528 15384 9540
rect 15436 9528 15442 9580
rect 12342 9460 12348 9512
rect 12400 9500 12406 9512
rect 12400 9472 13952 9500
rect 12400 9460 12406 9472
rect 13449 9435 13507 9441
rect 13449 9401 13461 9435
rect 13495 9432 13507 9435
rect 13814 9432 13820 9444
rect 13495 9404 13820 9432
rect 13495 9401 13507 9404
rect 13449 9395 13507 9401
rect 13814 9392 13820 9404
rect 13872 9392 13878 9444
rect 13924 9441 13952 9472
rect 14090 9460 14096 9512
rect 14148 9500 14154 9512
rect 14369 9503 14427 9509
rect 14369 9500 14381 9503
rect 14148 9472 14381 9500
rect 14148 9460 14154 9472
rect 14369 9469 14381 9472
rect 14415 9469 14427 9503
rect 14369 9463 14427 9469
rect 13909 9435 13967 9441
rect 13909 9401 13921 9435
rect 13955 9401 13967 9435
rect 14384 9432 14412 9463
rect 14550 9460 14556 9512
rect 14608 9460 14614 9512
rect 15562 9460 15568 9512
rect 15620 9460 15626 9512
rect 15746 9460 15752 9512
rect 15804 9460 15810 9512
rect 14642 9432 14648 9444
rect 14384 9404 14648 9432
rect 13909 9395 13967 9401
rect 14642 9392 14648 9404
rect 14700 9432 14706 9444
rect 16408 9441 16436 9608
rect 17494 9596 17500 9648
rect 17552 9636 17558 9648
rect 18046 9636 18052 9648
rect 17552 9608 18052 9636
rect 17552 9596 17558 9608
rect 18046 9596 18052 9608
rect 18104 9596 18110 9648
rect 19058 9596 19064 9648
rect 19116 9636 19122 9648
rect 20622 9636 20628 9648
rect 19116 9608 20628 9636
rect 19116 9596 19122 9608
rect 20622 9596 20628 9608
rect 20680 9596 20686 9648
rect 20254 9528 20260 9580
rect 20312 9528 20318 9580
rect 21008 9568 21036 9676
rect 21082 9664 21088 9716
rect 21140 9704 21146 9716
rect 22005 9707 22063 9713
rect 22005 9704 22017 9707
rect 21140 9676 22017 9704
rect 21140 9664 21146 9676
rect 22005 9673 22017 9676
rect 22051 9673 22063 9707
rect 22005 9667 22063 9673
rect 23308 9676 24256 9704
rect 21450 9596 21456 9648
rect 21508 9636 21514 9648
rect 23308 9636 23336 9676
rect 21508 9608 23336 9636
rect 21508 9596 21514 9608
rect 21008 9540 21956 9568
rect 16942 9460 16948 9512
rect 17000 9500 17006 9512
rect 17313 9503 17371 9509
rect 17313 9500 17325 9503
rect 17000 9472 17325 9500
rect 17000 9460 17006 9472
rect 17313 9469 17325 9472
rect 17359 9469 17371 9503
rect 18874 9500 18880 9512
rect 17313 9463 17371 9469
rect 17420 9472 18880 9500
rect 16117 9435 16175 9441
rect 16117 9432 16129 9435
rect 14700 9404 16129 9432
rect 14700 9392 14706 9404
rect 16117 9401 16129 9404
rect 16163 9401 16175 9435
rect 16117 9395 16175 9401
rect 16393 9435 16451 9441
rect 16393 9401 16405 9435
rect 16439 9432 16451 9435
rect 17420 9432 17448 9472
rect 18874 9460 18880 9472
rect 18932 9500 18938 9512
rect 21082 9500 21088 9512
rect 18932 9472 21088 9500
rect 18932 9460 18938 9472
rect 21082 9460 21088 9472
rect 21140 9460 21146 9512
rect 21174 9460 21180 9512
rect 21232 9460 21238 9512
rect 16439 9404 17448 9432
rect 21928 9432 21956 9540
rect 22094 9528 22100 9580
rect 22152 9568 22158 9580
rect 22646 9568 22652 9580
rect 22152 9540 22652 9568
rect 22152 9528 22158 9540
rect 22646 9528 22652 9540
rect 22704 9528 22710 9580
rect 24026 9528 24032 9580
rect 24084 9528 24090 9580
rect 24228 9568 24256 9676
rect 25041 9571 25099 9577
rect 25041 9568 25053 9571
rect 24228 9540 25053 9568
rect 25041 9537 25053 9540
rect 25087 9537 25099 9571
rect 25041 9531 25099 9537
rect 22925 9503 22983 9509
rect 22925 9469 22937 9503
rect 22971 9500 22983 9503
rect 23382 9500 23388 9512
rect 22971 9472 23388 9500
rect 22971 9469 22983 9472
rect 22925 9463 22983 9469
rect 23382 9460 23388 9472
rect 23440 9460 23446 9512
rect 24044 9500 24072 9528
rect 24394 9500 24400 9512
rect 24044 9472 24400 9500
rect 24394 9460 24400 9472
rect 24452 9500 24458 9512
rect 25317 9503 25375 9509
rect 25317 9500 25329 9503
rect 24452 9472 25329 9500
rect 24452 9460 24458 9472
rect 25317 9469 25329 9472
rect 25363 9469 25375 9503
rect 25317 9463 25375 9469
rect 22646 9432 22652 9444
rect 21928 9404 22652 9432
rect 16439 9401 16451 9404
rect 16393 9395 16451 9401
rect 22646 9392 22652 9404
rect 22704 9392 22710 9444
rect 11964 9367 12022 9373
rect 11964 9333 11976 9367
rect 12010 9364 12022 9367
rect 12342 9364 12348 9376
rect 12010 9336 12348 9364
rect 12010 9333 12022 9336
rect 11964 9327 12022 9333
rect 12342 9324 12348 9336
rect 12400 9324 12406 9376
rect 13722 9324 13728 9376
rect 13780 9364 13786 9376
rect 15105 9367 15163 9373
rect 15105 9364 15117 9367
rect 13780 9336 15117 9364
rect 13780 9324 13786 9336
rect 15105 9333 15117 9336
rect 15151 9333 15163 9367
rect 15105 9327 15163 9333
rect 15654 9324 15660 9376
rect 15712 9364 15718 9376
rect 15930 9364 15936 9376
rect 15712 9336 15936 9364
rect 15712 9324 15718 9336
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 16850 9324 16856 9376
rect 16908 9324 16914 9376
rect 17037 9367 17095 9373
rect 17037 9333 17049 9367
rect 17083 9364 17095 9367
rect 17126 9364 17132 9376
rect 17083 9336 17132 9364
rect 17083 9333 17095 9336
rect 17037 9327 17095 9333
rect 17126 9324 17132 9336
rect 17184 9324 17190 9376
rect 17586 9373 17592 9376
rect 17576 9367 17592 9373
rect 17576 9333 17588 9367
rect 17576 9327 17592 9333
rect 17586 9324 17592 9327
rect 17644 9324 17650 9376
rect 17954 9324 17960 9376
rect 18012 9364 18018 9376
rect 18874 9364 18880 9376
rect 18012 9336 18880 9364
rect 18012 9324 18018 9336
rect 18874 9324 18880 9336
rect 18932 9364 18938 9376
rect 19061 9367 19119 9373
rect 19061 9364 19073 9367
rect 18932 9336 19073 9364
rect 18932 9324 18938 9336
rect 19061 9333 19073 9336
rect 19107 9333 19119 9367
rect 19061 9327 19119 9333
rect 19429 9367 19487 9373
rect 19429 9333 19441 9367
rect 19475 9364 19487 9367
rect 19794 9364 19800 9376
rect 19475 9336 19800 9364
rect 19475 9333 19487 9336
rect 19429 9327 19487 9333
rect 19794 9324 19800 9336
rect 19852 9324 19858 9376
rect 22462 9324 22468 9376
rect 22520 9364 22526 9376
rect 24397 9367 24455 9373
rect 24397 9364 24409 9367
rect 22520 9336 24409 9364
rect 22520 9324 22526 9336
rect 24397 9333 24409 9336
rect 24443 9333 24455 9367
rect 24397 9327 24455 9333
rect 24854 9324 24860 9376
rect 24912 9324 24918 9376
rect 1104 9274 25852 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 25852 9274
rect 1104 9200 25852 9222
rect 10962 9120 10968 9172
rect 11020 9160 11026 9172
rect 11149 9163 11207 9169
rect 11149 9160 11161 9163
rect 11020 9132 11161 9160
rect 11020 9120 11026 9132
rect 11149 9129 11161 9132
rect 11195 9129 11207 9163
rect 11149 9123 11207 9129
rect 11882 9120 11888 9172
rect 11940 9160 11946 9172
rect 12621 9163 12679 9169
rect 12621 9160 12633 9163
rect 11940 9132 12633 9160
rect 11940 9120 11946 9132
rect 12621 9129 12633 9132
rect 12667 9129 12679 9163
rect 12621 9123 12679 9129
rect 12802 9120 12808 9172
rect 12860 9160 12866 9172
rect 14277 9163 14335 9169
rect 14277 9160 14289 9163
rect 12860 9132 14289 9160
rect 12860 9120 12866 9132
rect 14277 9129 14289 9132
rect 14323 9129 14335 9163
rect 14277 9123 14335 9129
rect 14642 9120 14648 9172
rect 14700 9160 14706 9172
rect 15102 9160 15108 9172
rect 14700 9132 15108 9160
rect 14700 9120 14706 9132
rect 15102 9120 15108 9132
rect 15160 9160 15166 9172
rect 15286 9160 15292 9172
rect 15160 9132 15292 9160
rect 15160 9120 15166 9132
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 17402 9160 17408 9172
rect 15580 9132 17408 9160
rect 15580 9104 15608 9132
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 17494 9120 17500 9172
rect 17552 9160 17558 9172
rect 18233 9163 18291 9169
rect 18233 9160 18245 9163
rect 17552 9132 18245 9160
rect 17552 9120 17558 9132
rect 18233 9129 18245 9132
rect 18279 9160 18291 9163
rect 20070 9160 20076 9172
rect 18279 9132 20076 9160
rect 18279 9129 18291 9132
rect 18233 9123 18291 9129
rect 20070 9120 20076 9132
rect 20128 9120 20134 9172
rect 20898 9120 20904 9172
rect 20956 9160 20962 9172
rect 21361 9163 21419 9169
rect 21361 9160 21373 9163
rect 20956 9132 21373 9160
rect 20956 9120 20962 9132
rect 21361 9129 21373 9132
rect 21407 9129 21419 9163
rect 21361 9123 21419 9129
rect 12989 9095 13047 9101
rect 12989 9061 13001 9095
rect 13035 9092 13047 9095
rect 13354 9092 13360 9104
rect 13035 9064 13360 9092
rect 13035 9061 13047 9064
rect 12989 9055 13047 9061
rect 13354 9052 13360 9064
rect 13412 9052 13418 9104
rect 15473 9095 15531 9101
rect 15473 9092 15485 9095
rect 13464 9064 15485 9092
rect 9125 9027 9183 9033
rect 9125 8993 9137 9027
rect 9171 9024 9183 9027
rect 11698 9024 11704 9036
rect 9171 8996 11704 9024
rect 9171 8993 9183 8996
rect 9125 8987 9183 8993
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 11882 8984 11888 9036
rect 11940 9024 11946 9036
rect 13464 9024 13492 9064
rect 15473 9061 15485 9064
rect 15519 9092 15531 9095
rect 15562 9092 15568 9104
rect 15519 9064 15568 9092
rect 15519 9061 15531 9064
rect 15473 9055 15531 9061
rect 15562 9052 15568 9064
rect 15620 9052 15626 9104
rect 15746 9052 15752 9104
rect 15804 9092 15810 9104
rect 19610 9092 19616 9104
rect 15804 9064 17632 9092
rect 15804 9052 15810 9064
rect 11940 8996 13492 9024
rect 11940 8984 11946 8996
rect 13538 8984 13544 9036
rect 13596 8984 13602 9036
rect 14550 8984 14556 9036
rect 14608 9024 14614 9036
rect 14829 9027 14887 9033
rect 14829 9024 14841 9027
rect 14608 8996 14841 9024
rect 14608 8984 14614 8996
rect 14829 8993 14841 8996
rect 14875 8993 14887 9027
rect 14829 8987 14887 8993
rect 16482 8984 16488 9036
rect 16540 8984 16546 9036
rect 17604 9024 17632 9064
rect 17880 9064 19616 9092
rect 17773 9027 17831 9033
rect 17773 9024 17785 9027
rect 17604 8996 17785 9024
rect 17773 8993 17785 8996
rect 17819 8993 17831 9027
rect 17773 8987 17831 8993
rect 2774 8916 2780 8968
rect 2832 8956 2838 8968
rect 4798 8956 4804 8968
rect 2832 8928 4804 8956
rect 2832 8916 2838 8928
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 10962 8956 10968 8968
rect 10534 8928 10968 8956
rect 10962 8916 10968 8928
rect 11020 8956 11026 8968
rect 12434 8956 12440 8968
rect 11020 8928 12440 8956
rect 11020 8916 11026 8928
rect 12434 8916 12440 8928
rect 12492 8916 12498 8968
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8956 13507 8959
rect 15838 8956 15844 8968
rect 13495 8928 15844 8956
rect 13495 8925 13507 8928
rect 13449 8919 13507 8925
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 15930 8916 15936 8968
rect 15988 8956 15994 8968
rect 16393 8959 16451 8965
rect 16393 8956 16405 8959
rect 15988 8928 16405 8956
rect 15988 8916 15994 8928
rect 16393 8925 16405 8928
rect 16439 8925 16451 8959
rect 16393 8919 16451 8925
rect 17126 8916 17132 8968
rect 17184 8956 17190 8968
rect 17589 8959 17647 8965
rect 17589 8956 17601 8959
rect 17184 8928 17601 8956
rect 17184 8916 17190 8928
rect 17589 8925 17601 8928
rect 17635 8956 17647 8959
rect 17880 8956 17908 9064
rect 19610 9052 19616 9064
rect 19668 9052 19674 9104
rect 24854 9092 24860 9104
rect 20916 9064 24860 9092
rect 17954 8984 17960 9036
rect 18012 9024 18018 9036
rect 20916 9024 20944 9064
rect 24854 9052 24860 9064
rect 24912 9052 24918 9104
rect 18012 8996 18736 9024
rect 18012 8984 18018 8996
rect 17635 8928 17908 8956
rect 18708 8956 18736 8996
rect 19306 8996 20944 9024
rect 21008 8996 22416 9024
rect 19306 8956 19334 8996
rect 18708 8928 19334 8956
rect 17635 8925 17647 8928
rect 17589 8919 17647 8925
rect 19610 8916 19616 8968
rect 19668 8916 19674 8968
rect 21008 8942 21036 8996
rect 22005 8959 22063 8965
rect 22005 8956 22017 8959
rect 21192 8928 22017 8956
rect 9401 8891 9459 8897
rect 9401 8857 9413 8891
rect 9447 8888 9459 8891
rect 9674 8888 9680 8900
rect 9447 8860 9680 8888
rect 9447 8857 9459 8860
rect 9401 8851 9459 8857
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 13357 8891 13415 8897
rect 13357 8857 13369 8891
rect 13403 8888 13415 8891
rect 13403 8860 17172 8888
rect 13403 8857 13415 8860
rect 13357 8851 13415 8857
rect 2406 8780 2412 8832
rect 2464 8820 2470 8832
rect 8570 8820 8576 8832
rect 2464 8792 8576 8820
rect 2464 8780 2470 8792
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 10873 8823 10931 8829
rect 10873 8789 10885 8823
rect 10919 8820 10931 8823
rect 10962 8820 10968 8832
rect 10919 8792 10968 8820
rect 10919 8789 10931 8792
rect 10873 8783 10931 8789
rect 10962 8780 10968 8792
rect 11020 8780 11026 8832
rect 14642 8780 14648 8832
rect 14700 8780 14706 8832
rect 14737 8823 14795 8829
rect 14737 8789 14749 8823
rect 14783 8820 14795 8823
rect 14826 8820 14832 8832
rect 14783 8792 14832 8820
rect 14783 8789 14795 8792
rect 14737 8783 14795 8789
rect 14826 8780 14832 8792
rect 14884 8820 14890 8832
rect 15010 8820 15016 8832
rect 14884 8792 15016 8820
rect 14884 8780 14890 8792
rect 15010 8780 15016 8792
rect 15068 8780 15074 8832
rect 15378 8780 15384 8832
rect 15436 8780 15442 8832
rect 15654 8780 15660 8832
rect 15712 8820 15718 8832
rect 15933 8823 15991 8829
rect 15933 8820 15945 8823
rect 15712 8792 15945 8820
rect 15712 8780 15718 8792
rect 15933 8789 15945 8792
rect 15979 8789 15991 8823
rect 15933 8783 15991 8789
rect 16301 8823 16359 8829
rect 16301 8789 16313 8823
rect 16347 8820 16359 8823
rect 16850 8820 16856 8832
rect 16347 8792 16856 8820
rect 16347 8789 16359 8792
rect 16301 8783 16359 8789
rect 16850 8780 16856 8792
rect 16908 8780 16914 8832
rect 17144 8829 17172 8860
rect 17494 8848 17500 8900
rect 17552 8848 17558 8900
rect 18690 8848 18696 8900
rect 18748 8848 18754 8900
rect 18877 8891 18935 8897
rect 18877 8857 18889 8891
rect 18923 8888 18935 8891
rect 19334 8888 19340 8900
rect 18923 8860 19340 8888
rect 18923 8857 18935 8860
rect 18877 8851 18935 8857
rect 19334 8848 19340 8860
rect 19392 8848 19398 8900
rect 19794 8848 19800 8900
rect 19852 8888 19858 8900
rect 19889 8891 19947 8897
rect 19889 8888 19901 8891
rect 19852 8860 19901 8888
rect 19852 8848 19858 8860
rect 19889 8857 19901 8860
rect 19935 8857 19947 8891
rect 19889 8851 19947 8857
rect 17129 8823 17187 8829
rect 17129 8789 17141 8823
rect 17175 8789 17187 8823
rect 17129 8783 17187 8789
rect 17770 8780 17776 8832
rect 17828 8820 17834 8832
rect 21192 8820 21220 8928
rect 22005 8925 22017 8928
rect 22051 8925 22063 8959
rect 22005 8919 22063 8925
rect 17828 8792 21220 8820
rect 17828 8780 17834 8792
rect 21450 8780 21456 8832
rect 21508 8820 21514 8832
rect 22388 8829 22416 8996
rect 22646 8916 22652 8968
rect 22704 8916 22710 8968
rect 24210 8916 24216 8968
rect 24268 8956 24274 8968
rect 24765 8959 24823 8965
rect 24765 8956 24777 8959
rect 24268 8928 24777 8956
rect 24268 8916 24274 8928
rect 24765 8925 24777 8928
rect 24811 8925 24823 8959
rect 24765 8919 24823 8925
rect 23845 8891 23903 8897
rect 23845 8857 23857 8891
rect 23891 8888 23903 8891
rect 24946 8888 24952 8900
rect 23891 8860 24952 8888
rect 23891 8857 23903 8860
rect 23845 8851 23903 8857
rect 24946 8848 24952 8860
rect 25004 8848 25010 8900
rect 21821 8823 21879 8829
rect 21821 8820 21833 8823
rect 21508 8792 21833 8820
rect 21508 8780 21514 8792
rect 21821 8789 21833 8792
rect 21867 8789 21879 8823
rect 21821 8783 21879 8789
rect 22373 8823 22431 8829
rect 22373 8789 22385 8823
rect 22419 8820 22431 8823
rect 24026 8820 24032 8832
rect 22419 8792 24032 8820
rect 22419 8789 22431 8792
rect 22373 8783 22431 8789
rect 24026 8780 24032 8792
rect 24084 8780 24090 8832
rect 24578 8780 24584 8832
rect 24636 8780 24642 8832
rect 1104 8730 25852 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 25852 8730
rect 1104 8656 25852 8678
rect 9674 8576 9680 8628
rect 9732 8616 9738 8628
rect 9950 8616 9956 8628
rect 9732 8588 9956 8616
rect 9732 8576 9738 8588
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 12618 8576 12624 8628
rect 12676 8616 12682 8628
rect 12805 8619 12863 8625
rect 12805 8616 12817 8619
rect 12676 8588 12817 8616
rect 12676 8576 12682 8588
rect 12805 8585 12817 8588
rect 12851 8616 12863 8619
rect 14461 8619 14519 8625
rect 12851 8588 13952 8616
rect 12851 8585 12863 8588
rect 12805 8579 12863 8585
rect 12526 8508 12532 8560
rect 12584 8548 12590 8560
rect 13722 8548 13728 8560
rect 12584 8520 13728 8548
rect 12584 8508 12590 8520
rect 13722 8508 13728 8520
rect 13780 8508 13786 8560
rect 13924 8557 13952 8588
rect 14461 8585 14473 8619
rect 14507 8616 14519 8619
rect 14550 8616 14556 8628
rect 14507 8588 14556 8616
rect 14507 8585 14519 8588
rect 14461 8579 14519 8585
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 15059 8619 15117 8625
rect 15059 8585 15071 8619
rect 15105 8616 15117 8619
rect 15105 8588 23980 8616
rect 15105 8585 15117 8588
rect 15059 8579 15117 8585
rect 13909 8551 13967 8557
rect 13909 8517 13921 8551
rect 13955 8517 13967 8551
rect 13909 8511 13967 8517
rect 14090 8508 14096 8560
rect 14148 8508 14154 8560
rect 16850 8508 16856 8560
rect 16908 8548 16914 8560
rect 23658 8548 23664 8560
rect 16908 8520 19196 8548
rect 16908 8508 16914 8520
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 14829 8483 14887 8489
rect 14829 8480 14841 8483
rect 14700 8452 14841 8480
rect 14700 8440 14706 8452
rect 14829 8449 14841 8452
rect 14875 8449 14887 8483
rect 14829 8443 14887 8449
rect 15102 8440 15108 8492
rect 15160 8480 15166 8492
rect 16117 8483 16175 8489
rect 16117 8480 16129 8483
rect 15160 8452 16129 8480
rect 15160 8440 15166 8452
rect 16117 8449 16129 8452
rect 16163 8449 16175 8483
rect 16117 8443 16175 8449
rect 17218 8440 17224 8492
rect 17276 8440 17282 8492
rect 17313 8483 17371 8489
rect 17313 8449 17325 8483
rect 17359 8480 17371 8483
rect 17957 8483 18015 8489
rect 17957 8480 17969 8483
rect 17359 8452 17969 8480
rect 17359 8449 17371 8452
rect 17313 8443 17371 8449
rect 17957 8449 17969 8452
rect 18003 8480 18015 8483
rect 18230 8480 18236 8492
rect 18003 8452 18236 8480
rect 18003 8449 18015 8452
rect 17957 8443 18015 8449
rect 11422 8372 11428 8424
rect 11480 8412 11486 8424
rect 11701 8415 11759 8421
rect 11701 8412 11713 8415
rect 11480 8384 11713 8412
rect 11480 8372 11486 8384
rect 11701 8381 11713 8384
rect 11747 8381 11759 8415
rect 11701 8375 11759 8381
rect 13173 8415 13231 8421
rect 13173 8381 13185 8415
rect 13219 8412 13231 8415
rect 13354 8412 13360 8424
rect 13219 8384 13360 8412
rect 13219 8381 13231 8384
rect 13173 8375 13231 8381
rect 13354 8372 13360 8384
rect 13412 8372 13418 8424
rect 17328 8412 17356 8443
rect 18230 8440 18236 8452
rect 18288 8440 18294 8492
rect 18414 8440 18420 8492
rect 18472 8440 18478 8492
rect 13464 8384 15240 8412
rect 12802 8304 12808 8356
rect 12860 8344 12866 8356
rect 13464 8344 13492 8384
rect 12860 8316 13492 8344
rect 15212 8344 15240 8384
rect 16408 8384 17356 8412
rect 16408 8344 16436 8384
rect 17402 8372 17408 8424
rect 17460 8372 17466 8424
rect 18874 8412 18880 8424
rect 18156 8384 18880 8412
rect 15212 8316 16436 8344
rect 16853 8347 16911 8353
rect 12860 8304 12866 8316
rect 16853 8313 16865 8347
rect 16899 8344 16911 8347
rect 17770 8344 17776 8356
rect 16899 8316 17776 8344
rect 16899 8313 16911 8316
rect 16853 8307 16911 8313
rect 17770 8304 17776 8316
rect 17828 8304 17834 8356
rect 18156 8344 18184 8384
rect 18874 8372 18880 8384
rect 18932 8372 18938 8424
rect 17880 8316 18184 8344
rect 11974 8236 11980 8288
rect 12032 8276 12038 8288
rect 17880 8276 17908 8316
rect 18230 8304 18236 8356
rect 18288 8344 18294 8356
rect 18506 8344 18512 8356
rect 18288 8316 18512 8344
rect 18288 8304 18294 8316
rect 18506 8304 18512 8316
rect 18564 8304 18570 8356
rect 19168 8344 19196 8520
rect 20272 8520 23664 8548
rect 20272 8489 20300 8520
rect 23658 8508 23664 8520
rect 23716 8508 23722 8560
rect 20257 8483 20315 8489
rect 20257 8449 20269 8483
rect 20303 8449 20315 8483
rect 20257 8443 20315 8449
rect 22186 8440 22192 8492
rect 22244 8440 22250 8492
rect 23952 8489 23980 8588
rect 23937 8483 23995 8489
rect 23937 8449 23949 8483
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 19429 8415 19487 8421
rect 19429 8381 19441 8415
rect 19475 8412 19487 8415
rect 20530 8412 20536 8424
rect 19475 8384 20536 8412
rect 19475 8381 19487 8384
rect 19429 8375 19487 8381
rect 20530 8372 20536 8384
rect 20588 8372 20594 8424
rect 21269 8415 21327 8421
rect 21269 8381 21281 8415
rect 21315 8412 21327 8415
rect 22278 8412 22284 8424
rect 21315 8384 22284 8412
rect 21315 8381 21327 8384
rect 21269 8375 21327 8381
rect 22278 8372 22284 8384
rect 22336 8372 22342 8424
rect 22462 8372 22468 8424
rect 22520 8412 22526 8424
rect 22557 8415 22615 8421
rect 22557 8412 22569 8415
rect 22520 8384 22569 8412
rect 22520 8372 22526 8384
rect 22557 8381 22569 8384
rect 22603 8381 22615 8415
rect 22557 8375 22615 8381
rect 24762 8372 24768 8424
rect 24820 8372 24826 8424
rect 20806 8344 20812 8356
rect 19168 8316 20812 8344
rect 20806 8304 20812 8316
rect 20864 8304 20870 8356
rect 12032 8248 17908 8276
rect 12032 8236 12038 8248
rect 17954 8236 17960 8288
rect 18012 8276 18018 8288
rect 22554 8276 22560 8288
rect 18012 8248 22560 8276
rect 18012 8236 18018 8248
rect 22554 8236 22560 8248
rect 22612 8236 22618 8288
rect 1104 8186 25852 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 25852 8186
rect 1104 8112 25852 8134
rect 11057 8075 11115 8081
rect 11057 8041 11069 8075
rect 11103 8072 11115 8075
rect 11790 8072 11796 8084
rect 11103 8044 11796 8072
rect 11103 8041 11115 8044
rect 11057 8035 11115 8041
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 12989 8075 13047 8081
rect 12989 8041 13001 8075
rect 13035 8072 13047 8075
rect 14277 8075 14335 8081
rect 13035 8044 14228 8072
rect 13035 8041 13047 8044
rect 12989 8035 13047 8041
rect 14200 8004 14228 8044
rect 14277 8041 14289 8075
rect 14323 8072 14335 8075
rect 14323 8044 15332 8072
rect 14323 8041 14335 8044
rect 14277 8035 14335 8041
rect 15304 8004 15332 8044
rect 15838 8032 15844 8084
rect 15896 8032 15902 8084
rect 16114 8032 16120 8084
rect 16172 8072 16178 8084
rect 16390 8072 16396 8084
rect 16172 8044 16396 8072
rect 16172 8032 16178 8044
rect 16390 8032 16396 8044
rect 16448 8032 16454 8084
rect 17770 8032 17776 8084
rect 17828 8072 17834 8084
rect 19058 8072 19064 8084
rect 17828 8044 19064 8072
rect 17828 8032 17834 8044
rect 19058 8032 19064 8044
rect 19116 8032 19122 8084
rect 25314 8072 25320 8084
rect 22066 8044 25320 8072
rect 18782 8004 18788 8016
rect 14200 7976 14964 8004
rect 15304 7976 18788 8004
rect 8386 7896 8392 7948
rect 8444 7936 8450 7948
rect 11701 7939 11759 7945
rect 8444 7908 11652 7936
rect 8444 7896 8450 7908
rect 11422 7828 11428 7880
rect 11480 7828 11486 7880
rect 10318 7760 10324 7812
rect 10376 7800 10382 7812
rect 11517 7803 11575 7809
rect 11517 7800 11529 7803
rect 10376 7772 11529 7800
rect 10376 7760 10382 7772
rect 11517 7769 11529 7772
rect 11563 7769 11575 7803
rect 11624 7800 11652 7908
rect 11701 7905 11713 7939
rect 11747 7936 11759 7939
rect 11974 7936 11980 7948
rect 11747 7908 11980 7936
rect 11747 7905 11759 7908
rect 11701 7899 11759 7905
rect 11974 7896 11980 7908
rect 12032 7896 12038 7948
rect 13633 7939 13691 7945
rect 13633 7905 13645 7939
rect 13679 7936 13691 7939
rect 13998 7936 14004 7948
rect 13679 7908 14004 7936
rect 13679 7905 13691 7908
rect 13633 7899 13691 7905
rect 13998 7896 14004 7908
rect 14056 7896 14062 7948
rect 14826 7896 14832 7948
rect 14884 7896 14890 7948
rect 13354 7828 13360 7880
rect 13412 7828 13418 7880
rect 13722 7828 13728 7880
rect 13780 7868 13786 7880
rect 14458 7868 14464 7880
rect 13780 7840 14464 7868
rect 13780 7828 13786 7840
rect 14458 7828 14464 7840
rect 14516 7828 14522 7880
rect 14642 7828 14648 7880
rect 14700 7828 14706 7880
rect 14936 7868 14964 7976
rect 18782 7964 18788 7976
rect 18840 7964 18846 8016
rect 19610 7964 19616 8016
rect 19668 8004 19674 8016
rect 21818 8004 21824 8016
rect 19668 7976 21824 8004
rect 19668 7964 19674 7976
rect 21818 7964 21824 7976
rect 21876 7964 21882 8016
rect 15746 7896 15752 7948
rect 15804 7936 15810 7948
rect 16393 7939 16451 7945
rect 16393 7936 16405 7939
rect 15804 7908 16405 7936
rect 15804 7896 15810 7908
rect 16393 7905 16405 7908
rect 16439 7905 16451 7939
rect 16393 7899 16451 7905
rect 18693 7939 18751 7945
rect 18693 7905 18705 7939
rect 18739 7936 18751 7939
rect 22066 7936 22094 8044
rect 25314 8032 25320 8044
rect 25372 8032 25378 8084
rect 24857 8007 24915 8013
rect 24857 7973 24869 8007
rect 24903 8004 24915 8007
rect 25038 8004 25044 8016
rect 24903 7976 25044 8004
rect 24903 7973 24915 7976
rect 24857 7967 24915 7973
rect 25038 7964 25044 7976
rect 25096 7964 25102 8016
rect 18739 7908 22094 7936
rect 18739 7905 18751 7908
rect 18693 7899 18751 7905
rect 22370 7896 22376 7948
rect 22428 7896 22434 7948
rect 16574 7868 16580 7880
rect 14936 7840 16580 7868
rect 16574 7828 16580 7840
rect 16632 7828 16638 7880
rect 17681 7871 17739 7877
rect 17681 7837 17693 7871
rect 17727 7868 17739 7871
rect 17954 7868 17960 7880
rect 17727 7840 17960 7868
rect 17727 7837 17739 7840
rect 17681 7831 17739 7837
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 20441 7871 20499 7877
rect 20441 7837 20453 7871
rect 20487 7868 20499 7871
rect 20487 7840 21128 7868
rect 20487 7837 20499 7840
rect 20441 7831 20499 7837
rect 13449 7803 13507 7809
rect 13449 7800 13461 7803
rect 11624 7772 13461 7800
rect 11517 7763 11575 7769
rect 13449 7769 13461 7772
rect 13495 7769 13507 7803
rect 14737 7803 14795 7809
rect 14737 7800 14749 7803
rect 13449 7763 13507 7769
rect 13740 7772 14749 7800
rect 12345 7735 12403 7741
rect 12345 7701 12357 7735
rect 12391 7732 12403 7735
rect 12618 7732 12624 7744
rect 12391 7704 12624 7732
rect 12391 7701 12403 7704
rect 12345 7695 12403 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 13354 7692 13360 7744
rect 13412 7732 13418 7744
rect 13740 7732 13768 7772
rect 14737 7769 14749 7772
rect 14783 7769 14795 7803
rect 14737 7763 14795 7769
rect 15286 7760 15292 7812
rect 15344 7800 15350 7812
rect 15381 7803 15439 7809
rect 15381 7800 15393 7803
rect 15344 7772 15393 7800
rect 15344 7760 15350 7772
rect 15381 7769 15393 7772
rect 15427 7800 15439 7803
rect 15838 7800 15844 7812
rect 15427 7772 15844 7800
rect 15427 7769 15439 7772
rect 15381 7763 15439 7769
rect 15838 7760 15844 7772
rect 15896 7760 15902 7812
rect 16209 7803 16267 7809
rect 16209 7769 16221 7803
rect 16255 7800 16267 7803
rect 20714 7800 20720 7812
rect 16255 7772 20720 7800
rect 16255 7769 16267 7772
rect 16209 7763 16267 7769
rect 20714 7760 20720 7772
rect 20772 7760 20778 7812
rect 13412 7704 13768 7732
rect 13412 7692 13418 7704
rect 13998 7692 14004 7744
rect 14056 7732 14062 7744
rect 15194 7732 15200 7744
rect 14056 7704 15200 7732
rect 14056 7692 14062 7704
rect 15194 7692 15200 7704
rect 15252 7692 15258 7744
rect 15654 7692 15660 7744
rect 15712 7732 15718 7744
rect 16301 7735 16359 7741
rect 16301 7732 16313 7735
rect 15712 7704 16313 7732
rect 15712 7692 15718 7704
rect 16301 7701 16313 7704
rect 16347 7701 16359 7735
rect 16301 7695 16359 7701
rect 18782 7692 18788 7744
rect 18840 7732 18846 7744
rect 19429 7735 19487 7741
rect 19429 7732 19441 7735
rect 18840 7704 19441 7732
rect 18840 7692 18846 7704
rect 19429 7701 19441 7704
rect 19475 7701 19487 7735
rect 19429 7695 19487 7701
rect 19886 7692 19892 7744
rect 19944 7692 19950 7744
rect 21100 7732 21128 7840
rect 21818 7828 21824 7880
rect 21876 7868 21882 7880
rect 22094 7868 22100 7880
rect 21876 7840 22100 7868
rect 21876 7828 21882 7840
rect 22094 7828 22100 7840
rect 22152 7828 22158 7880
rect 24026 7868 24032 7880
rect 23506 7840 24032 7868
rect 24026 7828 24032 7840
rect 24084 7868 24090 7880
rect 24210 7868 24216 7880
rect 24084 7840 24216 7868
rect 24084 7828 24090 7840
rect 24210 7828 24216 7840
rect 24268 7828 24274 7880
rect 21453 7803 21511 7809
rect 21453 7769 21465 7803
rect 21499 7800 21511 7803
rect 21634 7800 21640 7812
rect 21499 7772 21640 7800
rect 21499 7769 21511 7772
rect 21453 7763 21511 7769
rect 21634 7760 21640 7772
rect 21692 7760 21698 7812
rect 24673 7803 24731 7809
rect 24673 7800 24685 7803
rect 23676 7772 24685 7800
rect 22370 7732 22376 7744
rect 21100 7704 22376 7732
rect 22370 7692 22376 7704
rect 22428 7692 22434 7744
rect 23382 7692 23388 7744
rect 23440 7732 23446 7744
rect 23676 7732 23704 7772
rect 24673 7769 24685 7772
rect 24719 7769 24731 7803
rect 24673 7763 24731 7769
rect 23440 7704 23704 7732
rect 23440 7692 23446 7704
rect 23842 7692 23848 7744
rect 23900 7692 23906 7744
rect 24210 7692 24216 7744
rect 24268 7692 24274 7744
rect 1104 7642 25852 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 25852 7642
rect 1104 7568 25852 7590
rect 11974 7488 11980 7540
rect 12032 7488 12038 7540
rect 12618 7488 12624 7540
rect 12676 7488 12682 7540
rect 13630 7488 13636 7540
rect 13688 7528 13694 7540
rect 15473 7531 15531 7537
rect 15473 7528 15485 7531
rect 13688 7500 15485 7528
rect 13688 7488 13694 7500
rect 15473 7497 15485 7500
rect 15519 7497 15531 7531
rect 15473 7491 15531 7497
rect 17773 7531 17831 7537
rect 17773 7497 17785 7531
rect 17819 7528 17831 7531
rect 18322 7528 18328 7540
rect 17819 7500 18328 7528
rect 17819 7497 17831 7500
rect 17773 7491 17831 7497
rect 18322 7488 18328 7500
rect 18380 7488 18386 7540
rect 19058 7488 19064 7540
rect 19116 7528 19122 7540
rect 21177 7531 21235 7537
rect 21177 7528 21189 7531
rect 19116 7500 21189 7528
rect 19116 7488 19122 7500
rect 21177 7497 21189 7500
rect 21223 7497 21235 7531
rect 21177 7491 21235 7497
rect 23474 7488 23480 7540
rect 23532 7488 23538 7540
rect 11057 7463 11115 7469
rect 11057 7460 11069 7463
rect 10534 7432 11069 7460
rect 11057 7429 11069 7432
rect 11103 7460 11115 7463
rect 11514 7460 11520 7472
rect 11103 7432 11520 7460
rect 11103 7429 11115 7432
rect 11057 7423 11115 7429
rect 11514 7420 11520 7432
rect 11572 7420 11578 7472
rect 12066 7420 12072 7472
rect 12124 7460 12130 7472
rect 14274 7460 14280 7472
rect 12124 7432 14280 7460
rect 12124 7420 12130 7432
rect 14274 7420 14280 7432
rect 14332 7420 14338 7472
rect 14458 7420 14464 7472
rect 14516 7420 14522 7472
rect 16117 7463 16175 7469
rect 16117 7429 16129 7463
rect 16163 7460 16175 7463
rect 16298 7460 16304 7472
rect 16163 7432 16304 7460
rect 16163 7429 16175 7432
rect 16117 7423 16175 7429
rect 16298 7420 16304 7432
rect 16356 7460 16362 7472
rect 16853 7463 16911 7469
rect 16853 7460 16865 7463
rect 16356 7432 16865 7460
rect 16356 7420 16362 7432
rect 16853 7429 16865 7432
rect 16899 7429 16911 7463
rect 16853 7423 16911 7429
rect 17681 7463 17739 7469
rect 17681 7429 17693 7463
rect 17727 7460 17739 7463
rect 18874 7460 18880 7472
rect 17727 7432 18880 7460
rect 17727 7429 17739 7432
rect 17681 7423 17739 7429
rect 18874 7420 18880 7432
rect 18932 7420 18938 7472
rect 20346 7420 20352 7472
rect 20404 7460 20410 7472
rect 20533 7463 20591 7469
rect 20533 7460 20545 7463
rect 20404 7432 20545 7460
rect 20404 7420 20410 7432
rect 20533 7429 20545 7432
rect 20579 7460 20591 7463
rect 21085 7463 21143 7469
rect 21085 7460 21097 7463
rect 20579 7432 21097 7460
rect 20579 7429 20591 7432
rect 20533 7423 20591 7429
rect 21085 7429 21097 7432
rect 21131 7429 21143 7463
rect 23492 7460 23520 7488
rect 21085 7423 21143 7429
rect 22296 7432 23520 7460
rect 19886 7352 19892 7404
rect 19944 7352 19950 7404
rect 20714 7352 20720 7404
rect 20772 7392 20778 7404
rect 21910 7392 21916 7404
rect 20772 7364 21916 7392
rect 20772 7352 20778 7364
rect 21910 7352 21916 7364
rect 21968 7392 21974 7404
rect 22296 7401 22324 7432
rect 25130 7420 25136 7472
rect 25188 7420 25194 7472
rect 22281 7395 22339 7401
rect 21968 7364 22094 7392
rect 21968 7352 21974 7364
rect 9030 7284 9036 7336
rect 9088 7284 9094 7336
rect 9309 7327 9367 7333
rect 9309 7293 9321 7327
rect 9355 7324 9367 7327
rect 10962 7324 10968 7336
rect 9355 7296 10968 7324
rect 9355 7293 9367 7296
rect 9309 7287 9367 7293
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11146 7284 11152 7336
rect 11204 7324 11210 7336
rect 12713 7327 12771 7333
rect 12713 7324 12725 7327
rect 11204 7296 12725 7324
rect 11204 7284 11210 7296
rect 12713 7293 12725 7296
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7293 12863 7327
rect 12805 7287 12863 7293
rect 13725 7327 13783 7333
rect 13725 7293 13737 7327
rect 13771 7293 13783 7327
rect 13725 7287 13783 7293
rect 14001 7327 14059 7333
rect 14001 7293 14013 7327
rect 14047 7324 14059 7327
rect 16666 7324 16672 7336
rect 14047 7296 16672 7324
rect 14047 7293 14059 7296
rect 14001 7287 14059 7293
rect 10778 7216 10784 7268
rect 10836 7256 10842 7268
rect 12820 7256 12848 7287
rect 10836 7228 12848 7256
rect 10836 7216 10842 7228
rect 12253 7191 12311 7197
rect 12253 7157 12265 7191
rect 12299 7188 12311 7191
rect 13446 7188 13452 7200
rect 12299 7160 13452 7188
rect 12299 7157 12311 7160
rect 12253 7151 12311 7157
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 13740 7188 13768 7287
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 17586 7284 17592 7336
rect 17644 7324 17650 7336
rect 17865 7327 17923 7333
rect 17865 7324 17877 7327
rect 17644 7296 17877 7324
rect 17644 7284 17650 7296
rect 17865 7293 17877 7296
rect 17911 7293 17923 7327
rect 17865 7287 17923 7293
rect 16301 7259 16359 7265
rect 16301 7225 16313 7259
rect 16347 7256 16359 7259
rect 17770 7256 17776 7268
rect 16347 7228 17776 7256
rect 16347 7225 16359 7228
rect 16301 7219 16359 7225
rect 17770 7216 17776 7228
rect 17828 7216 17834 7268
rect 15102 7188 15108 7200
rect 13740 7160 15108 7188
rect 15102 7148 15108 7160
rect 15160 7148 15166 7200
rect 16666 7148 16672 7200
rect 16724 7148 16730 7200
rect 17034 7148 17040 7200
rect 17092 7188 17098 7200
rect 17313 7191 17371 7197
rect 17313 7188 17325 7191
rect 17092 7160 17325 7188
rect 17092 7148 17098 7160
rect 17313 7157 17325 7160
rect 17359 7157 17371 7191
rect 17880 7188 17908 7287
rect 18506 7284 18512 7336
rect 18564 7284 18570 7336
rect 18785 7327 18843 7333
rect 18785 7293 18797 7327
rect 18831 7324 18843 7327
rect 19242 7324 19248 7336
rect 18831 7296 19248 7324
rect 18831 7293 18843 7296
rect 18785 7287 18843 7293
rect 19242 7284 19248 7296
rect 19300 7284 19306 7336
rect 19794 7284 19800 7336
rect 19852 7324 19858 7336
rect 21269 7327 21327 7333
rect 21269 7324 21281 7327
rect 19852 7296 21281 7324
rect 19852 7284 19858 7296
rect 21269 7293 21281 7296
rect 21315 7293 21327 7327
rect 21269 7287 21327 7293
rect 22066 7256 22094 7364
rect 22281 7361 22293 7395
rect 22327 7361 22339 7395
rect 22281 7355 22339 7361
rect 23474 7352 23480 7404
rect 23532 7392 23538 7404
rect 23937 7395 23995 7401
rect 23937 7392 23949 7395
rect 23532 7364 23949 7392
rect 23532 7352 23538 7364
rect 23937 7361 23949 7364
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 23293 7327 23351 7333
rect 23293 7293 23305 7327
rect 23339 7324 23351 7327
rect 24854 7324 24860 7336
rect 23339 7296 24860 7324
rect 23339 7293 23351 7296
rect 23293 7287 23351 7293
rect 24854 7284 24860 7296
rect 24912 7284 24918 7336
rect 23566 7256 23572 7268
rect 22066 7228 23572 7256
rect 23566 7216 23572 7228
rect 23624 7216 23630 7268
rect 20257 7191 20315 7197
rect 20257 7188 20269 7191
rect 17880 7160 20269 7188
rect 17313 7151 17371 7157
rect 20257 7157 20269 7160
rect 20303 7157 20315 7191
rect 20257 7151 20315 7157
rect 20717 7191 20775 7197
rect 20717 7157 20729 7191
rect 20763 7188 20775 7191
rect 22830 7188 22836 7200
rect 20763 7160 22836 7188
rect 20763 7157 20775 7160
rect 20717 7151 20775 7157
rect 22830 7148 22836 7160
rect 22888 7148 22894 7200
rect 1104 7098 25852 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 25852 7098
rect 1104 7024 25852 7046
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 12529 6987 12587 6993
rect 12529 6984 12541 6987
rect 12400 6956 12541 6984
rect 12400 6944 12406 6956
rect 12529 6953 12541 6956
rect 12575 6984 12587 6987
rect 14826 6984 14832 6996
rect 12575 6956 14832 6984
rect 12575 6953 12587 6956
rect 12529 6947 12587 6953
rect 14826 6944 14832 6956
rect 14884 6944 14890 6996
rect 19886 6984 19892 6996
rect 18432 6956 19892 6984
rect 14642 6916 14648 6928
rect 14476 6888 14648 6916
rect 10781 6851 10839 6857
rect 10781 6817 10793 6851
rect 10827 6848 10839 6851
rect 11698 6848 11704 6860
rect 10827 6820 11704 6848
rect 10827 6817 10839 6820
rect 10781 6811 10839 6817
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 14182 6808 14188 6860
rect 14240 6848 14246 6860
rect 14476 6848 14504 6888
rect 14642 6876 14648 6888
rect 14700 6876 14706 6928
rect 14240 6820 14504 6848
rect 14240 6808 14246 6820
rect 17402 6808 17408 6860
rect 17460 6808 17466 6860
rect 17862 6808 17868 6860
rect 17920 6848 17926 6860
rect 18432 6848 18460 6956
rect 19886 6944 19892 6956
rect 19944 6984 19950 6996
rect 20162 6984 20168 6996
rect 19944 6956 20168 6984
rect 19944 6944 19950 6956
rect 20162 6944 20168 6956
rect 20220 6984 20226 6996
rect 20441 6987 20499 6993
rect 20441 6984 20453 6987
rect 20220 6956 20453 6984
rect 20220 6944 20226 6956
rect 20441 6953 20453 6956
rect 20487 6953 20499 6987
rect 20441 6947 20499 6953
rect 18506 6876 18512 6928
rect 18564 6916 18570 6928
rect 19610 6916 19616 6928
rect 18564 6888 19616 6916
rect 18564 6876 18570 6888
rect 19610 6876 19616 6888
rect 19668 6876 19674 6928
rect 19794 6876 19800 6928
rect 19852 6876 19858 6928
rect 23842 6876 23848 6928
rect 23900 6916 23906 6928
rect 23900 6888 25176 6916
rect 23900 6876 23906 6888
rect 17920 6820 18460 6848
rect 18877 6851 18935 6857
rect 17920 6808 17926 6820
rect 18877 6817 18889 6851
rect 18923 6848 18935 6851
rect 19812 6848 19840 6876
rect 18923 6820 19840 6848
rect 18923 6817 18935 6820
rect 18877 6811 18935 6817
rect 19886 6808 19892 6860
rect 19944 6808 19950 6860
rect 20073 6851 20131 6857
rect 20073 6817 20085 6851
rect 20119 6817 20131 6851
rect 20073 6811 20131 6817
rect 13722 6740 13728 6792
rect 13780 6740 13786 6792
rect 15470 6740 15476 6792
rect 15528 6740 15534 6792
rect 16942 6740 16948 6792
rect 17000 6780 17006 6792
rect 17129 6783 17187 6789
rect 17129 6780 17141 6783
rect 17000 6752 17141 6780
rect 17000 6740 17006 6752
rect 17129 6749 17141 6752
rect 17175 6749 17187 6783
rect 19518 6780 19524 6792
rect 17129 6743 17187 6749
rect 19306 6752 19524 6780
rect 11054 6672 11060 6724
rect 11112 6672 11118 6724
rect 11514 6712 11520 6724
rect 11440 6684 11520 6712
rect 11440 6644 11468 6684
rect 11514 6672 11520 6684
rect 11572 6672 11578 6724
rect 14642 6672 14648 6724
rect 14700 6672 14706 6724
rect 16485 6715 16543 6721
rect 16485 6681 16497 6715
rect 16531 6681 16543 6715
rect 16485 6675 16543 6681
rect 12434 6644 12440 6656
rect 11440 6616 12440 6644
rect 12434 6604 12440 6616
rect 12492 6644 12498 6656
rect 12805 6647 12863 6653
rect 12805 6644 12817 6647
rect 12492 6616 12817 6644
rect 12492 6604 12498 6616
rect 12805 6613 12817 6616
rect 12851 6613 12863 6647
rect 12805 6607 12863 6613
rect 13538 6604 13544 6656
rect 13596 6604 13602 6656
rect 14274 6604 14280 6656
rect 14332 6644 14338 6656
rect 14737 6647 14795 6653
rect 14737 6644 14749 6647
rect 14332 6616 14749 6644
rect 14332 6604 14338 6616
rect 14737 6613 14749 6616
rect 14783 6613 14795 6647
rect 16500 6644 16528 6675
rect 16666 6672 16672 6724
rect 16724 6712 16730 6724
rect 17862 6712 17868 6724
rect 16724 6684 17868 6712
rect 16724 6672 16730 6684
rect 17862 6672 17868 6684
rect 17920 6672 17926 6724
rect 19306 6644 19334 6752
rect 19518 6740 19524 6752
rect 19576 6740 19582 6792
rect 20088 6780 20116 6811
rect 20438 6808 20444 6860
rect 20496 6848 20502 6860
rect 20496 6820 22692 6848
rect 20496 6808 20502 6820
rect 20254 6780 20260 6792
rect 20088 6752 20260 6780
rect 20254 6740 20260 6752
rect 20312 6740 20318 6792
rect 20901 6783 20959 6789
rect 20901 6749 20913 6783
rect 20947 6780 20959 6783
rect 21542 6780 21548 6792
rect 20947 6752 21548 6780
rect 20947 6749 20959 6752
rect 20901 6743 20959 6749
rect 21542 6740 21548 6752
rect 21600 6740 21606 6792
rect 21726 6740 21732 6792
rect 21784 6780 21790 6792
rect 21910 6780 21916 6792
rect 21784 6752 21916 6780
rect 21784 6740 21790 6752
rect 21910 6740 21916 6752
rect 21968 6740 21974 6792
rect 22664 6789 22692 6820
rect 23290 6808 23296 6860
rect 23348 6848 23354 6860
rect 24026 6848 24032 6860
rect 23348 6820 24032 6848
rect 23348 6808 23354 6820
rect 24026 6808 24032 6820
rect 24084 6808 24090 6860
rect 24486 6808 24492 6860
rect 24544 6848 24550 6860
rect 25148 6857 25176 6888
rect 25041 6851 25099 6857
rect 25041 6848 25053 6851
rect 24544 6820 25053 6848
rect 24544 6808 24550 6820
rect 25041 6817 25053 6820
rect 25087 6817 25099 6851
rect 25041 6811 25099 6817
rect 25133 6851 25191 6857
rect 25133 6817 25145 6851
rect 25179 6817 25191 6851
rect 25133 6811 25191 6817
rect 22649 6783 22707 6789
rect 22649 6749 22661 6783
rect 22695 6749 22707 6783
rect 22649 6743 22707 6749
rect 21821 6715 21879 6721
rect 21821 6681 21833 6715
rect 21867 6712 21879 6715
rect 23845 6715 23903 6721
rect 21867 6684 21956 6712
rect 21867 6681 21879 6684
rect 21821 6675 21879 6681
rect 16500 6616 19334 6644
rect 19429 6647 19487 6653
rect 14737 6607 14795 6613
rect 19429 6613 19441 6647
rect 19475 6644 19487 6647
rect 19518 6644 19524 6656
rect 19475 6616 19524 6644
rect 19475 6613 19487 6616
rect 19429 6607 19487 6613
rect 19518 6604 19524 6616
rect 19576 6604 19582 6656
rect 19794 6604 19800 6656
rect 19852 6604 19858 6656
rect 21928 6644 21956 6684
rect 23845 6681 23857 6715
rect 23891 6712 23903 6715
rect 25130 6712 25136 6724
rect 23891 6684 25136 6712
rect 23891 6681 23903 6684
rect 23845 6675 23903 6681
rect 25130 6672 25136 6684
rect 25188 6672 25194 6724
rect 23290 6644 23296 6656
rect 21928 6616 23296 6644
rect 23290 6604 23296 6616
rect 23348 6604 23354 6656
rect 23382 6604 23388 6656
rect 23440 6644 23446 6656
rect 24581 6647 24639 6653
rect 24581 6644 24593 6647
rect 23440 6616 24593 6644
rect 23440 6604 23446 6616
rect 24581 6613 24593 6616
rect 24627 6613 24639 6647
rect 24581 6607 24639 6613
rect 24854 6604 24860 6656
rect 24912 6644 24918 6656
rect 24949 6647 25007 6653
rect 24949 6644 24961 6647
rect 24912 6616 24961 6644
rect 24912 6604 24918 6616
rect 24949 6613 24961 6616
rect 24995 6613 25007 6647
rect 24949 6607 25007 6613
rect 1104 6554 25852 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 25852 6554
rect 1104 6480 25852 6502
rect 10413 6443 10471 6449
rect 10413 6409 10425 6443
rect 10459 6440 10471 6443
rect 11146 6440 11152 6452
rect 10459 6412 11152 6440
rect 10459 6409 10471 6412
rect 10413 6403 10471 6409
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 12161 6443 12219 6449
rect 12161 6409 12173 6443
rect 12207 6440 12219 6443
rect 12802 6440 12808 6452
rect 12207 6412 12808 6440
rect 12207 6409 12219 6412
rect 12161 6403 12219 6409
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 13357 6443 13415 6449
rect 13357 6409 13369 6443
rect 13403 6440 13415 6443
rect 17313 6443 17371 6449
rect 17313 6440 17325 6443
rect 13403 6412 17325 6440
rect 13403 6409 13415 6412
rect 13357 6403 13415 6409
rect 17313 6409 17325 6412
rect 17359 6409 17371 6443
rect 17313 6403 17371 6409
rect 17862 6400 17868 6452
rect 17920 6440 17926 6452
rect 17957 6443 18015 6449
rect 17957 6440 17969 6443
rect 17920 6412 17969 6440
rect 17920 6400 17926 6412
rect 17957 6409 17969 6412
rect 18003 6409 18015 6443
rect 17957 6403 18015 6409
rect 18322 6400 18328 6452
rect 18380 6440 18386 6452
rect 18380 6412 19334 6440
rect 18380 6400 18386 6412
rect 10873 6375 10931 6381
rect 10873 6341 10885 6375
rect 10919 6372 10931 6375
rect 10919 6344 12434 6372
rect 10919 6341 10931 6344
rect 10873 6335 10931 6341
rect 6362 6264 6368 6316
rect 6420 6304 6426 6316
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 6420 6276 10793 6304
rect 6420 6264 6426 6276
rect 10781 6273 10793 6276
rect 10827 6273 10839 6307
rect 10781 6267 10839 6273
rect 11146 6264 11152 6316
rect 11204 6304 11210 6316
rect 12069 6307 12127 6313
rect 12069 6304 12081 6307
rect 11204 6276 12081 6304
rect 11204 6264 11210 6276
rect 12069 6273 12081 6276
rect 12115 6273 12127 6307
rect 12069 6267 12127 6273
rect 10962 6196 10968 6248
rect 11020 6196 11026 6248
rect 12250 6196 12256 6248
rect 12308 6196 12314 6248
rect 12406 6236 12434 6344
rect 13998 6332 14004 6384
rect 14056 6372 14062 6384
rect 19306 6372 19334 6412
rect 19518 6400 19524 6452
rect 19576 6440 19582 6452
rect 20346 6440 20352 6452
rect 19576 6412 20352 6440
rect 19576 6400 19582 6412
rect 20346 6400 20352 6412
rect 20404 6400 20410 6452
rect 22646 6440 22652 6452
rect 20548 6412 22652 6440
rect 20438 6372 20444 6384
rect 14056 6344 18276 6372
rect 19306 6344 20444 6372
rect 14056 6332 14062 6344
rect 12710 6264 12716 6316
rect 12768 6304 12774 6316
rect 13725 6307 13783 6313
rect 13725 6304 13737 6307
rect 12768 6276 13737 6304
rect 12768 6264 12774 6276
rect 13725 6273 13737 6276
rect 13771 6273 13783 6307
rect 13725 6267 13783 6273
rect 13817 6307 13875 6313
rect 13817 6273 13829 6307
rect 13863 6304 13875 6307
rect 14182 6304 14188 6316
rect 13863 6276 14188 6304
rect 13863 6273 13875 6276
rect 13817 6267 13875 6273
rect 14182 6264 14188 6276
rect 14240 6304 14246 6316
rect 14369 6307 14427 6313
rect 14369 6304 14381 6307
rect 14240 6276 14381 6304
rect 14240 6264 14246 6276
rect 14369 6273 14381 6276
rect 14415 6273 14427 6307
rect 14369 6267 14427 6273
rect 15105 6307 15163 6313
rect 15105 6273 15117 6307
rect 15151 6304 15163 6307
rect 15151 6276 17172 6304
rect 15151 6273 15163 6276
rect 15105 6267 15163 6273
rect 12406 6208 13492 6236
rect 2682 6128 2688 6180
rect 2740 6168 2746 6180
rect 10318 6168 10324 6180
rect 2740 6140 10324 6168
rect 2740 6128 2746 6140
rect 10318 6128 10324 6140
rect 10376 6128 10382 6180
rect 11701 6171 11759 6177
rect 11701 6137 11713 6171
rect 11747 6168 11759 6171
rect 13354 6168 13360 6180
rect 11747 6140 13360 6168
rect 11747 6137 11759 6140
rect 11701 6131 11759 6137
rect 13354 6128 13360 6140
rect 13412 6128 13418 6180
rect 12989 6103 13047 6109
rect 12989 6069 13001 6103
rect 13035 6100 13047 6103
rect 13464 6100 13492 6208
rect 13630 6196 13636 6248
rect 13688 6236 13694 6248
rect 13909 6239 13967 6245
rect 13909 6236 13921 6239
rect 13688 6208 13921 6236
rect 13688 6196 13694 6208
rect 13909 6205 13921 6208
rect 13955 6205 13967 6239
rect 13909 6199 13967 6205
rect 16114 6196 16120 6248
rect 16172 6196 16178 6248
rect 13722 6128 13728 6180
rect 13780 6168 13786 6180
rect 16853 6171 16911 6177
rect 16853 6168 16865 6171
rect 13780 6140 16865 6168
rect 13780 6128 13786 6140
rect 16853 6137 16865 6140
rect 16899 6137 16911 6171
rect 17144 6168 17172 6276
rect 17218 6264 17224 6316
rect 17276 6264 17282 6316
rect 18248 6313 18276 6344
rect 20438 6332 20444 6344
rect 20496 6332 20502 6384
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 20257 6307 20315 6313
rect 20257 6273 20269 6307
rect 20303 6304 20315 6307
rect 20548 6304 20576 6412
rect 22646 6400 22652 6412
rect 22704 6400 22710 6452
rect 23750 6400 23756 6452
rect 23808 6440 23814 6452
rect 24581 6443 24639 6449
rect 24581 6440 24593 6443
rect 23808 6412 24593 6440
rect 23808 6400 23814 6412
rect 24581 6409 24593 6412
rect 24627 6409 24639 6443
rect 24581 6403 24639 6409
rect 22554 6372 22560 6384
rect 20303 6276 20576 6304
rect 20640 6344 22560 6372
rect 20303 6273 20315 6276
rect 20257 6267 20315 6273
rect 17310 6196 17316 6248
rect 17368 6236 17374 6248
rect 17405 6239 17463 6245
rect 17405 6236 17417 6239
rect 17368 6208 17417 6236
rect 17368 6196 17374 6208
rect 17405 6205 17417 6208
rect 17451 6205 17463 6239
rect 17405 6199 17463 6205
rect 19429 6239 19487 6245
rect 19429 6205 19441 6239
rect 19475 6236 19487 6239
rect 20640 6236 20668 6344
rect 22554 6332 22560 6344
rect 22612 6332 22618 6384
rect 22002 6264 22008 6316
rect 22060 6264 22066 6316
rect 23414 6276 23980 6304
rect 19475 6208 20668 6236
rect 21269 6239 21327 6245
rect 19475 6205 19487 6208
rect 19429 6199 19487 6205
rect 21269 6205 21281 6239
rect 21315 6236 21327 6239
rect 21726 6236 21732 6248
rect 21315 6208 21732 6236
rect 21315 6205 21327 6208
rect 21269 6199 21327 6205
rect 21726 6196 21732 6208
rect 21784 6196 21790 6248
rect 22281 6239 22339 6245
rect 22281 6205 22293 6239
rect 22327 6236 22339 6239
rect 23842 6236 23848 6248
rect 22327 6208 23848 6236
rect 22327 6205 22339 6208
rect 22281 6199 22339 6205
rect 23842 6196 23848 6208
rect 23900 6196 23906 6248
rect 22002 6168 22008 6180
rect 17144 6140 22008 6168
rect 16853 6131 16911 6137
rect 22002 6128 22008 6140
rect 22060 6128 22066 6180
rect 23952 6168 23980 6276
rect 24118 6264 24124 6316
rect 24176 6304 24182 6316
rect 24765 6307 24823 6313
rect 24765 6304 24777 6307
rect 24176 6276 24777 6304
rect 24176 6264 24182 6276
rect 24765 6273 24777 6276
rect 24811 6273 24823 6307
rect 24765 6267 24823 6273
rect 23952 6140 24164 6168
rect 24136 6112 24164 6140
rect 15194 6100 15200 6112
rect 13035 6072 15200 6100
rect 13035 6069 13047 6072
rect 12989 6063 13047 6069
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 15654 6060 15660 6112
rect 15712 6100 15718 6112
rect 19610 6100 19616 6112
rect 15712 6072 19616 6100
rect 15712 6060 15718 6072
rect 19610 6060 19616 6072
rect 19668 6060 19674 6112
rect 19794 6060 19800 6112
rect 19852 6100 19858 6112
rect 20254 6100 20260 6112
rect 19852 6072 20260 6100
rect 19852 6060 19858 6072
rect 20254 6060 20260 6072
rect 20312 6100 20318 6112
rect 23753 6103 23811 6109
rect 23753 6100 23765 6103
rect 20312 6072 23765 6100
rect 20312 6060 20318 6072
rect 23753 6069 23765 6072
rect 23799 6069 23811 6103
rect 23753 6063 23811 6069
rect 23842 6060 23848 6112
rect 23900 6100 23906 6112
rect 24029 6103 24087 6109
rect 24029 6100 24041 6103
rect 23900 6072 24041 6100
rect 23900 6060 23906 6072
rect 24029 6069 24041 6072
rect 24075 6069 24087 6103
rect 24029 6063 24087 6069
rect 24118 6060 24124 6112
rect 24176 6100 24182 6112
rect 24213 6103 24271 6109
rect 24213 6100 24225 6103
rect 24176 6072 24225 6100
rect 24176 6060 24182 6072
rect 24213 6069 24225 6072
rect 24259 6069 24271 6103
rect 24213 6063 24271 6069
rect 1104 6010 25852 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 25852 6010
rect 1104 5936 25852 5958
rect 11054 5856 11060 5908
rect 11112 5896 11118 5908
rect 11793 5899 11851 5905
rect 11793 5896 11805 5899
rect 11112 5868 11805 5896
rect 11112 5856 11118 5868
rect 11793 5865 11805 5868
rect 11839 5896 11851 5899
rect 12250 5896 12256 5908
rect 11839 5868 12256 5896
rect 11839 5865 11851 5868
rect 11793 5859 11851 5865
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 13541 5899 13599 5905
rect 13541 5865 13553 5899
rect 13587 5896 13599 5899
rect 13998 5896 14004 5908
rect 13587 5868 14004 5896
rect 13587 5865 13599 5868
rect 13541 5859 13599 5865
rect 13998 5856 14004 5868
rect 14056 5856 14062 5908
rect 14185 5899 14243 5905
rect 14185 5865 14197 5899
rect 14231 5896 14243 5899
rect 14366 5896 14372 5908
rect 14231 5868 14372 5896
rect 14231 5865 14243 5868
rect 14185 5859 14243 5865
rect 14366 5856 14372 5868
rect 14424 5856 14430 5908
rect 14737 5899 14795 5905
rect 14737 5865 14749 5899
rect 14783 5896 14795 5899
rect 14783 5868 17264 5896
rect 14783 5865 14795 5868
rect 14737 5859 14795 5865
rect 11330 5788 11336 5840
rect 11388 5828 11394 5840
rect 15930 5828 15936 5840
rect 11388 5800 15936 5828
rect 11388 5788 11394 5800
rect 15930 5788 15936 5800
rect 15988 5788 15994 5840
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5760 10379 5763
rect 10778 5760 10784 5772
rect 10367 5732 10784 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 10778 5720 10784 5732
rect 10836 5720 10842 5772
rect 12158 5720 12164 5772
rect 12216 5760 12222 5772
rect 12253 5763 12311 5769
rect 12253 5760 12265 5763
rect 12216 5732 12265 5760
rect 12216 5720 12222 5732
rect 12253 5729 12265 5732
rect 12299 5729 12311 5763
rect 14461 5763 14519 5769
rect 12253 5723 12311 5729
rect 12406 5732 13768 5760
rect 9030 5652 9036 5704
rect 9088 5692 9094 5704
rect 9582 5692 9588 5704
rect 9088 5664 9588 5692
rect 9088 5652 9094 5664
rect 9582 5652 9588 5664
rect 9640 5692 9646 5704
rect 10045 5695 10103 5701
rect 10045 5692 10057 5695
rect 9640 5664 10057 5692
rect 9640 5652 9646 5664
rect 10045 5661 10057 5664
rect 10091 5661 10103 5695
rect 10045 5655 10103 5661
rect 11606 5652 11612 5704
rect 11664 5692 11670 5704
rect 12406 5692 12434 5732
rect 11664 5664 12434 5692
rect 11664 5652 11670 5664
rect 12526 5652 12532 5704
rect 12584 5652 12590 5704
rect 13740 5701 13768 5732
rect 14461 5729 14473 5763
rect 14507 5760 14519 5763
rect 15194 5760 15200 5772
rect 14507 5732 15200 5760
rect 14507 5729 14519 5732
rect 14461 5723 14519 5729
rect 15194 5720 15200 5732
rect 15252 5720 15258 5772
rect 15378 5720 15384 5772
rect 15436 5720 15442 5772
rect 16942 5760 16948 5772
rect 15948 5732 16948 5760
rect 13725 5695 13783 5701
rect 13725 5661 13737 5695
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 15102 5652 15108 5704
rect 15160 5692 15166 5704
rect 15948 5701 15976 5732
rect 16942 5720 16948 5732
rect 17000 5720 17006 5772
rect 17236 5760 17264 5868
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 17460 5868 17693 5896
rect 17460 5856 17466 5868
rect 17681 5865 17693 5868
rect 17727 5865 17739 5899
rect 17681 5859 17739 5865
rect 19978 5856 19984 5908
rect 20036 5896 20042 5908
rect 21542 5896 21548 5908
rect 20036 5868 21548 5896
rect 20036 5856 20042 5868
rect 21542 5856 21548 5868
rect 21600 5856 21606 5908
rect 21910 5856 21916 5908
rect 21968 5896 21974 5908
rect 23845 5899 23903 5905
rect 23845 5896 23857 5899
rect 21968 5868 23857 5896
rect 21968 5856 21974 5868
rect 23845 5865 23857 5868
rect 23891 5865 23903 5899
rect 23845 5859 23903 5865
rect 25222 5856 25228 5908
rect 25280 5856 25286 5908
rect 18141 5831 18199 5837
rect 18141 5797 18153 5831
rect 18187 5828 18199 5831
rect 18187 5800 20576 5828
rect 18187 5797 18199 5800
rect 18141 5791 18199 5797
rect 18601 5763 18659 5769
rect 18601 5760 18613 5763
rect 17236 5732 18613 5760
rect 18601 5729 18613 5732
rect 18647 5729 18659 5763
rect 18601 5723 18659 5729
rect 18693 5763 18751 5769
rect 18693 5729 18705 5763
rect 18739 5760 18751 5763
rect 18739 5732 18920 5760
rect 18739 5729 18751 5732
rect 18693 5723 18751 5729
rect 15933 5695 15991 5701
rect 15933 5692 15945 5695
rect 15160 5664 15945 5692
rect 15160 5652 15166 5664
rect 15933 5661 15945 5664
rect 15979 5661 15991 5695
rect 15933 5655 15991 5661
rect 18509 5695 18567 5701
rect 18509 5661 18521 5695
rect 18555 5692 18567 5695
rect 18782 5692 18788 5704
rect 18555 5664 18788 5692
rect 18555 5661 18567 5664
rect 18509 5655 18567 5661
rect 18782 5652 18788 5664
rect 18840 5652 18846 5704
rect 11054 5584 11060 5636
rect 11112 5584 11118 5636
rect 13446 5584 13452 5636
rect 13504 5624 13510 5636
rect 16209 5627 16267 5633
rect 13504 5596 15148 5624
rect 13504 5584 13510 5596
rect 15120 5565 15148 5596
rect 16209 5593 16221 5627
rect 16255 5593 16267 5627
rect 16209 5587 16267 5593
rect 15105 5559 15163 5565
rect 15105 5525 15117 5559
rect 15151 5525 15163 5559
rect 16224 5556 16252 5587
rect 16666 5584 16672 5636
rect 16724 5584 16730 5636
rect 16850 5556 16856 5568
rect 16224 5528 16856 5556
rect 15105 5519 15163 5525
rect 16850 5516 16856 5528
rect 16908 5556 16914 5568
rect 18892 5556 18920 5732
rect 19886 5720 19892 5772
rect 19944 5720 19950 5772
rect 19613 5695 19671 5701
rect 19613 5661 19625 5695
rect 19659 5692 19671 5695
rect 19659 5664 20208 5692
rect 19659 5661 19671 5664
rect 19613 5655 19671 5661
rect 16908 5528 18920 5556
rect 20180 5556 20208 5664
rect 20548 5624 20576 5800
rect 22002 5788 22008 5840
rect 22060 5828 22066 5840
rect 24857 5831 24915 5837
rect 24857 5828 24869 5831
rect 22060 5800 24869 5828
rect 22060 5788 22066 5800
rect 24857 5797 24869 5800
rect 24903 5797 24915 5831
rect 24857 5791 24915 5797
rect 21729 5763 21787 5769
rect 21729 5760 21741 5763
rect 20640 5732 21741 5760
rect 20640 5704 20668 5732
rect 21729 5729 21741 5732
rect 21775 5729 21787 5763
rect 21729 5723 21787 5729
rect 20622 5652 20628 5704
rect 20680 5652 20686 5704
rect 21450 5652 21456 5704
rect 21508 5652 21514 5704
rect 22738 5652 22744 5704
rect 22796 5692 22802 5704
rect 23201 5695 23259 5701
rect 23201 5692 23213 5695
rect 22796 5664 23213 5692
rect 22796 5652 22802 5664
rect 23201 5661 23213 5664
rect 23247 5692 23259 5695
rect 23842 5692 23848 5704
rect 23247 5664 23848 5692
rect 23247 5661 23259 5664
rect 23201 5655 23259 5661
rect 23842 5652 23848 5664
rect 23900 5652 23906 5704
rect 23934 5652 23940 5704
rect 23992 5692 23998 5704
rect 24029 5695 24087 5701
rect 24029 5692 24041 5695
rect 23992 5664 24041 5692
rect 23992 5652 23998 5664
rect 24029 5661 24041 5664
rect 24075 5661 24087 5695
rect 24029 5655 24087 5661
rect 24578 5652 24584 5704
rect 24636 5692 24642 5704
rect 24673 5695 24731 5701
rect 24673 5692 24685 5695
rect 24636 5664 24685 5692
rect 24636 5652 24642 5664
rect 24673 5661 24685 5664
rect 24719 5661 24731 5695
rect 24673 5655 24731 5661
rect 23385 5627 23443 5633
rect 20548 5596 22094 5624
rect 20898 5556 20904 5568
rect 20180 5528 20904 5556
rect 16908 5516 16914 5528
rect 20898 5516 20904 5528
rect 20956 5516 20962 5568
rect 22066 5556 22094 5596
rect 23385 5593 23397 5627
rect 23431 5624 23443 5627
rect 23750 5624 23756 5636
rect 23431 5596 23756 5624
rect 23431 5593 23443 5596
rect 23385 5587 23443 5593
rect 23750 5584 23756 5596
rect 23808 5584 23814 5636
rect 25130 5624 25136 5636
rect 23860 5596 25136 5624
rect 23860 5556 23888 5596
rect 25130 5584 25136 5596
rect 25188 5584 25194 5636
rect 22066 5528 23888 5556
rect 24578 5516 24584 5568
rect 24636 5556 24642 5568
rect 25317 5559 25375 5565
rect 25317 5556 25329 5559
rect 24636 5528 25329 5556
rect 24636 5516 24642 5528
rect 25317 5525 25329 5528
rect 25363 5525 25375 5559
rect 25317 5519 25375 5525
rect 1104 5466 25852 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 25852 5466
rect 1104 5392 25852 5414
rect 3418 5312 3424 5364
rect 3476 5352 3482 5364
rect 10686 5352 10692 5364
rect 3476 5324 10692 5352
rect 3476 5312 3482 5324
rect 10686 5312 10692 5324
rect 10744 5312 10750 5364
rect 10965 5355 11023 5361
rect 10965 5321 10977 5355
rect 11011 5352 11023 5355
rect 11606 5352 11612 5364
rect 11011 5324 11612 5352
rect 11011 5321 11023 5324
rect 10965 5315 11023 5321
rect 11606 5312 11612 5324
rect 11664 5312 11670 5364
rect 13630 5352 13636 5364
rect 13464 5324 13636 5352
rect 11054 5244 11060 5296
rect 11112 5284 11118 5296
rect 11514 5284 11520 5296
rect 11112 5256 11520 5284
rect 11112 5244 11118 5256
rect 11514 5244 11520 5256
rect 11572 5244 11578 5296
rect 11698 5244 11704 5296
rect 11756 5284 11762 5296
rect 13464 5293 13492 5324
rect 13630 5312 13636 5324
rect 13688 5312 13694 5364
rect 14182 5312 14188 5364
rect 14240 5352 14246 5364
rect 14921 5355 14979 5361
rect 14921 5352 14933 5355
rect 14240 5324 14933 5352
rect 14240 5312 14246 5324
rect 14921 5321 14933 5324
rect 14967 5352 14979 5355
rect 17310 5352 17316 5364
rect 14967 5324 17316 5352
rect 14967 5321 14979 5324
rect 14921 5315 14979 5321
rect 17310 5312 17316 5324
rect 17368 5312 17374 5364
rect 18432 5324 20392 5352
rect 13449 5287 13507 5293
rect 11756 5256 12572 5284
rect 11756 5244 11762 5256
rect 10689 5219 10747 5225
rect 10689 5185 10701 5219
rect 10735 5216 10747 5219
rect 11149 5219 11207 5225
rect 11149 5216 11161 5219
rect 10735 5188 11161 5216
rect 10735 5185 10747 5188
rect 10689 5179 10747 5185
rect 11149 5185 11161 5188
rect 11195 5216 11207 5219
rect 11422 5216 11428 5228
rect 11195 5188 11428 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 11422 5176 11428 5188
rect 11480 5176 11486 5228
rect 12544 5216 12572 5256
rect 13449 5253 13461 5287
rect 13495 5253 13507 5287
rect 13449 5247 13507 5253
rect 14458 5244 14464 5296
rect 14516 5244 14522 5296
rect 17862 5244 17868 5296
rect 17920 5244 17926 5296
rect 13173 5219 13231 5225
rect 13173 5216 13185 5219
rect 12544 5188 13185 5216
rect 11793 5151 11851 5157
rect 11793 5117 11805 5151
rect 11839 5148 11851 5151
rect 11882 5148 11888 5160
rect 11839 5120 11888 5148
rect 11839 5117 11851 5120
rect 11793 5111 11851 5117
rect 11882 5108 11888 5120
rect 11940 5108 11946 5160
rect 12066 5108 12072 5160
rect 12124 5148 12130 5160
rect 12161 5151 12219 5157
rect 12161 5148 12173 5151
rect 12124 5120 12173 5148
rect 12124 5108 12130 5120
rect 12161 5117 12173 5120
rect 12207 5117 12219 5151
rect 12161 5111 12219 5117
rect 12544 5012 12572 5188
rect 13173 5185 13185 5188
rect 13219 5185 13231 5219
rect 13173 5179 13231 5185
rect 17129 5219 17187 5225
rect 17129 5185 17141 5219
rect 17175 5216 17187 5219
rect 18432 5216 18460 5324
rect 17175 5188 18460 5216
rect 17175 5185 17187 5188
rect 17129 5179 17187 5185
rect 18506 5176 18512 5228
rect 18564 5216 18570 5228
rect 18785 5219 18843 5225
rect 18785 5216 18797 5219
rect 18564 5188 18797 5216
rect 18564 5176 18570 5188
rect 18785 5185 18797 5188
rect 18831 5185 18843 5219
rect 18785 5179 18843 5185
rect 20162 5176 20168 5228
rect 20220 5176 20226 5228
rect 20364 5216 20392 5324
rect 20438 5312 20444 5364
rect 20496 5352 20502 5364
rect 20533 5355 20591 5361
rect 20533 5352 20545 5355
rect 20496 5324 20545 5352
rect 20496 5312 20502 5324
rect 20533 5321 20545 5324
rect 20579 5321 20591 5355
rect 21910 5352 21916 5364
rect 20533 5315 20591 5321
rect 20640 5324 21916 5352
rect 20640 5216 20668 5324
rect 21910 5312 21916 5324
rect 21968 5312 21974 5364
rect 20806 5244 20812 5296
rect 20864 5284 20870 5296
rect 20864 5256 21220 5284
rect 20864 5244 20870 5256
rect 20364 5188 20668 5216
rect 21082 5176 21088 5228
rect 21140 5176 21146 5228
rect 21192 5216 21220 5256
rect 21542 5244 21548 5296
rect 21600 5244 21606 5296
rect 22002 5216 22008 5228
rect 21192 5188 22008 5216
rect 22002 5176 22008 5188
rect 22060 5176 22066 5228
rect 22094 5176 22100 5228
rect 22152 5176 22158 5228
rect 23750 5176 23756 5228
rect 23808 5216 23814 5228
rect 23845 5219 23903 5225
rect 23845 5216 23857 5219
rect 23808 5188 23857 5216
rect 23808 5176 23814 5188
rect 23845 5185 23857 5188
rect 23891 5185 23903 5219
rect 23845 5179 23903 5185
rect 15194 5108 15200 5160
rect 15252 5148 15258 5160
rect 15473 5151 15531 5157
rect 15473 5148 15485 5151
rect 15252 5120 15485 5148
rect 15252 5108 15258 5120
rect 15473 5117 15485 5120
rect 15519 5117 15531 5151
rect 15473 5111 15531 5117
rect 15746 5108 15752 5160
rect 15804 5108 15810 5160
rect 19061 5151 19119 5157
rect 19061 5117 19073 5151
rect 19107 5148 19119 5151
rect 21266 5148 21272 5160
rect 19107 5120 21272 5148
rect 19107 5117 19119 5120
rect 19061 5111 19119 5117
rect 21266 5108 21272 5120
rect 21324 5108 21330 5160
rect 21542 5108 21548 5160
rect 21600 5148 21606 5160
rect 22465 5151 22523 5157
rect 22465 5148 22477 5151
rect 21600 5120 22477 5148
rect 21600 5108 21606 5120
rect 22465 5117 22477 5120
rect 22511 5117 22523 5151
rect 22465 5111 22523 5117
rect 23474 5108 23480 5160
rect 23532 5148 23538 5160
rect 24305 5151 24363 5157
rect 24305 5148 24317 5151
rect 23532 5120 24317 5148
rect 23532 5108 23538 5120
rect 24305 5117 24317 5120
rect 24351 5117 24363 5151
rect 24305 5111 24363 5117
rect 14918 5040 14924 5092
rect 14976 5080 14982 5092
rect 18414 5080 18420 5092
rect 14976 5052 18420 5080
rect 14976 5040 14982 5052
rect 18414 5040 18420 5052
rect 18472 5040 18478 5092
rect 20162 5040 20168 5092
rect 20220 5080 20226 5092
rect 24210 5080 24216 5092
rect 20220 5052 24216 5080
rect 20220 5040 20226 5052
rect 24210 5040 24216 5052
rect 24268 5040 24274 5092
rect 13906 5012 13912 5024
rect 12544 4984 13912 5012
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 15470 4972 15476 5024
rect 15528 5012 15534 5024
rect 21177 5015 21235 5021
rect 21177 5012 21189 5015
rect 15528 4984 21189 5012
rect 15528 4972 15534 4984
rect 21177 4981 21189 4984
rect 21223 4981 21235 5015
rect 21177 4975 21235 4981
rect 1104 4922 25852 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 25852 4922
rect 1104 4848 25852 4870
rect 10134 4768 10140 4820
rect 10192 4768 10198 4820
rect 11238 4768 11244 4820
rect 11296 4808 11302 4820
rect 11422 4808 11428 4820
rect 11296 4780 11428 4808
rect 11296 4768 11302 4780
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 11882 4768 11888 4820
rect 11940 4808 11946 4820
rect 20162 4808 20168 4820
rect 11940 4780 20168 4808
rect 11940 4768 11946 4780
rect 20162 4768 20168 4780
rect 20220 4768 20226 4820
rect 21266 4768 21272 4820
rect 21324 4768 21330 4820
rect 22370 4768 22376 4820
rect 22428 4808 22434 4820
rect 24765 4811 24823 4817
rect 24765 4808 24777 4811
rect 22428 4780 24777 4808
rect 22428 4768 22434 4780
rect 24765 4777 24777 4780
rect 24811 4777 24823 4811
rect 24765 4771 24823 4777
rect 10413 4743 10471 4749
rect 10413 4709 10425 4743
rect 10459 4740 10471 4743
rect 10459 4712 15240 4740
rect 10459 4709 10471 4712
rect 10413 4703 10471 4709
rect 1486 4632 1492 4684
rect 1544 4672 1550 4684
rect 2041 4675 2099 4681
rect 2041 4672 2053 4675
rect 1544 4644 2053 4672
rect 1544 4632 1550 4644
rect 2041 4641 2053 4644
rect 2087 4641 2099 4675
rect 2041 4635 2099 4641
rect 5077 4675 5135 4681
rect 5077 4641 5089 4675
rect 5123 4672 5135 4675
rect 9582 4672 9588 4684
rect 5123 4644 9588 4672
rect 5123 4641 5135 4644
rect 5077 4635 5135 4641
rect 9582 4632 9588 4644
rect 9640 4632 9646 4684
rect 11238 4672 11244 4684
rect 10612 4644 11244 4672
rect 1762 4564 1768 4616
rect 1820 4564 1826 4616
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 3988 4536 4016 4567
rect 7098 4564 7104 4616
rect 7156 4564 7162 4616
rect 10612 4613 10640 4644
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 11333 4675 11391 4681
rect 11333 4641 11345 4675
rect 11379 4672 11391 4675
rect 14918 4672 14924 4684
rect 11379 4644 14924 4672
rect 11379 4641 11391 4644
rect 11333 4635 11391 4641
rect 14918 4632 14924 4644
rect 14976 4632 14982 4684
rect 15102 4632 15108 4684
rect 15160 4632 15166 4684
rect 15212 4672 15240 4712
rect 16850 4700 16856 4752
rect 16908 4700 16914 4752
rect 16960 4712 19656 4740
rect 15470 4672 15476 4684
rect 15212 4644 15476 4672
rect 15470 4632 15476 4644
rect 15528 4632 15534 4684
rect 15838 4632 15844 4684
rect 15896 4672 15902 4684
rect 16960 4672 16988 4712
rect 15896 4644 16988 4672
rect 15896 4632 15902 4644
rect 18506 4632 18512 4684
rect 18564 4672 18570 4684
rect 19521 4675 19579 4681
rect 19521 4672 19533 4675
rect 18564 4644 19533 4672
rect 18564 4632 18570 4644
rect 19521 4641 19533 4644
rect 19567 4641 19579 4675
rect 19628 4672 19656 4712
rect 22066 4712 23704 4740
rect 22066 4672 22094 4712
rect 19628 4644 22094 4672
rect 19521 4635 19579 4641
rect 9861 4607 9919 4613
rect 9861 4573 9873 4607
rect 9907 4604 9919 4607
rect 10597 4607 10655 4613
rect 10597 4604 10609 4607
rect 9907 4576 10609 4604
rect 9907 4573 9919 4576
rect 9861 4567 9919 4573
rect 10597 4573 10609 4576
rect 10643 4573 10655 4607
rect 10597 4567 10655 4573
rect 11057 4607 11115 4613
rect 11057 4573 11069 4607
rect 11103 4573 11115 4607
rect 11057 4567 11115 4573
rect 12529 4607 12587 4613
rect 12529 4573 12541 4607
rect 12575 4604 12587 4607
rect 14274 4604 14280 4616
rect 12575 4576 14280 4604
rect 12575 4573 12587 4576
rect 12529 4567 12587 4573
rect 1596 4508 4016 4536
rect 4617 4539 4675 4545
rect 1596 4477 1624 4508
rect 4617 4505 4629 4539
rect 4663 4536 4675 4539
rect 5353 4539 5411 4545
rect 5353 4536 5365 4539
rect 4663 4508 5365 4536
rect 4663 4505 4675 4508
rect 4617 4499 4675 4505
rect 5353 4505 5365 4508
rect 5399 4505 5411 4539
rect 7377 4539 7435 4545
rect 7377 4536 7389 4539
rect 6578 4508 7389 4536
rect 5353 4499 5411 4505
rect 7377 4505 7389 4508
rect 7423 4505 7435 4539
rect 7377 4499 7435 4505
rect 9769 4539 9827 4545
rect 9769 4505 9781 4539
rect 9815 4536 9827 4539
rect 10686 4536 10692 4548
rect 9815 4508 10692 4536
rect 9815 4505 9827 4508
rect 9769 4499 9827 4505
rect 1581 4471 1639 4477
rect 1581 4437 1593 4471
rect 1627 4437 1639 4471
rect 7392 4468 7420 4499
rect 10686 4496 10692 4508
rect 10744 4496 10750 4548
rect 11072 4536 11100 4567
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14461 4607 14519 4613
rect 14461 4573 14473 4607
rect 14507 4604 14519 4607
rect 14734 4604 14740 4616
rect 14507 4576 14740 4604
rect 14507 4573 14519 4576
rect 14461 4567 14519 4573
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 17589 4607 17647 4613
rect 17589 4573 17601 4607
rect 17635 4604 17647 4607
rect 17635 4576 18552 4604
rect 17635 4573 17647 4576
rect 17589 4567 17647 4573
rect 13541 4539 13599 4545
rect 11072 4508 12434 4536
rect 11054 4468 11060 4480
rect 7392 4440 11060 4468
rect 1581 4431 1639 4437
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 12406 4468 12434 4508
rect 13541 4505 13553 4539
rect 13587 4536 13599 4539
rect 14918 4536 14924 4548
rect 13587 4508 14924 4536
rect 13587 4505 13599 4508
rect 13541 4499 13599 4505
rect 14918 4496 14924 4508
rect 14976 4496 14982 4548
rect 15378 4496 15384 4548
rect 15436 4496 15442 4548
rect 15838 4536 15844 4548
rect 15764 4508 15844 4536
rect 13446 4468 13452 4480
rect 12406 4440 13452 4468
rect 13446 4428 13452 4440
rect 13504 4428 13510 4480
rect 14277 4471 14335 4477
rect 14277 4437 14289 4471
rect 14323 4468 14335 4471
rect 14458 4468 14464 4480
rect 14323 4440 14464 4468
rect 14323 4437 14335 4440
rect 14277 4431 14335 4437
rect 14458 4428 14464 4440
rect 14516 4428 14522 4480
rect 14550 4428 14556 4480
rect 14608 4468 14614 4480
rect 14737 4471 14795 4477
rect 14737 4468 14749 4471
rect 14608 4440 14749 4468
rect 14608 4428 14614 4440
rect 14737 4437 14749 4440
rect 14783 4468 14795 4471
rect 15764 4468 15792 4508
rect 15838 4496 15844 4508
rect 15896 4496 15902 4548
rect 18322 4496 18328 4548
rect 18380 4496 18386 4548
rect 18524 4536 18552 4576
rect 21818 4564 21824 4616
rect 21876 4564 21882 4616
rect 22002 4564 22008 4616
rect 22060 4604 22066 4616
rect 23676 4613 23704 4712
rect 24026 4700 24032 4752
rect 24084 4740 24090 4752
rect 25317 4743 25375 4749
rect 25317 4740 25329 4743
rect 24084 4712 25329 4740
rect 24084 4700 24090 4712
rect 25317 4709 25329 4712
rect 25363 4709 25375 4743
rect 25317 4703 25375 4709
rect 23661 4607 23719 4613
rect 22060 4576 23612 4604
rect 22060 4564 22066 4576
rect 19702 4536 19708 4548
rect 18524 4508 19708 4536
rect 19702 4496 19708 4508
rect 19760 4496 19766 4548
rect 19794 4496 19800 4548
rect 19852 4496 19858 4548
rect 20254 4496 20260 4548
rect 20312 4496 20318 4548
rect 22649 4539 22707 4545
rect 22649 4505 22661 4539
rect 22695 4505 22707 4539
rect 23584 4536 23612 4576
rect 23661 4573 23673 4607
rect 23707 4604 23719 4607
rect 24121 4607 24179 4613
rect 24121 4604 24133 4607
rect 23707 4576 24133 4604
rect 23707 4573 23719 4576
rect 23661 4567 23719 4573
rect 24121 4573 24133 4576
rect 24167 4573 24179 4607
rect 24121 4567 24179 4573
rect 24673 4539 24731 4545
rect 24673 4536 24685 4539
rect 23584 4508 24685 4536
rect 22649 4499 22707 4505
rect 24673 4505 24685 4508
rect 24719 4536 24731 4539
rect 25133 4539 25191 4545
rect 25133 4536 25145 4539
rect 24719 4508 25145 4536
rect 24719 4505 24731 4508
rect 24673 4499 24731 4505
rect 25133 4505 25145 4508
rect 25179 4505 25191 4539
rect 25133 4499 25191 4505
rect 16666 4468 16672 4480
rect 14783 4440 16672 4468
rect 14783 4437 14795 4440
rect 14737 4431 14795 4437
rect 16666 4428 16672 4440
rect 16724 4428 16730 4480
rect 19978 4428 19984 4480
rect 20036 4468 20042 4480
rect 22664 4468 22692 4499
rect 20036 4440 22692 4468
rect 20036 4428 20042 4440
rect 23750 4428 23756 4480
rect 23808 4428 23814 4480
rect 1104 4378 25852 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 25852 4378
rect 1104 4304 25852 4326
rect 1762 4224 1768 4276
rect 1820 4264 1826 4276
rect 2225 4267 2283 4273
rect 2225 4264 2237 4267
rect 1820 4236 2237 4264
rect 1820 4224 1826 4236
rect 2225 4233 2237 4236
rect 2271 4233 2283 4267
rect 2225 4227 2283 4233
rect 14550 4224 14556 4276
rect 14608 4224 14614 4276
rect 15470 4224 15476 4276
rect 15528 4264 15534 4276
rect 15657 4267 15715 4273
rect 15657 4264 15669 4267
rect 15528 4236 15669 4264
rect 15528 4224 15534 4236
rect 15657 4233 15669 4236
rect 15703 4233 15715 4267
rect 15657 4227 15715 4233
rect 16117 4267 16175 4273
rect 16117 4233 16129 4267
rect 16163 4264 16175 4267
rect 17218 4264 17224 4276
rect 16163 4236 17224 4264
rect 16163 4233 16175 4236
rect 16117 4227 16175 4233
rect 17218 4224 17224 4236
rect 17276 4224 17282 4276
rect 20254 4224 20260 4276
rect 20312 4264 20318 4276
rect 21545 4267 21603 4273
rect 21545 4264 21557 4267
rect 20312 4236 21557 4264
rect 20312 4224 20318 4236
rect 21545 4233 21557 4236
rect 21591 4264 21603 4267
rect 22005 4267 22063 4273
rect 22005 4264 22017 4267
rect 21591 4236 22017 4264
rect 21591 4233 21603 4236
rect 21545 4227 21603 4233
rect 22005 4233 22017 4236
rect 22051 4233 22063 4267
rect 22005 4227 22063 4233
rect 24670 4224 24676 4276
rect 24728 4224 24734 4276
rect 12176 4168 12388 4196
rect 1486 4088 1492 4140
rect 1544 4128 1550 4140
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 1544 4100 1593 4128
rect 1544 4088 1550 4100
rect 1581 4097 1593 4100
rect 1627 4097 1639 4131
rect 1581 4091 1639 4097
rect 1854 4088 1860 4140
rect 1912 4128 1918 4140
rect 2869 4131 2927 4137
rect 2869 4128 2881 4131
rect 1912 4100 2881 4128
rect 1912 4088 1918 4100
rect 2869 4097 2881 4100
rect 2915 4128 2927 4131
rect 3145 4131 3203 4137
rect 3145 4128 3157 4131
rect 2915 4100 3157 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 3145 4097 3157 4100
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 4341 4131 4399 4137
rect 4341 4128 4353 4131
rect 4120 4100 4353 4128
rect 4120 4088 4126 4100
rect 4341 4097 4353 4100
rect 4387 4097 4399 4131
rect 4341 4091 4399 4097
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 9493 4131 9551 4137
rect 9493 4128 9505 4131
rect 9272 4100 9505 4128
rect 9272 4088 9278 4100
rect 9493 4097 9505 4100
rect 9539 4097 9551 4131
rect 9493 4091 9551 4097
rect 10244 4100 10548 4128
rect 10244 4060 10272 4100
rect 9324 4032 10272 4060
rect 2682 3952 2688 4004
rect 2740 3952 2746 4004
rect 4157 3995 4215 4001
rect 4157 3961 4169 3995
rect 4203 3992 4215 3995
rect 7282 3992 7288 4004
rect 4203 3964 7288 3992
rect 4203 3961 4215 3964
rect 4157 3955 4215 3961
rect 7282 3952 7288 3964
rect 7340 3952 7346 4004
rect 9324 4001 9352 4032
rect 10318 4020 10324 4072
rect 10376 4020 10382 4072
rect 10520 4060 10548 4100
rect 10594 4088 10600 4140
rect 10652 4088 10658 4140
rect 12176 4128 12204 4168
rect 11532 4100 12204 4128
rect 11532 4060 11560 4100
rect 12250 4088 12256 4140
rect 12308 4088 12314 4140
rect 12360 4128 12388 4168
rect 14182 4156 14188 4208
rect 14240 4156 14246 4208
rect 14568 4196 14596 4224
rect 14568 4168 14674 4196
rect 15562 4156 15568 4208
rect 15620 4196 15626 4208
rect 22465 4199 22523 4205
rect 22465 4196 22477 4199
rect 15620 4168 22477 4196
rect 15620 4156 15626 4168
rect 22465 4165 22477 4168
rect 22511 4165 22523 4199
rect 22465 4159 22523 4165
rect 13354 4128 13360 4140
rect 12360 4100 13360 4128
rect 13354 4088 13360 4100
rect 13412 4088 13418 4140
rect 13906 4088 13912 4140
rect 13964 4088 13970 4140
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 17083 4100 17724 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 10520 4032 11560 4060
rect 11609 4063 11667 4069
rect 11609 4029 11621 4063
rect 11655 4060 11667 4063
rect 12618 4060 12624 4072
rect 11655 4032 12624 4060
rect 11655 4029 11667 4032
rect 11609 4023 11667 4029
rect 12618 4020 12624 4032
rect 12676 4020 12682 4072
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4029 13323 4063
rect 13265 4023 13323 4029
rect 9309 3995 9367 4001
rect 9309 3961 9321 3995
rect 9355 3961 9367 3995
rect 9309 3955 9367 3961
rect 9861 3995 9919 4001
rect 9861 3961 9873 3995
rect 9907 3992 9919 3995
rect 11698 3992 11704 4004
rect 9907 3964 11704 3992
rect 9907 3961 9919 3964
rect 9861 3955 9919 3961
rect 11698 3952 11704 3964
rect 11756 3952 11762 4004
rect 3881 3927 3939 3933
rect 3881 3893 3893 3927
rect 3927 3924 3939 3927
rect 4062 3924 4068 3936
rect 3927 3896 4068 3924
rect 3927 3893 3939 3896
rect 3881 3887 3939 3893
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 4798 3884 4804 3936
rect 4856 3884 4862 3936
rect 5258 3884 5264 3936
rect 5316 3924 5322 3936
rect 6089 3927 6147 3933
rect 6089 3924 6101 3927
rect 5316 3896 6101 3924
rect 5316 3884 5322 3896
rect 6089 3893 6101 3896
rect 6135 3893 6147 3927
rect 6089 3887 6147 3893
rect 7006 3884 7012 3936
rect 7064 3884 7070 3936
rect 9033 3927 9091 3933
rect 9033 3893 9045 3927
rect 9079 3924 9091 3927
rect 9214 3924 9220 3936
rect 9079 3896 9220 3924
rect 9079 3893 9091 3896
rect 9033 3887 9091 3893
rect 9214 3884 9220 3896
rect 9272 3884 9278 3936
rect 10042 3884 10048 3936
rect 10100 3884 10106 3936
rect 11793 3927 11851 3933
rect 11793 3893 11805 3927
rect 11839 3924 11851 3927
rect 12158 3924 12164 3936
rect 11839 3896 12164 3924
rect 11839 3893 11851 3896
rect 11793 3887 11851 3893
rect 12158 3884 12164 3896
rect 12216 3884 12222 3936
rect 13280 3924 13308 4023
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 17313 4063 17371 4069
rect 17313 4060 17325 4063
rect 16264 4032 17325 4060
rect 16264 4020 16270 4032
rect 17313 4029 17325 4032
rect 17359 4029 17371 4063
rect 17313 4023 17371 4029
rect 17696 3992 17724 4100
rect 17770 4088 17776 4140
rect 17828 4128 17834 4140
rect 18693 4131 18751 4137
rect 18693 4128 18705 4131
rect 17828 4100 18705 4128
rect 17828 4088 17834 4100
rect 18693 4097 18705 4100
rect 18739 4097 18751 4131
rect 18693 4091 18751 4097
rect 20898 4088 20904 4140
rect 20956 4088 20962 4140
rect 20990 4088 20996 4140
rect 21048 4088 21054 4140
rect 21818 4088 21824 4140
rect 21876 4088 21882 4140
rect 22002 4088 22008 4140
rect 22060 4128 22066 4140
rect 25133 4131 25191 4137
rect 25133 4128 25145 4131
rect 22060 4100 25145 4128
rect 22060 4088 22066 4100
rect 25133 4097 25145 4100
rect 25179 4097 25191 4131
rect 25133 4091 25191 4097
rect 18414 4020 18420 4072
rect 18472 4060 18478 4072
rect 19153 4063 19211 4069
rect 19153 4060 19165 4063
rect 18472 4032 19165 4060
rect 18472 4020 18478 4032
rect 19153 4029 19165 4032
rect 19199 4029 19211 4063
rect 19153 4023 19211 4029
rect 21177 4063 21235 4069
rect 21177 4029 21189 4063
rect 21223 4060 21235 4063
rect 21266 4060 21272 4072
rect 21223 4032 21272 4060
rect 21223 4029 21235 4032
rect 21177 4023 21235 4029
rect 21266 4020 21272 4032
rect 21324 4020 21330 4072
rect 21910 4020 21916 4072
rect 21968 4020 21974 4072
rect 24118 4020 24124 4072
rect 24176 4020 24182 4072
rect 19058 3992 19064 4004
rect 17696 3964 19064 3992
rect 19058 3952 19064 3964
rect 19116 3952 19122 4004
rect 21928 3992 21956 4020
rect 22554 3992 22560 4004
rect 21928 3964 22560 3992
rect 22554 3952 22560 3964
rect 22612 3952 22618 4004
rect 17494 3924 17500 3936
rect 13280 3896 17500 3924
rect 17494 3884 17500 3896
rect 17552 3884 17558 3936
rect 19150 3884 19156 3936
rect 19208 3924 19214 3936
rect 19886 3924 19892 3936
rect 19208 3896 19892 3924
rect 19208 3884 19214 3896
rect 19886 3884 19892 3896
rect 19944 3884 19950 3936
rect 20533 3927 20591 3933
rect 20533 3893 20545 3927
rect 20579 3924 20591 3927
rect 21450 3924 21456 3936
rect 20579 3896 21456 3924
rect 20579 3893 20591 3896
rect 20533 3887 20591 3893
rect 21450 3884 21456 3896
rect 21508 3884 21514 3936
rect 21910 3884 21916 3936
rect 21968 3924 21974 3936
rect 22094 3924 22100 3936
rect 21968 3896 22100 3924
rect 21968 3884 21974 3896
rect 22094 3884 22100 3896
rect 22152 3884 22158 3936
rect 23750 3884 23756 3936
rect 23808 3924 23814 3936
rect 25317 3927 25375 3933
rect 25317 3924 25329 3927
rect 23808 3896 25329 3924
rect 23808 3884 23814 3896
rect 25317 3893 25329 3896
rect 25363 3893 25375 3927
rect 25317 3887 25375 3893
rect 1104 3834 25852 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 25852 3834
rect 1104 3760 25852 3782
rect 2869 3723 2927 3729
rect 2869 3689 2881 3723
rect 2915 3720 2927 3723
rect 3326 3720 3332 3732
rect 2915 3692 3332 3720
rect 2915 3689 2927 3692
rect 2869 3683 2927 3689
rect 3326 3680 3332 3692
rect 3384 3680 3390 3732
rect 4249 3723 4307 3729
rect 4249 3689 4261 3723
rect 4295 3720 4307 3723
rect 7834 3720 7840 3732
rect 4295 3692 7840 3720
rect 4295 3689 4307 3692
rect 4249 3683 4307 3689
rect 7834 3680 7840 3692
rect 7892 3680 7898 3732
rect 8386 3680 8392 3732
rect 8444 3680 8450 3732
rect 10413 3723 10471 3729
rect 10413 3689 10425 3723
rect 10459 3720 10471 3723
rect 10502 3720 10508 3732
rect 10459 3692 10508 3720
rect 10459 3689 10471 3692
rect 10413 3683 10471 3689
rect 10502 3680 10508 3692
rect 10560 3680 10566 3732
rect 13814 3720 13820 3732
rect 13556 3692 13820 3720
rect 1872 3624 5304 3652
rect 1872 3593 1900 3624
rect 1857 3587 1915 3593
rect 1857 3553 1869 3587
rect 1903 3553 1915 3587
rect 1857 3547 1915 3553
rect 5166 3544 5172 3596
rect 5224 3544 5230 3596
rect 5276 3584 5304 3624
rect 6362 3612 6368 3664
rect 6420 3612 6426 3664
rect 7101 3655 7159 3661
rect 7101 3621 7113 3655
rect 7147 3652 7159 3655
rect 8846 3652 8852 3664
rect 7147 3624 8852 3652
rect 7147 3621 7159 3624
rect 7101 3615 7159 3621
rect 8846 3612 8852 3624
rect 8904 3612 8910 3664
rect 9677 3655 9735 3661
rect 9677 3621 9689 3655
rect 9723 3652 9735 3655
rect 13556 3652 13584 3692
rect 13814 3680 13820 3692
rect 13872 3680 13878 3732
rect 14918 3680 14924 3732
rect 14976 3720 14982 3732
rect 18506 3720 18512 3732
rect 14976 3692 18512 3720
rect 14976 3680 14982 3692
rect 18506 3680 18512 3692
rect 18564 3680 18570 3732
rect 20254 3680 20260 3732
rect 20312 3720 20318 3732
rect 21542 3720 21548 3732
rect 20312 3692 21548 3720
rect 20312 3680 20318 3692
rect 21542 3680 21548 3692
rect 21600 3680 21606 3732
rect 22646 3680 22652 3732
rect 22704 3720 22710 3732
rect 23845 3723 23903 3729
rect 23845 3720 23857 3723
rect 22704 3692 23857 3720
rect 22704 3680 22710 3692
rect 23845 3689 23857 3692
rect 23891 3689 23903 3723
rect 23845 3683 23903 3689
rect 14366 3652 14372 3664
rect 9723 3624 13584 3652
rect 13648 3624 14372 3652
rect 9723 3621 9735 3624
rect 9677 3615 9735 3621
rect 8386 3584 8392 3596
rect 5276 3556 8392 3584
rect 8386 3544 8392 3556
rect 8444 3544 8450 3596
rect 10042 3544 10048 3596
rect 10100 3584 10106 3596
rect 11057 3587 11115 3593
rect 11057 3584 11069 3587
rect 10100 3556 11069 3584
rect 10100 3544 10106 3556
rect 11057 3553 11069 3556
rect 11103 3584 11115 3587
rect 12526 3584 12532 3596
rect 11103 3556 12532 3584
rect 11103 3553 11115 3556
rect 11057 3547 11115 3553
rect 12526 3544 12532 3556
rect 12584 3544 12590 3596
rect 12802 3544 12808 3596
rect 12860 3544 12866 3596
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3485 1639 3519
rect 1581 3479 1639 3485
rect 1596 3448 1624 3479
rect 2222 3476 2228 3528
rect 2280 3516 2286 3528
rect 3053 3519 3111 3525
rect 3053 3516 3065 3519
rect 2280 3488 3065 3516
rect 2280 3476 2286 3488
rect 3053 3485 3065 3488
rect 3099 3516 3111 3519
rect 3513 3519 3571 3525
rect 3513 3516 3525 3519
rect 3099 3488 3525 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 3513 3485 3525 3488
rect 3559 3485 3571 3519
rect 3513 3479 3571 3485
rect 4430 3476 4436 3528
rect 4488 3476 4494 3528
rect 4798 3476 4804 3528
rect 4856 3516 4862 3528
rect 4893 3519 4951 3525
rect 4893 3516 4905 3519
rect 4856 3488 4905 3516
rect 4856 3476 4862 3488
rect 4893 3485 4905 3488
rect 4939 3485 4951 3519
rect 6549 3519 6607 3525
rect 6549 3516 6561 3519
rect 4893 3479 4951 3485
rect 6288 3488 6561 3516
rect 1596 3420 3832 3448
rect 3804 3392 3832 3420
rect 6288 3392 6316 3488
rect 6549 3485 6561 3488
rect 6595 3485 6607 3519
rect 6549 3479 6607 3485
rect 7006 3476 7012 3528
rect 7064 3516 7070 3528
rect 7285 3519 7343 3525
rect 7285 3516 7297 3519
rect 7064 3488 7297 3516
rect 7064 3476 7070 3488
rect 7285 3485 7297 3488
rect 7331 3485 7343 3519
rect 7285 3479 7343 3485
rect 8478 3476 8484 3528
rect 8536 3516 8542 3528
rect 8573 3519 8631 3525
rect 8573 3516 8585 3519
rect 8536 3488 8585 3516
rect 8536 3476 8542 3488
rect 8573 3485 8585 3488
rect 8619 3516 8631 3519
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8619 3488 8953 3516
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 9861 3519 9919 3525
rect 9861 3516 9873 3519
rect 8941 3479 8999 3485
rect 9600 3488 9873 3516
rect 7374 3408 7380 3460
rect 7432 3448 7438 3460
rect 7837 3451 7895 3457
rect 7837 3448 7849 3451
rect 7432 3420 7849 3448
rect 7432 3408 7438 3420
rect 7837 3417 7849 3420
rect 7883 3417 7895 3451
rect 7837 3411 7895 3417
rect 9600 3392 9628 3488
rect 9861 3485 9873 3488
rect 9907 3485 9919 3519
rect 9861 3479 9919 3485
rect 10597 3519 10655 3525
rect 10597 3485 10609 3519
rect 10643 3516 10655 3519
rect 10686 3516 10692 3528
rect 10643 3488 10692 3516
rect 10643 3485 10655 3488
rect 10597 3479 10655 3485
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3485 11391 3519
rect 11333 3479 11391 3485
rect 12437 3519 12495 3525
rect 12437 3485 12449 3519
rect 12483 3516 12495 3519
rect 13648 3516 13676 3624
rect 14366 3612 14372 3624
rect 14424 3612 14430 3664
rect 17402 3612 17408 3664
rect 17460 3652 17466 3664
rect 18322 3652 18328 3664
rect 17460 3624 18328 3652
rect 17460 3612 17466 3624
rect 18322 3612 18328 3624
rect 18380 3612 18386 3664
rect 18782 3612 18788 3664
rect 18840 3652 18846 3664
rect 18840 3624 21772 3652
rect 18840 3612 18846 3624
rect 13998 3544 14004 3596
rect 14056 3584 14062 3596
rect 14737 3587 14795 3593
rect 14737 3584 14749 3587
rect 14056 3556 14749 3584
rect 14056 3544 14062 3556
rect 14737 3553 14749 3556
rect 14783 3553 14795 3587
rect 14737 3547 14795 3553
rect 15470 3544 15476 3596
rect 15528 3584 15534 3596
rect 16577 3587 16635 3593
rect 16577 3584 16589 3587
rect 15528 3556 16589 3584
rect 15528 3544 15534 3556
rect 16577 3553 16589 3556
rect 16623 3553 16635 3587
rect 16577 3547 16635 3553
rect 17678 3544 17684 3596
rect 17736 3544 17742 3596
rect 18049 3587 18107 3593
rect 18049 3553 18061 3587
rect 18095 3584 18107 3587
rect 18690 3584 18696 3596
rect 18095 3556 18696 3584
rect 18095 3553 18107 3556
rect 18049 3547 18107 3553
rect 18690 3544 18696 3556
rect 18748 3544 18754 3596
rect 19518 3584 19524 3596
rect 19168 3556 19524 3584
rect 12483 3488 13676 3516
rect 14461 3519 14519 3525
rect 12483 3485 12495 3488
rect 12437 3479 12495 3485
rect 14461 3485 14473 3519
rect 14507 3516 14519 3519
rect 16022 3516 16028 3528
rect 14507 3488 16028 3516
rect 14507 3485 14519 3488
rect 14461 3479 14519 3485
rect 11348 3448 11376 3479
rect 16022 3476 16028 3488
rect 16080 3476 16086 3528
rect 16301 3519 16359 3525
rect 16301 3485 16313 3519
rect 16347 3516 16359 3519
rect 17696 3516 17724 3544
rect 16347 3488 17724 3516
rect 18325 3519 18383 3525
rect 16347 3485 16359 3488
rect 16301 3479 16359 3485
rect 18325 3485 18337 3519
rect 18371 3516 18383 3519
rect 19168 3516 19196 3556
rect 19518 3544 19524 3556
rect 19576 3544 19582 3596
rect 19889 3587 19947 3593
rect 19889 3553 19901 3587
rect 19935 3553 19947 3587
rect 19889 3547 19947 3553
rect 18371 3488 19196 3516
rect 18371 3485 18383 3488
rect 18325 3479 18383 3485
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 19392 3488 19441 3516
rect 19392 3476 19398 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 19429 3479 19487 3485
rect 15010 3448 15016 3460
rect 11348 3420 15016 3448
rect 15010 3408 15016 3420
rect 15068 3408 15074 3460
rect 17126 3448 17132 3460
rect 16316 3420 17132 3448
rect 3326 3340 3332 3392
rect 3384 3340 3390 3392
rect 3786 3340 3792 3392
rect 3844 3340 3850 3392
rect 6089 3383 6147 3389
rect 6089 3349 6101 3383
rect 6135 3380 6147 3383
rect 6270 3380 6276 3392
rect 6135 3352 6276 3380
rect 6135 3349 6147 3352
rect 6089 3343 6147 3349
rect 6270 3340 6276 3352
rect 6328 3340 6334 3392
rect 7742 3340 7748 3392
rect 7800 3340 7806 3392
rect 9217 3383 9275 3389
rect 9217 3349 9229 3383
rect 9263 3380 9275 3383
rect 9306 3380 9312 3392
rect 9263 3352 9312 3380
rect 9263 3349 9275 3352
rect 9217 3343 9275 3349
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 9401 3383 9459 3389
rect 9401 3349 9413 3383
rect 9447 3380 9459 3383
rect 9582 3380 9588 3392
rect 9447 3352 9588 3380
rect 9447 3349 9459 3352
rect 9401 3343 9459 3349
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 10318 3340 10324 3392
rect 10376 3380 10382 3392
rect 16316 3380 16344 3420
rect 17126 3408 17132 3420
rect 17184 3408 17190 3460
rect 17678 3408 17684 3460
rect 17736 3448 17742 3460
rect 19904 3448 19932 3547
rect 20070 3544 20076 3596
rect 20128 3584 20134 3596
rect 21744 3593 21772 3624
rect 21729 3587 21787 3593
rect 20128 3556 21496 3584
rect 20128 3544 20134 3556
rect 21358 3476 21364 3528
rect 21416 3476 21422 3528
rect 21468 3516 21496 3556
rect 21729 3553 21741 3587
rect 21775 3553 21787 3587
rect 21729 3547 21787 3553
rect 22738 3544 22744 3596
rect 22796 3584 22802 3596
rect 23201 3587 23259 3593
rect 23201 3584 23213 3587
rect 22796 3556 23213 3584
rect 22796 3544 22802 3556
rect 23201 3553 23213 3556
rect 23247 3553 23259 3587
rect 23201 3547 23259 3553
rect 21468 3488 23060 3516
rect 23032 3460 23060 3488
rect 24026 3476 24032 3528
rect 24084 3476 24090 3528
rect 24302 3476 24308 3528
rect 24360 3516 24366 3528
rect 24578 3516 24584 3528
rect 24360 3488 24584 3516
rect 24360 3476 24366 3488
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 17736 3420 19932 3448
rect 17736 3408 17742 3420
rect 21634 3408 21640 3460
rect 21692 3448 21698 3460
rect 22830 3448 22836 3460
rect 21692 3420 22836 3448
rect 21692 3408 21698 3420
rect 22830 3408 22836 3420
rect 22888 3408 22894 3460
rect 23014 3408 23020 3460
rect 23072 3448 23078 3460
rect 23750 3448 23756 3460
rect 23072 3420 23756 3448
rect 23072 3408 23078 3420
rect 23750 3408 23756 3420
rect 23808 3408 23814 3460
rect 10376 3352 16344 3380
rect 10376 3340 10382 3352
rect 16390 3340 16396 3392
rect 16448 3380 16454 3392
rect 20438 3380 20444 3392
rect 16448 3352 20444 3380
rect 16448 3340 16454 3352
rect 20438 3340 20444 3352
rect 20496 3340 20502 3392
rect 20530 3340 20536 3392
rect 20588 3380 20594 3392
rect 23106 3380 23112 3392
rect 20588 3352 23112 3380
rect 20588 3340 20594 3352
rect 23106 3340 23112 3352
rect 23164 3340 23170 3392
rect 24578 3340 24584 3392
rect 24636 3380 24642 3392
rect 25225 3383 25283 3389
rect 25225 3380 25237 3383
rect 24636 3352 25237 3380
rect 24636 3340 24642 3352
rect 25225 3349 25237 3352
rect 25271 3349 25283 3383
rect 25225 3343 25283 3349
rect 1104 3290 25852 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 25852 3290
rect 1104 3216 25852 3238
rect 7193 3179 7251 3185
rect 7193 3145 7205 3179
rect 7239 3176 7251 3179
rect 9122 3176 9128 3188
rect 7239 3148 9128 3176
rect 7239 3145 7251 3148
rect 7193 3139 7251 3145
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 9674 3136 9680 3188
rect 9732 3136 9738 3188
rect 10318 3136 10324 3188
rect 10376 3136 10382 3188
rect 10965 3179 11023 3185
rect 10965 3145 10977 3179
rect 11011 3176 11023 3179
rect 11330 3176 11336 3188
rect 11011 3148 11336 3176
rect 11011 3145 11023 3148
rect 10965 3139 11023 3145
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 13906 3176 13912 3188
rect 12406 3148 13912 3176
rect 9401 3111 9459 3117
rect 9401 3077 9413 3111
rect 9447 3108 9459 3111
rect 12406 3108 12434 3148
rect 13906 3136 13912 3148
rect 13964 3136 13970 3188
rect 14182 3136 14188 3188
rect 14240 3176 14246 3188
rect 16482 3176 16488 3188
rect 14240 3148 16488 3176
rect 14240 3136 14246 3148
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 17862 3136 17868 3188
rect 17920 3176 17926 3188
rect 17920 3148 20760 3176
rect 17920 3136 17926 3148
rect 14200 3108 14228 3136
rect 9447 3080 11192 3108
rect 9447 3077 9459 3080
rect 9401 3071 9459 3077
rect 2406 3000 2412 3052
rect 2464 3000 2470 3052
rect 3694 3000 3700 3052
rect 3752 3000 3758 3052
rect 5442 3000 5448 3052
rect 5500 3000 5506 3052
rect 6638 3000 6644 3052
rect 6696 3040 6702 3052
rect 6733 3043 6791 3049
rect 6733 3040 6745 3043
rect 6696 3012 6745 3040
rect 6696 3000 6702 3012
rect 6733 3009 6745 3012
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 7374 3000 7380 3052
rect 7432 3000 7438 3052
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3040 9091 3043
rect 9861 3043 9919 3049
rect 9861 3040 9873 3043
rect 9079 3012 9873 3040
rect 9079 3009 9091 3012
rect 9033 3003 9091 3009
rect 9861 3009 9873 3012
rect 9907 3040 9919 3043
rect 10318 3040 10324 3052
rect 9907 3012 10324 3040
rect 9907 3009 9919 3012
rect 9861 3003 9919 3009
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 10505 3043 10563 3049
rect 10505 3009 10517 3043
rect 10551 3040 10563 3043
rect 11054 3040 11060 3052
rect 10551 3012 11060 3040
rect 10551 3009 10563 3012
rect 10505 3003 10563 3009
rect 2133 2975 2191 2981
rect 2133 2941 2145 2975
rect 2179 2972 2191 2975
rect 2590 2972 2596 2984
rect 2179 2944 2596 2972
rect 2179 2941 2191 2944
rect 2133 2935 2191 2941
rect 2590 2932 2596 2944
rect 2648 2932 2654 2984
rect 3326 2932 3332 2984
rect 3384 2972 3390 2984
rect 3421 2975 3479 2981
rect 3421 2972 3433 2975
rect 3384 2944 3433 2972
rect 3384 2932 3390 2944
rect 3421 2941 3433 2944
rect 3467 2941 3479 2975
rect 3421 2935 3479 2941
rect 5166 2932 5172 2984
rect 5224 2932 5230 2984
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 7837 2975 7895 2981
rect 7837 2972 7849 2975
rect 7800 2944 7849 2972
rect 7800 2932 7806 2944
rect 7837 2941 7849 2944
rect 7883 2941 7895 2975
rect 7837 2935 7895 2941
rect 9217 2975 9275 2981
rect 9217 2941 9229 2975
rect 9263 2972 9275 2975
rect 10520 2972 10548 3003
rect 11054 3000 11060 3012
rect 11112 3000 11118 3052
rect 11164 3049 11192 3080
rect 11992 3080 12434 3108
rect 13188 3080 14228 3108
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3040 11207 3043
rect 11790 3040 11796 3052
rect 11195 3012 11796 3040
rect 11195 3009 11207 3012
rect 11149 3003 11207 3009
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 11992 3049 12020 3080
rect 13188 3049 13216 3080
rect 16574 3068 16580 3120
rect 16632 3108 16638 3120
rect 16632 3080 19196 3108
rect 16632 3068 16638 3080
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3009 13231 3043
rect 13173 3003 13231 3009
rect 14090 3000 14096 3052
rect 14148 3040 14154 3052
rect 14829 3043 14887 3049
rect 14829 3040 14841 3043
rect 14148 3012 14841 3040
rect 14148 3000 14154 3012
rect 14829 3009 14841 3012
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3040 17095 3043
rect 18598 3040 18604 3052
rect 17083 3012 18604 3040
rect 17083 3009 17095 3012
rect 17037 3003 17095 3009
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 18877 3043 18935 3049
rect 18877 3009 18889 3043
rect 18923 3040 18935 3043
rect 18966 3040 18972 3052
rect 18923 3012 18972 3040
rect 18923 3009 18935 3012
rect 18877 3003 18935 3009
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 9263 2944 10548 2972
rect 9263 2941 9275 2944
rect 9217 2935 9275 2941
rect 11422 2932 11428 2984
rect 11480 2972 11486 2984
rect 11698 2972 11704 2984
rect 11480 2944 11704 2972
rect 11480 2932 11486 2944
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 13630 2932 13636 2984
rect 13688 2932 13694 2984
rect 14734 2932 14740 2984
rect 14792 2972 14798 2984
rect 15289 2975 15347 2981
rect 15289 2972 15301 2975
rect 14792 2944 15301 2972
rect 14792 2932 14798 2944
rect 15289 2941 15301 2944
rect 15335 2941 15347 2975
rect 15289 2935 15347 2941
rect 15838 2932 15844 2984
rect 15896 2972 15902 2984
rect 19168 2981 19196 3080
rect 20530 3068 20536 3120
rect 20588 3108 20594 3120
rect 20625 3111 20683 3117
rect 20625 3108 20637 3111
rect 20588 3080 20637 3108
rect 20588 3068 20594 3080
rect 20625 3077 20637 3080
rect 20671 3077 20683 3111
rect 20625 3071 20683 3077
rect 20732 3040 20760 3148
rect 20898 3136 20904 3188
rect 20956 3176 20962 3188
rect 21269 3179 21327 3185
rect 21269 3176 21281 3179
rect 20956 3148 21281 3176
rect 20956 3136 20962 3148
rect 21269 3145 21281 3148
rect 21315 3145 21327 3179
rect 21269 3139 21327 3145
rect 22186 3136 22192 3188
rect 22244 3136 22250 3188
rect 22554 3136 22560 3188
rect 22612 3176 22618 3188
rect 22925 3179 22983 3185
rect 22925 3176 22937 3179
rect 22612 3148 22937 3176
rect 22612 3136 22618 3148
rect 22925 3145 22937 3148
rect 22971 3145 22983 3179
rect 22925 3139 22983 3145
rect 23658 3136 23664 3188
rect 23716 3136 23722 3188
rect 24210 3136 24216 3188
rect 24268 3136 24274 3188
rect 20809 3111 20867 3117
rect 20809 3077 20821 3111
rect 20855 3108 20867 3111
rect 21910 3108 21916 3120
rect 20855 3080 21916 3108
rect 20855 3077 20867 3080
rect 20809 3071 20867 3077
rect 21910 3068 21916 3080
rect 21968 3068 21974 3120
rect 22094 3068 22100 3120
rect 22152 3068 22158 3120
rect 22833 3111 22891 3117
rect 22833 3077 22845 3111
rect 22879 3108 22891 3111
rect 23014 3108 23020 3120
rect 22879 3080 23020 3108
rect 22879 3077 22891 3080
rect 22833 3071 22891 3077
rect 23014 3068 23020 3080
rect 23072 3068 23078 3120
rect 23566 3068 23572 3120
rect 23624 3068 23630 3120
rect 23750 3068 23756 3120
rect 23808 3108 23814 3120
rect 25409 3111 25467 3117
rect 25409 3108 25421 3111
rect 23808 3080 25421 3108
rect 23808 3068 23814 3080
rect 25409 3077 25421 3080
rect 25455 3077 25467 3111
rect 25409 3071 25467 3077
rect 21818 3040 21824 3052
rect 20732 3012 21824 3040
rect 21818 3000 21824 3012
rect 21876 3000 21882 3052
rect 22922 3000 22928 3052
rect 22980 3040 22986 3052
rect 24397 3043 24455 3049
rect 24397 3040 24409 3043
rect 22980 3012 24409 3040
rect 22980 3000 22986 3012
rect 24397 3009 24409 3012
rect 24443 3009 24455 3043
rect 24397 3003 24455 3009
rect 25130 3000 25136 3052
rect 25188 3000 25194 3052
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 15896 2944 17325 2972
rect 15896 2932 15902 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 19153 2975 19211 2981
rect 19153 2941 19165 2975
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 21358 2932 21364 2984
rect 21416 2972 21422 2984
rect 23474 2972 23480 2984
rect 21416 2944 23480 2972
rect 21416 2932 21422 2944
rect 23474 2932 23480 2944
rect 23532 2932 23538 2984
rect 6549 2907 6607 2913
rect 6549 2873 6561 2907
rect 6595 2904 6607 2907
rect 11146 2904 11152 2916
rect 6595 2876 11152 2904
rect 6595 2873 6607 2876
rect 6549 2867 6607 2873
rect 11146 2864 11152 2876
rect 11204 2864 11210 2916
rect 15102 2864 15108 2916
rect 15160 2904 15166 2916
rect 17218 2904 17224 2916
rect 15160 2876 17224 2904
rect 15160 2864 15166 2876
rect 17218 2864 17224 2876
rect 17276 2864 17282 2916
rect 19518 2864 19524 2916
rect 19576 2904 19582 2916
rect 22094 2904 22100 2916
rect 19576 2876 22100 2904
rect 19576 2864 19582 2876
rect 22094 2864 22100 2876
rect 22152 2864 22158 2916
rect 24946 2864 24952 2916
rect 25004 2864 25010 2916
rect 4430 2796 4436 2848
rect 4488 2836 4494 2848
rect 4525 2839 4583 2845
rect 4525 2836 4537 2839
rect 4488 2808 4537 2836
rect 4488 2796 4494 2808
rect 4525 2805 4537 2808
rect 4571 2805 4583 2839
rect 4525 2799 4583 2805
rect 4890 2796 4896 2848
rect 4948 2796 4954 2848
rect 8067 2839 8125 2845
rect 8067 2805 8079 2839
rect 8113 2836 8125 2839
rect 14826 2836 14832 2848
rect 8113 2808 14832 2836
rect 8113 2805 8125 2808
rect 8067 2799 8125 2805
rect 14826 2796 14832 2808
rect 14884 2796 14890 2848
rect 16942 2796 16948 2848
rect 17000 2836 17006 2848
rect 19886 2836 19892 2848
rect 17000 2808 19892 2836
rect 17000 2796 17006 2808
rect 19886 2796 19892 2808
rect 19944 2796 19950 2848
rect 1104 2746 25852 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 25852 2746
rect 1104 2672 25852 2694
rect 8389 2635 8447 2641
rect 8389 2601 8401 2635
rect 8435 2632 8447 2635
rect 8570 2632 8576 2644
rect 8435 2604 8576 2632
rect 8435 2601 8447 2604
rect 8389 2595 8447 2601
rect 8570 2592 8576 2604
rect 8628 2592 8634 2644
rect 15746 2632 15752 2644
rect 9876 2604 15752 2632
rect 9766 2564 9772 2576
rect 2884 2536 9772 2564
rect 2884 2505 2912 2536
rect 9766 2524 9772 2536
rect 9824 2524 9830 2576
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2465 2927 2499
rect 2869 2459 2927 2465
rect 5442 2456 5448 2508
rect 5500 2456 5506 2508
rect 6825 2499 6883 2505
rect 6825 2465 6837 2499
rect 6871 2496 6883 2499
rect 6871 2468 8340 2496
rect 6871 2465 6883 2468
rect 6825 2459 6883 2465
rect 8312 2440 8340 2468
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 2958 2428 2964 2440
rect 2639 2400 2964 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 2958 2388 2964 2400
rect 3016 2428 3022 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3016 2400 3985 2428
rect 3016 2388 3022 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 4249 2363 4307 2369
rect 4249 2329 4261 2363
rect 4295 2360 4307 2363
rect 4724 2360 4752 2391
rect 4890 2388 4896 2440
rect 4948 2428 4954 2440
rect 5169 2431 5227 2437
rect 5169 2428 5181 2431
rect 4948 2400 5181 2428
rect 4948 2388 4954 2400
rect 5169 2397 5181 2400
rect 5215 2428 5227 2431
rect 5534 2428 5540 2440
rect 5215 2400 5540 2428
rect 5215 2397 5227 2400
rect 5169 2391 5227 2397
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 6641 2431 6699 2437
rect 6641 2397 6653 2431
rect 6687 2428 6699 2431
rect 7285 2431 7343 2437
rect 7285 2428 7297 2431
rect 6687 2400 7297 2428
rect 6687 2397 6699 2400
rect 6641 2391 6699 2397
rect 7285 2397 7297 2400
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 5902 2360 5908 2372
rect 4295 2332 5908 2360
rect 4295 2329 4307 2332
rect 4249 2323 4307 2329
rect 5902 2320 5908 2332
rect 5960 2320 5966 2372
rect 7300 2360 7328 2391
rect 7834 2388 7840 2440
rect 7892 2428 7898 2440
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 7892 2400 7941 2428
rect 7892 2388 7898 2400
rect 7929 2397 7941 2400
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 8294 2388 8300 2440
rect 8352 2428 8358 2440
rect 8573 2431 8631 2437
rect 8573 2428 8585 2431
rect 8352 2400 8585 2428
rect 8352 2388 8358 2400
rect 8573 2397 8585 2400
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 9306 2388 9312 2440
rect 9364 2388 9370 2440
rect 9876 2437 9904 2604
rect 15746 2592 15752 2604
rect 15804 2592 15810 2644
rect 16022 2592 16028 2644
rect 16080 2632 16086 2644
rect 16117 2635 16175 2641
rect 16117 2632 16129 2635
rect 16080 2604 16129 2632
rect 16080 2592 16086 2604
rect 16117 2601 16129 2604
rect 16163 2601 16175 2635
rect 16117 2595 16175 2601
rect 16408 2604 18644 2632
rect 13446 2524 13452 2576
rect 13504 2564 13510 2576
rect 16408 2564 16436 2604
rect 18616 2564 18644 2604
rect 18690 2592 18696 2644
rect 18748 2592 18754 2644
rect 22278 2592 22284 2644
rect 22336 2632 22342 2644
rect 23198 2632 23204 2644
rect 22336 2604 23204 2632
rect 22336 2592 22342 2604
rect 23198 2592 23204 2604
rect 23256 2592 23262 2644
rect 21269 2567 21327 2573
rect 21269 2564 21281 2567
rect 13504 2536 16436 2564
rect 16546 2536 18552 2564
rect 18616 2536 21281 2564
rect 13504 2524 13510 2536
rect 10965 2499 11023 2505
rect 10965 2465 10977 2499
rect 11011 2496 11023 2499
rect 11011 2468 14228 2496
rect 11011 2465 11023 2468
rect 10965 2459 11023 2465
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2397 9919 2431
rect 9861 2391 9919 2397
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2428 11943 2431
rect 12158 2428 12164 2440
rect 11931 2400 12164 2428
rect 11931 2397 11943 2400
rect 11885 2391 11943 2397
rect 12158 2388 12164 2400
rect 12216 2388 12222 2440
rect 12434 2388 12440 2440
rect 12492 2388 12498 2440
rect 14090 2388 14096 2440
rect 14148 2388 14154 2440
rect 8846 2360 8852 2372
rect 7300 2332 8852 2360
rect 8846 2320 8852 2332
rect 8904 2320 8910 2372
rect 9324 2360 9352 2388
rect 9950 2360 9956 2372
rect 9324 2332 9956 2360
rect 9950 2320 9956 2332
rect 10008 2320 10014 2372
rect 11974 2360 11980 2372
rect 10520 2332 11980 2360
rect 2590 2252 2596 2304
rect 2648 2292 2654 2304
rect 3789 2295 3847 2301
rect 3789 2292 3801 2295
rect 2648 2264 3801 2292
rect 2648 2252 2654 2264
rect 3789 2261 3801 2264
rect 3835 2261 3847 2295
rect 3789 2255 3847 2261
rect 4522 2252 4528 2304
rect 4580 2252 4586 2304
rect 6457 2295 6515 2301
rect 6457 2261 6469 2295
rect 6503 2292 6515 2295
rect 6638 2292 6644 2304
rect 6503 2264 6644 2292
rect 6503 2261 6515 2264
rect 6457 2255 6515 2261
rect 6638 2252 6644 2264
rect 6696 2252 6702 2304
rect 7098 2252 7104 2304
rect 7156 2252 7162 2304
rect 7745 2295 7803 2301
rect 7745 2261 7757 2295
rect 7791 2292 7803 2295
rect 8386 2292 8392 2304
rect 7791 2264 8392 2292
rect 7791 2261 7803 2264
rect 7745 2255 7803 2261
rect 8386 2252 8392 2264
rect 8444 2252 8450 2304
rect 9125 2295 9183 2301
rect 9125 2261 9137 2295
rect 9171 2292 9183 2295
rect 10520 2292 10548 2332
rect 11974 2320 11980 2332
rect 12032 2320 12038 2372
rect 13262 2320 13268 2372
rect 13320 2320 13326 2372
rect 14200 2360 14228 2468
rect 14366 2456 14372 2508
rect 14424 2496 14430 2508
rect 14921 2499 14979 2505
rect 14921 2496 14933 2499
rect 14424 2468 14933 2496
rect 14424 2456 14430 2468
rect 14921 2465 14933 2468
rect 14967 2465 14979 2499
rect 14921 2459 14979 2465
rect 16022 2456 16028 2508
rect 16080 2496 16086 2508
rect 16393 2499 16451 2505
rect 16393 2496 16405 2499
rect 16080 2468 16405 2496
rect 16080 2456 16086 2468
rect 16393 2465 16405 2468
rect 16439 2465 16451 2499
rect 16393 2459 16451 2465
rect 14458 2388 14464 2440
rect 14516 2388 14522 2440
rect 16114 2388 16120 2440
rect 16172 2428 16178 2440
rect 16546 2428 16574 2536
rect 17310 2456 17316 2508
rect 17368 2456 17374 2508
rect 18524 2496 18552 2536
rect 21269 2533 21281 2536
rect 21315 2533 21327 2567
rect 22186 2564 22192 2576
rect 21269 2527 21327 2533
rect 21376 2536 22192 2564
rect 18524 2468 19564 2496
rect 16172 2400 16574 2428
rect 16172 2388 16178 2400
rect 16758 2388 16764 2440
rect 16816 2428 16822 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16816 2400 16865 2428
rect 16816 2388 16822 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 18877 2431 18935 2437
rect 18877 2397 18889 2431
rect 18923 2397 18935 2431
rect 18877 2391 18935 2397
rect 18892 2360 18920 2391
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 19536 2428 19564 2468
rect 19886 2456 19892 2508
rect 19944 2456 19950 2508
rect 21376 2428 21404 2536
rect 22186 2524 22192 2536
rect 22244 2524 22250 2576
rect 22094 2456 22100 2508
rect 22152 2496 22158 2508
rect 22465 2499 22523 2505
rect 22465 2496 22477 2499
rect 22152 2468 22477 2496
rect 22152 2456 22158 2468
rect 22465 2465 22477 2468
rect 22511 2465 22523 2499
rect 22465 2459 22523 2465
rect 23845 2499 23903 2505
rect 23845 2465 23857 2499
rect 23891 2496 23903 2499
rect 24854 2496 24860 2508
rect 23891 2468 24860 2496
rect 23891 2465 23903 2468
rect 23845 2459 23903 2465
rect 24854 2456 24860 2468
rect 24912 2456 24918 2508
rect 19536 2400 21404 2428
rect 21450 2388 21456 2440
rect 21508 2388 21514 2440
rect 22189 2431 22247 2437
rect 22189 2397 22201 2431
rect 22235 2397 22247 2431
rect 22189 2391 22247 2397
rect 22204 2360 22232 2391
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 25130 2360 25136 2372
rect 14200 2332 16574 2360
rect 18892 2332 22140 2360
rect 22204 2332 25136 2360
rect 9171 2264 10548 2292
rect 11701 2295 11759 2301
rect 9171 2261 9183 2264
rect 9125 2255 9183 2261
rect 11701 2261 11713 2295
rect 11747 2292 11759 2295
rect 15654 2292 15660 2304
rect 11747 2264 15660 2292
rect 11747 2261 11759 2264
rect 11701 2255 11759 2261
rect 15654 2252 15660 2264
rect 15712 2252 15718 2304
rect 16546 2292 16574 2332
rect 21174 2292 21180 2304
rect 16546 2264 21180 2292
rect 21174 2252 21180 2264
rect 21232 2252 21238 2304
rect 22112 2292 22140 2332
rect 25130 2320 25136 2332
rect 25188 2320 25194 2372
rect 23290 2292 23296 2304
rect 22112 2264 23296 2292
rect 23290 2252 23296 2264
rect 23348 2252 23354 2304
rect 25222 2252 25228 2304
rect 25280 2252 25286 2304
rect 1104 2202 25852 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 25852 2202
rect 1104 2128 25852 2150
rect 4522 2048 4528 2100
rect 4580 2088 4586 2100
rect 4580 2060 6914 2088
rect 4580 2048 4586 2060
rect 6886 2020 6914 2060
rect 8386 2048 8392 2100
rect 8444 2088 8450 2100
rect 15194 2088 15200 2100
rect 8444 2060 15200 2088
rect 8444 2048 8450 2060
rect 15194 2048 15200 2060
rect 15252 2048 15258 2100
rect 11330 2020 11336 2032
rect 6886 1992 11336 2020
rect 11330 1980 11336 1992
rect 11388 1980 11394 2032
rect 7834 1912 7840 1964
rect 7892 1952 7898 1964
rect 17034 1952 17040 1964
rect 7892 1924 17040 1952
rect 7892 1912 7898 1924
rect 17034 1912 17040 1924
rect 17092 1912 17098 1964
rect 7098 1844 7104 1896
rect 7156 1884 7162 1896
rect 12710 1884 12716 1896
rect 7156 1856 12716 1884
rect 7156 1844 7162 1856
rect 12710 1844 12716 1856
rect 12768 1844 12774 1896
rect 11238 1776 11244 1828
rect 11296 1816 11302 1828
rect 25222 1816 25228 1828
rect 11296 1788 25228 1816
rect 11296 1776 11302 1788
rect 25222 1776 25228 1788
rect 25280 1776 25286 1828
<< via1 >>
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 13820 54315 13872 54324
rect 13820 54281 13829 54315
rect 13829 54281 13863 54315
rect 13863 54281 13872 54315
rect 13820 54272 13872 54281
rect 4068 54136 4120 54188
rect 4804 54179 4856 54188
rect 4804 54145 4813 54179
rect 4813 54145 4847 54179
rect 4847 54145 4856 54179
rect 4804 54136 4856 54145
rect 7380 54179 7432 54188
rect 7380 54145 7389 54179
rect 7389 54145 7423 54179
rect 7423 54145 7432 54179
rect 7380 54136 7432 54145
rect 9588 54179 9640 54188
rect 9588 54145 9597 54179
rect 9597 54145 9631 54179
rect 9631 54145 9640 54179
rect 9588 54136 9640 54145
rect 11704 54136 11756 54188
rect 2412 54068 2464 54120
rect 5172 54111 5224 54120
rect 5172 54077 5181 54111
rect 5181 54077 5215 54111
rect 5215 54077 5224 54111
rect 5172 54068 5224 54077
rect 7840 54111 7892 54120
rect 7840 54077 7849 54111
rect 7849 54077 7883 54111
rect 7883 54077 7892 54111
rect 7840 54068 7892 54077
rect 9312 54068 9364 54120
rect 12348 54068 12400 54120
rect 14832 54136 14884 54188
rect 16580 54136 16632 54188
rect 17592 54136 17644 54188
rect 18972 54315 19024 54324
rect 18972 54281 18981 54315
rect 18981 54281 19015 54315
rect 19015 54281 19024 54315
rect 18972 54272 19024 54281
rect 20720 54179 20772 54188
rect 20720 54145 20729 54179
rect 20729 54145 20763 54179
rect 20763 54145 20772 54179
rect 20720 54136 20772 54145
rect 21732 54136 21784 54188
rect 23112 54136 23164 54188
rect 25872 54136 25924 54188
rect 8576 54000 8628 54052
rect 13912 54000 13964 54052
rect 15660 54000 15712 54052
rect 20168 54000 20220 54052
rect 12716 53932 12768 53984
rect 15568 53932 15620 53984
rect 16948 53932 17000 53984
rect 22100 53932 22152 53984
rect 25044 53932 25096 53984
rect 25320 53975 25372 53984
rect 25320 53941 25329 53975
rect 25329 53941 25363 53975
rect 25363 53941 25372 53975
rect 25320 53932 25372 53941
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 24492 53771 24544 53780
rect 24492 53737 24501 53771
rect 24501 53737 24535 53771
rect 24535 53737 24544 53771
rect 24492 53728 24544 53737
rect 24768 53771 24820 53780
rect 24768 53737 24777 53771
rect 24777 53737 24811 53771
rect 24811 53737 24820 53771
rect 24768 53728 24820 53737
rect 10692 53660 10744 53712
rect 1032 53592 1084 53644
rect 3792 53592 3844 53644
rect 6552 53592 6604 53644
rect 4160 53567 4212 53576
rect 4160 53533 4169 53567
rect 4169 53533 4203 53567
rect 4203 53533 4212 53567
rect 4160 53524 4212 53533
rect 7840 53524 7892 53576
rect 10692 53524 10744 53576
rect 23388 53524 23440 53576
rect 24492 53524 24544 53576
rect 25044 53567 25096 53576
rect 25044 53533 25053 53567
rect 25053 53533 25087 53567
rect 25087 53533 25096 53567
rect 25044 53524 25096 53533
rect 5540 53456 5592 53508
rect 22836 53388 22888 53440
rect 23940 53431 23992 53440
rect 23940 53397 23949 53431
rect 23949 53397 23983 53431
rect 23983 53397 23992 53431
rect 23940 53388 23992 53397
rect 25872 53388 25924 53440
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 4068 53184 4120 53236
rect 7748 53048 7800 53100
rect 24768 53048 24820 53100
rect 25044 53091 25096 53100
rect 25044 53057 25053 53091
rect 25053 53057 25087 53091
rect 25087 53057 25096 53091
rect 25044 53048 25096 53057
rect 24400 52980 24452 53032
rect 18696 52912 18748 52964
rect 23756 52887 23808 52896
rect 23756 52853 23765 52887
rect 23765 52853 23799 52887
rect 23799 52853 23808 52887
rect 23756 52844 23808 52853
rect 24492 52887 24544 52896
rect 24492 52853 24501 52887
rect 24501 52853 24535 52887
rect 24535 52853 24544 52887
rect 24492 52844 24544 52853
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 4160 52640 4212 52692
rect 24400 52640 24452 52692
rect 9496 52436 9548 52488
rect 26516 52436 26568 52488
rect 24952 52411 25004 52420
rect 24952 52377 24961 52411
rect 24961 52377 24995 52411
rect 24995 52377 25004 52411
rect 24952 52368 25004 52377
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 25044 52096 25096 52148
rect 25320 52003 25372 52012
rect 25320 51969 25329 52003
rect 25329 51969 25363 52003
rect 25363 51969 25372 52003
rect 25320 51960 25372 51969
rect 23388 51756 23440 51808
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 7380 51552 7432 51604
rect 7840 51484 7892 51536
rect 4804 51348 4856 51400
rect 8484 51391 8536 51400
rect 8484 51357 8493 51391
rect 8493 51357 8527 51391
rect 8527 51357 8536 51391
rect 8484 51348 8536 51357
rect 10508 51348 10560 51400
rect 10784 51280 10836 51332
rect 24952 51323 25004 51332
rect 24952 51289 24961 51323
rect 24961 51289 24995 51323
rect 24995 51289 25004 51323
rect 24952 51280 25004 51289
rect 26608 51280 26660 51332
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 24952 50915 25004 50924
rect 24952 50881 24961 50915
rect 24961 50881 24995 50915
rect 24995 50881 25004 50915
rect 24952 50872 25004 50881
rect 18604 50668 18656 50720
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 5540 50464 5592 50516
rect 8392 50464 8444 50516
rect 9588 50507 9640 50516
rect 9588 50473 9597 50507
rect 9597 50473 9631 50507
rect 9631 50473 9640 50507
rect 9588 50464 9640 50473
rect 7748 50396 7800 50448
rect 8576 50328 8628 50380
rect 9588 50192 9640 50244
rect 25504 50167 25556 50176
rect 25504 50133 25513 50167
rect 25513 50133 25547 50167
rect 25547 50133 25556 50167
rect 25504 50124 25556 50133
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 25504 49784 25556 49836
rect 24676 49716 24728 49768
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 10692 49351 10744 49360
rect 10692 49317 10701 49351
rect 10701 49317 10735 49351
rect 10735 49317 10744 49351
rect 10692 49308 10744 49317
rect 11704 49351 11756 49360
rect 11704 49317 11713 49351
rect 11713 49317 11747 49351
rect 11747 49317 11756 49351
rect 11704 49308 11756 49317
rect 10232 49104 10284 49156
rect 10876 49104 10928 49156
rect 25136 49147 25188 49156
rect 25136 49113 25145 49147
rect 25145 49113 25179 49147
rect 25179 49113 25188 49147
rect 25136 49104 25188 49113
rect 20076 49036 20128 49088
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 9128 48832 9180 48884
rect 8300 48628 8352 48680
rect 8392 48671 8444 48680
rect 8392 48637 8401 48671
rect 8401 48637 8435 48671
rect 8435 48637 8444 48671
rect 8392 48628 8444 48637
rect 9956 48560 10008 48612
rect 9128 48492 9180 48544
rect 25136 48492 25188 48544
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 7748 48084 7800 48136
rect 23388 48127 23440 48136
rect 23388 48093 23397 48127
rect 23397 48093 23431 48127
rect 23431 48093 23440 48127
rect 23388 48084 23440 48093
rect 25136 48127 25188 48136
rect 25136 48093 25145 48127
rect 25145 48093 25179 48127
rect 25179 48093 25188 48127
rect 25136 48084 25188 48093
rect 17592 48016 17644 48068
rect 12624 47948 12676 48000
rect 24032 47991 24084 48000
rect 24032 47957 24041 47991
rect 24041 47957 24075 47991
rect 24075 47957 24084 47991
rect 24032 47948 24084 47957
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 9220 47744 9272 47796
rect 9496 47744 9548 47796
rect 8576 47676 8628 47728
rect 10968 47676 11020 47728
rect 25320 47651 25372 47660
rect 25320 47617 25329 47651
rect 25329 47617 25363 47651
rect 25363 47617 25372 47651
rect 25320 47608 25372 47617
rect 8300 47404 8352 47456
rect 9496 47447 9548 47456
rect 9496 47413 9505 47447
rect 9505 47413 9539 47447
rect 9539 47413 9548 47447
rect 9496 47404 9548 47413
rect 24952 47404 25004 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 9220 46996 9272 47048
rect 13728 46928 13780 46980
rect 25320 46860 25372 46912
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 10784 46699 10836 46708
rect 10784 46665 10793 46699
rect 10793 46665 10827 46699
rect 10827 46665 10836 46699
rect 10784 46656 10836 46665
rect 10968 46656 11020 46708
rect 13728 46588 13780 46640
rect 10784 46520 10836 46572
rect 13912 46563 13964 46572
rect 13912 46529 13921 46563
rect 13921 46529 13955 46563
rect 13955 46529 13964 46563
rect 13912 46520 13964 46529
rect 25320 46563 25372 46572
rect 25320 46529 25329 46563
rect 25329 46529 25363 46563
rect 25363 46529 25372 46563
rect 25320 46520 25372 46529
rect 15752 46495 15804 46504
rect 15752 46461 15761 46495
rect 15761 46461 15795 46495
rect 15795 46461 15804 46495
rect 15752 46452 15804 46461
rect 10784 46384 10836 46436
rect 10416 46359 10468 46368
rect 10416 46325 10425 46359
rect 10425 46325 10459 46359
rect 10459 46325 10468 46359
rect 10416 46316 10468 46325
rect 15016 46316 15068 46368
rect 25688 46316 25740 46368
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 8484 46155 8536 46164
rect 8484 46121 8493 46155
rect 8493 46121 8527 46155
rect 8527 46121 8536 46155
rect 8484 46112 8536 46121
rect 7748 45976 7800 46028
rect 15568 46044 15620 46096
rect 15016 46019 15068 46028
rect 15016 45985 15025 46019
rect 15025 45985 15059 46019
rect 15059 45985 15068 46019
rect 15016 45976 15068 45985
rect 16488 46019 16540 46028
rect 16488 45985 16497 46019
rect 16497 45985 16531 46019
rect 16531 45985 16540 46019
rect 16488 45976 16540 45985
rect 7840 45908 7892 45960
rect 12532 45908 12584 45960
rect 25320 45951 25372 45960
rect 25320 45917 25329 45951
rect 25329 45917 25363 45951
rect 25363 45917 25372 45951
rect 25320 45908 25372 45917
rect 15108 45772 15160 45824
rect 26056 45772 26108 45824
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 10508 45500 10560 45552
rect 12532 45500 12584 45552
rect 12624 45500 12676 45552
rect 12716 45475 12768 45484
rect 12716 45441 12725 45475
rect 12725 45441 12759 45475
rect 12759 45441 12768 45475
rect 12716 45432 12768 45441
rect 14556 45407 14608 45416
rect 14556 45373 14565 45407
rect 14565 45373 14599 45407
rect 14599 45373 14608 45407
rect 14556 45364 14608 45373
rect 25320 45228 25372 45280
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 9496 45024 9548 45076
rect 9956 44888 10008 44940
rect 9128 44863 9180 44872
rect 9128 44829 9137 44863
rect 9137 44829 9171 44863
rect 9171 44829 9180 44863
rect 9128 44820 9180 44829
rect 9680 44752 9732 44804
rect 15660 44931 15712 44940
rect 15660 44897 15669 44931
rect 15669 44897 15703 44931
rect 15703 44897 15712 44931
rect 15660 44888 15712 44897
rect 25320 44863 25372 44872
rect 25320 44829 25329 44863
rect 25329 44829 25363 44863
rect 25363 44829 25372 44863
rect 25320 44820 25372 44829
rect 11520 44752 11572 44804
rect 15108 44752 15160 44804
rect 19984 44752 20036 44804
rect 10416 44684 10468 44736
rect 11704 44684 11756 44736
rect 25228 44684 25280 44736
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 9588 44523 9640 44532
rect 9588 44489 9597 44523
rect 9597 44489 9631 44523
rect 9631 44489 9640 44523
rect 9588 44480 9640 44489
rect 9220 44344 9272 44396
rect 10784 44344 10836 44396
rect 24768 44387 24820 44396
rect 24768 44353 24777 44387
rect 24777 44353 24811 44387
rect 24811 44353 24820 44387
rect 24768 44344 24820 44353
rect 9036 44276 9088 44328
rect 10508 44208 10560 44260
rect 10692 44183 10744 44192
rect 10692 44149 10701 44183
rect 10701 44149 10735 44183
rect 10735 44149 10744 44183
rect 10692 44140 10744 44149
rect 10968 44140 11020 44192
rect 16856 44140 16908 44192
rect 22836 44140 22888 44192
rect 24860 44140 24912 44192
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 16580 43936 16632 43988
rect 24032 43800 24084 43852
rect 19524 43732 19576 43784
rect 21088 43664 21140 43716
rect 25504 43639 25556 43648
rect 25504 43605 25513 43639
rect 25513 43605 25547 43639
rect 25547 43605 25556 43639
rect 25504 43596 25556 43605
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 25504 43324 25556 43376
rect 24216 43052 24268 43104
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 10232 42755 10284 42764
rect 10232 42721 10241 42755
rect 10241 42721 10275 42755
rect 10275 42721 10284 42755
rect 10232 42712 10284 42721
rect 8944 42644 8996 42696
rect 10600 42644 10652 42696
rect 25136 42619 25188 42628
rect 25136 42585 25145 42619
rect 25145 42585 25179 42619
rect 25179 42585 25188 42619
rect 25136 42576 25188 42585
rect 24308 42508 24360 42560
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 9680 42304 9732 42356
rect 11520 42236 11572 42288
rect 9128 42100 9180 42152
rect 9772 42100 9824 42152
rect 10692 42100 10744 42152
rect 15568 42032 15620 42084
rect 24492 42032 24544 42084
rect 11520 42007 11572 42016
rect 11520 41973 11529 42007
rect 11529 41973 11563 42007
rect 11563 41973 11572 42007
rect 11520 41964 11572 41973
rect 11704 42007 11756 42016
rect 11704 41973 11713 42007
rect 11713 41973 11747 42007
rect 11747 41973 11756 42007
rect 11704 41964 11756 41973
rect 25136 41964 25188 42016
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 10876 41803 10928 41812
rect 10876 41769 10885 41803
rect 10885 41769 10919 41803
rect 10919 41769 10928 41803
rect 10876 41760 10928 41769
rect 16212 41692 16264 41744
rect 18696 41692 18748 41744
rect 10968 41624 11020 41676
rect 10232 41599 10284 41608
rect 10232 41565 10241 41599
rect 10241 41565 10275 41599
rect 10275 41565 10284 41599
rect 10232 41556 10284 41565
rect 25136 41599 25188 41608
rect 25136 41565 25145 41599
rect 25145 41565 25179 41599
rect 25179 41565 25188 41599
rect 25136 41556 25188 41565
rect 21364 41488 21416 41540
rect 20260 41420 20312 41472
rect 24676 41420 24728 41472
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 25320 41123 25372 41132
rect 25320 41089 25329 41123
rect 25329 41089 25363 41123
rect 25363 41089 25372 41123
rect 25320 41080 25372 41089
rect 25044 40876 25096 40928
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 25504 40375 25556 40384
rect 25504 40341 25513 40375
rect 25513 40341 25547 40375
rect 25547 40341 25556 40375
rect 25504 40332 25556 40341
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 23296 40128 23348 40180
rect 25504 40060 25556 40112
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 25320 39423 25372 39432
rect 25320 39389 25329 39423
rect 25329 39389 25363 39423
rect 25363 39389 25372 39423
rect 25320 39380 25372 39389
rect 21916 39244 21968 39296
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 25320 38700 25372 38752
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 25320 38335 25372 38344
rect 25320 38301 25329 38335
rect 25329 38301 25363 38335
rect 25363 38301 25372 38335
rect 25320 38292 25372 38301
rect 25412 38156 25464 38208
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 7840 37952 7892 38004
rect 8852 37859 8904 37868
rect 8852 37825 8861 37859
rect 8861 37825 8895 37859
rect 8895 37825 8904 37859
rect 8852 37816 8904 37825
rect 25136 37859 25188 37868
rect 25136 37825 25145 37859
rect 25145 37825 25179 37859
rect 25179 37825 25188 37859
rect 25136 37816 25188 37825
rect 25780 37680 25832 37732
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 16304 37272 16356 37324
rect 18604 37272 18656 37324
rect 25504 37111 25556 37120
rect 25504 37077 25513 37111
rect 25513 37077 25547 37111
rect 25547 37077 25556 37111
rect 25504 37068 25556 37077
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 25504 36796 25556 36848
rect 25596 36592 25648 36644
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 25320 36159 25372 36168
rect 25320 36125 25329 36159
rect 25329 36125 25363 36159
rect 25363 36125 25372 36159
rect 25320 36116 25372 36125
rect 25136 36023 25188 36032
rect 25136 35989 25145 36023
rect 25145 35989 25179 36023
rect 25179 35989 25188 36023
rect 25136 35980 25188 35989
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 11704 35776 11756 35828
rect 26056 35776 26108 35828
rect 11520 35751 11572 35760
rect 11520 35717 11529 35751
rect 11529 35717 11563 35751
rect 11563 35717 11572 35751
rect 11520 35708 11572 35717
rect 12164 35708 12216 35760
rect 25688 35708 25740 35760
rect 9680 35615 9732 35624
rect 9680 35581 9689 35615
rect 9689 35581 9723 35615
rect 9723 35581 9732 35615
rect 9680 35572 9732 35581
rect 9772 35572 9824 35624
rect 11796 35479 11848 35488
rect 11796 35445 11805 35479
rect 11805 35445 11839 35479
rect 11839 35445 11848 35479
rect 11796 35436 11848 35445
rect 15752 35436 15804 35488
rect 21824 35640 21876 35692
rect 22192 35572 22244 35624
rect 22560 35615 22612 35624
rect 22560 35581 22569 35615
rect 22569 35581 22603 35615
rect 22603 35581 22612 35615
rect 22560 35572 22612 35581
rect 20628 35436 20680 35488
rect 21180 35436 21232 35488
rect 22008 35479 22060 35488
rect 22008 35445 22017 35479
rect 22017 35445 22051 35479
rect 22051 35445 22060 35479
rect 22008 35436 22060 35445
rect 25320 35436 25372 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 22744 35096 22796 35148
rect 25228 35028 25280 35080
rect 25320 35071 25372 35080
rect 25320 35037 25329 35071
rect 25329 35037 25363 35071
rect 25363 35037 25372 35071
rect 25320 35028 25372 35037
rect 19984 34960 20036 35012
rect 20444 34960 20496 35012
rect 16488 34892 16540 34944
rect 21824 34935 21876 34944
rect 21824 34901 21833 34935
rect 21833 34901 21867 34935
rect 21867 34901 21876 34935
rect 21824 34892 21876 34901
rect 22468 34892 22520 34944
rect 25688 34892 25740 34944
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 20812 34688 20864 34740
rect 25320 34595 25372 34604
rect 25320 34561 25329 34595
rect 25329 34561 25363 34595
rect 25363 34561 25372 34595
rect 25320 34552 25372 34561
rect 21088 34348 21140 34400
rect 21364 34391 21416 34400
rect 21364 34357 21373 34391
rect 21373 34357 21407 34391
rect 21407 34357 21416 34391
rect 21364 34348 21416 34357
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 9036 34144 9088 34196
rect 11796 34008 11848 34060
rect 19708 34008 19760 34060
rect 22284 34008 22336 34060
rect 9220 33940 9272 33992
rect 19432 33983 19484 33992
rect 19432 33949 19441 33983
rect 19441 33949 19475 33983
rect 19475 33949 19484 33983
rect 19432 33940 19484 33949
rect 25320 33983 25372 33992
rect 25320 33949 25329 33983
rect 25329 33949 25363 33983
rect 25363 33949 25372 33983
rect 25320 33940 25372 33949
rect 15384 33872 15436 33924
rect 19800 33872 19852 33924
rect 21364 33872 21416 33924
rect 21180 33847 21232 33856
rect 21180 33813 21189 33847
rect 21189 33813 21223 33847
rect 21223 33813 21232 33847
rect 21180 33804 21232 33813
rect 22928 33804 22980 33856
rect 23204 33804 23256 33856
rect 23664 33847 23716 33856
rect 23664 33813 23673 33847
rect 23673 33813 23707 33847
rect 23707 33813 23716 33847
rect 23664 33804 23716 33813
rect 26240 33804 26292 33856
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 22560 33600 22612 33652
rect 23204 33600 23256 33652
rect 21364 33532 21416 33584
rect 19524 33507 19576 33516
rect 19524 33473 19533 33507
rect 19533 33473 19567 33507
rect 19567 33473 19576 33507
rect 19524 33464 19576 33473
rect 22284 33532 22336 33584
rect 23664 33532 23716 33584
rect 19800 33396 19852 33448
rect 20536 33396 20588 33448
rect 22376 33396 22428 33448
rect 22928 33396 22980 33448
rect 21364 33260 21416 33312
rect 23664 33260 23716 33312
rect 24676 33260 24728 33312
rect 24768 33260 24820 33312
rect 25964 33260 26016 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 16764 33099 16816 33108
rect 16764 33065 16773 33099
rect 16773 33065 16807 33099
rect 16807 33065 16816 33099
rect 16764 33056 16816 33065
rect 22376 33056 22428 33108
rect 22744 33056 22796 33108
rect 16120 32963 16172 32972
rect 16120 32929 16129 32963
rect 16129 32929 16163 32963
rect 16163 32929 16172 32963
rect 16580 32963 16632 32972
rect 16120 32920 16172 32929
rect 16580 32929 16589 32963
rect 16589 32929 16623 32963
rect 16623 32929 16632 32963
rect 16580 32920 16632 32929
rect 16764 32852 16816 32904
rect 17132 32852 17184 32904
rect 17868 32920 17920 32972
rect 19432 32852 19484 32904
rect 12624 32716 12676 32768
rect 17040 32716 17092 32768
rect 21824 32716 21876 32768
rect 22284 32963 22336 32972
rect 22284 32929 22293 32963
rect 22293 32929 22327 32963
rect 22327 32929 22336 32963
rect 22284 32920 22336 32929
rect 25320 32988 25372 33040
rect 25044 32963 25096 32972
rect 25044 32929 25053 32963
rect 25053 32929 25087 32963
rect 25087 32929 25096 32963
rect 25044 32920 25096 32929
rect 25228 32963 25280 32972
rect 25228 32929 25237 32963
rect 25237 32929 25271 32963
rect 25271 32929 25280 32963
rect 25228 32920 25280 32929
rect 23664 32852 23716 32904
rect 24952 32852 25004 32904
rect 25412 32852 25464 32904
rect 24676 32784 24728 32836
rect 23848 32716 23900 32768
rect 24860 32716 24912 32768
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 17040 32555 17092 32564
rect 15384 32487 15436 32496
rect 15384 32453 15393 32487
rect 15393 32453 15427 32487
rect 15427 32453 15436 32487
rect 17040 32521 17049 32555
rect 17049 32521 17083 32555
rect 17083 32521 17092 32555
rect 17040 32512 17092 32521
rect 15384 32444 15436 32453
rect 16672 32444 16724 32496
rect 23940 32512 23992 32564
rect 25320 32512 25372 32564
rect 26056 32512 26108 32564
rect 22284 32444 22336 32496
rect 13360 32308 13412 32360
rect 16764 32308 16816 32360
rect 16580 32172 16632 32224
rect 18972 32172 19024 32224
rect 21180 32308 21232 32360
rect 19432 32172 19484 32224
rect 20904 32172 20956 32224
rect 21824 32376 21876 32428
rect 24768 32444 24820 32496
rect 25228 32308 25280 32360
rect 21456 32240 21508 32292
rect 21364 32172 21416 32224
rect 21824 32172 21876 32224
rect 26516 32172 26568 32224
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 18512 31968 18564 32020
rect 18972 31968 19024 32020
rect 21456 31968 21508 32020
rect 22192 31968 22244 32020
rect 12532 31900 12584 31952
rect 16120 31875 16172 31884
rect 16120 31841 16129 31875
rect 16129 31841 16163 31875
rect 16163 31841 16172 31875
rect 16120 31832 16172 31841
rect 17684 31832 17736 31884
rect 19708 31875 19760 31884
rect 19708 31841 19717 31875
rect 19717 31841 19751 31875
rect 19751 31841 19760 31875
rect 19708 31832 19760 31841
rect 21916 31832 21968 31884
rect 16580 31764 16632 31816
rect 16764 31807 16816 31816
rect 16764 31773 16773 31807
rect 16773 31773 16807 31807
rect 16807 31773 16816 31807
rect 16764 31764 16816 31773
rect 19432 31807 19484 31816
rect 19432 31773 19441 31807
rect 19441 31773 19475 31807
rect 19475 31773 19484 31807
rect 19432 31764 19484 31773
rect 16672 31628 16724 31680
rect 21364 31696 21416 31748
rect 22560 31696 22612 31748
rect 22744 31900 22796 31952
rect 25044 31900 25096 31952
rect 23296 31832 23348 31884
rect 23020 31764 23072 31816
rect 25320 31807 25372 31816
rect 25320 31773 25329 31807
rect 25329 31773 25363 31807
rect 25363 31773 25372 31807
rect 25320 31764 25372 31773
rect 18972 31628 19024 31680
rect 20996 31628 21048 31680
rect 21640 31671 21692 31680
rect 21640 31637 21649 31671
rect 21649 31637 21683 31671
rect 21683 31637 21692 31671
rect 21640 31628 21692 31637
rect 22008 31671 22060 31680
rect 22008 31637 22017 31671
rect 22017 31637 22051 31671
rect 22051 31637 22060 31671
rect 22008 31628 22060 31637
rect 24768 31628 24820 31680
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 19708 31424 19760 31476
rect 21364 31467 21416 31476
rect 21364 31433 21373 31467
rect 21373 31433 21407 31467
rect 21407 31433 21416 31467
rect 21364 31424 21416 31433
rect 21732 31424 21784 31476
rect 22008 31424 22060 31476
rect 23572 31424 23624 31476
rect 25504 31424 25556 31476
rect 14924 31356 14976 31408
rect 18972 31356 19024 31408
rect 22652 31356 22704 31408
rect 23020 31356 23072 31408
rect 16764 31288 16816 31340
rect 20444 31331 20496 31340
rect 20444 31297 20453 31331
rect 20453 31297 20487 31331
rect 20487 31297 20496 31331
rect 20444 31288 20496 31297
rect 13360 31263 13412 31272
rect 13360 31229 13369 31263
rect 13369 31229 13403 31263
rect 13403 31229 13412 31263
rect 13360 31220 13412 31229
rect 16120 31220 16172 31272
rect 17684 31263 17736 31272
rect 17684 31229 17693 31263
rect 17693 31229 17727 31263
rect 17727 31229 17736 31263
rect 17684 31220 17736 31229
rect 18696 31220 18748 31272
rect 22284 31288 22336 31340
rect 23848 31288 23900 31340
rect 25504 31288 25556 31340
rect 25136 31220 25188 31272
rect 25872 31220 25924 31272
rect 13820 31084 13872 31136
rect 16580 31084 16632 31136
rect 16764 31127 16816 31136
rect 16764 31093 16773 31127
rect 16773 31093 16807 31127
rect 16807 31093 16816 31127
rect 16764 31084 16816 31093
rect 17500 31084 17552 31136
rect 20444 31084 20496 31136
rect 21180 31084 21232 31136
rect 23848 31084 23900 31136
rect 24768 31084 24820 31136
rect 25136 31127 25188 31136
rect 25136 31093 25145 31127
rect 25145 31093 25179 31127
rect 25179 31093 25188 31127
rect 25136 31084 25188 31093
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 10232 30880 10284 30932
rect 15384 30880 15436 30932
rect 18696 30880 18748 30932
rect 18972 30880 19024 30932
rect 22652 30880 22704 30932
rect 19432 30744 19484 30796
rect 21364 30744 21416 30796
rect 8760 30676 8812 30728
rect 14096 30676 14148 30728
rect 15384 30676 15436 30728
rect 23848 30880 23900 30932
rect 25504 30923 25556 30932
rect 25504 30889 25513 30923
rect 25513 30889 25547 30923
rect 25547 30889 25556 30923
rect 25504 30880 25556 30889
rect 15108 30651 15160 30660
rect 15108 30617 15117 30651
rect 15117 30617 15151 30651
rect 15151 30617 15160 30651
rect 15108 30608 15160 30617
rect 18972 30608 19024 30660
rect 20996 30651 21048 30660
rect 20996 30617 21005 30651
rect 21005 30617 21039 30651
rect 21039 30617 21048 30651
rect 20996 30608 21048 30617
rect 22652 30608 22704 30660
rect 18788 30540 18840 30592
rect 20076 30583 20128 30592
rect 20076 30549 20085 30583
rect 20085 30549 20119 30583
rect 20119 30549 20128 30583
rect 20076 30540 20128 30549
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 13360 30336 13412 30388
rect 16580 30336 16632 30388
rect 7656 30200 7708 30252
rect 12716 30268 12768 30320
rect 14096 30311 14148 30320
rect 14096 30277 14105 30311
rect 14105 30277 14139 30311
rect 14139 30277 14148 30311
rect 14096 30268 14148 30277
rect 14556 30268 14608 30320
rect 16856 30243 16908 30252
rect 16856 30209 16865 30243
rect 16865 30209 16899 30243
rect 16899 30209 16908 30243
rect 16856 30200 16908 30209
rect 12072 30175 12124 30184
rect 12072 30141 12081 30175
rect 12081 30141 12115 30175
rect 12115 30141 12124 30175
rect 12072 30132 12124 30141
rect 12164 30132 12216 30184
rect 12716 30132 12768 30184
rect 13360 30132 13412 30184
rect 16028 30175 16080 30184
rect 16028 30141 16037 30175
rect 16037 30141 16071 30175
rect 16071 30141 16080 30175
rect 16028 30132 16080 30141
rect 18972 30379 19024 30388
rect 18972 30345 18981 30379
rect 18981 30345 19015 30379
rect 19015 30345 19024 30379
rect 18972 30336 19024 30345
rect 20076 30336 20128 30388
rect 18328 30268 18380 30320
rect 21916 30268 21968 30320
rect 22468 30311 22520 30320
rect 22468 30277 22477 30311
rect 22477 30277 22511 30311
rect 22511 30277 22520 30311
rect 22468 30268 22520 30277
rect 22836 30268 22888 30320
rect 24860 30268 24912 30320
rect 19984 30132 20036 30184
rect 20536 30175 20588 30184
rect 20536 30141 20545 30175
rect 20545 30141 20579 30175
rect 20579 30141 20588 30175
rect 20536 30132 20588 30141
rect 8944 30107 8996 30116
rect 8944 30073 8953 30107
rect 8953 30073 8987 30107
rect 8987 30073 8996 30107
rect 8944 30064 8996 30073
rect 16488 30064 16540 30116
rect 22100 30064 22152 30116
rect 11520 29996 11572 30048
rect 13636 29996 13688 30048
rect 15936 29996 15988 30048
rect 19800 29996 19852 30048
rect 21916 29996 21968 30048
rect 22836 30132 22888 30184
rect 23572 30175 23624 30184
rect 23572 30141 23581 30175
rect 23581 30141 23615 30175
rect 23615 30141 23624 30175
rect 23572 30132 23624 30141
rect 25228 30132 25280 30184
rect 26148 30064 26200 30116
rect 24860 29996 24912 30048
rect 25228 29996 25280 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 12072 29792 12124 29844
rect 13820 29792 13872 29844
rect 11428 29656 11480 29708
rect 13360 29656 13412 29708
rect 16028 29656 16080 29708
rect 15660 29588 15712 29640
rect 16488 29767 16540 29776
rect 16488 29733 16497 29767
rect 16497 29733 16531 29767
rect 16531 29733 16540 29767
rect 16488 29724 16540 29733
rect 18420 29724 18472 29776
rect 19340 29656 19392 29708
rect 11336 29520 11388 29572
rect 12716 29520 12768 29572
rect 14924 29452 14976 29504
rect 15200 29495 15252 29504
rect 15200 29461 15209 29495
rect 15209 29461 15243 29495
rect 15243 29461 15252 29495
rect 15200 29452 15252 29461
rect 16120 29452 16172 29504
rect 16488 29452 16540 29504
rect 18328 29520 18380 29572
rect 18880 29588 18932 29640
rect 26148 29792 26200 29844
rect 23388 29724 23440 29776
rect 26608 29656 26660 29708
rect 20812 29588 20864 29640
rect 24492 29588 24544 29640
rect 25320 29631 25372 29640
rect 25320 29597 25329 29631
rect 25329 29597 25363 29631
rect 25363 29597 25372 29631
rect 25320 29588 25372 29597
rect 24860 29520 24912 29572
rect 18788 29495 18840 29504
rect 18788 29461 18797 29495
rect 18797 29461 18831 29495
rect 18831 29461 18840 29495
rect 18788 29452 18840 29461
rect 19156 29452 19208 29504
rect 19984 29452 20036 29504
rect 22468 29452 22520 29504
rect 24492 29495 24544 29504
rect 24492 29461 24501 29495
rect 24501 29461 24535 29495
rect 24535 29461 24544 29495
rect 24492 29452 24544 29461
rect 25228 29452 25280 29504
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 8852 29248 8904 29300
rect 10416 29248 10468 29300
rect 12440 29248 12492 29300
rect 12624 29291 12676 29300
rect 12624 29257 12633 29291
rect 12633 29257 12667 29291
rect 12667 29257 12676 29291
rect 12624 29248 12676 29257
rect 13820 29248 13872 29300
rect 13912 29248 13964 29300
rect 9680 29180 9732 29232
rect 10876 29044 10928 29096
rect 11796 29044 11848 29096
rect 14924 29180 14976 29232
rect 13360 29155 13412 29164
rect 13360 29121 13369 29155
rect 13369 29121 13403 29155
rect 13403 29121 13412 29155
rect 13360 29112 13412 29121
rect 15200 29248 15252 29300
rect 17500 29248 17552 29300
rect 17868 29248 17920 29300
rect 19156 29291 19208 29300
rect 19156 29257 19165 29291
rect 19165 29257 19199 29291
rect 19199 29257 19208 29291
rect 19156 29248 19208 29257
rect 20628 29248 20680 29300
rect 15936 29223 15988 29232
rect 15936 29189 15945 29223
rect 15945 29189 15979 29223
rect 15979 29189 15988 29223
rect 15936 29180 15988 29189
rect 17040 29180 17092 29232
rect 19984 29223 20036 29232
rect 19984 29189 19993 29223
rect 19993 29189 20027 29223
rect 20027 29189 20036 29223
rect 19984 29180 20036 29189
rect 20352 29180 20404 29232
rect 24124 29248 24176 29300
rect 24584 29248 24636 29300
rect 25320 29248 25372 29300
rect 17408 29112 17460 29164
rect 13636 29044 13688 29096
rect 17868 29112 17920 29164
rect 20904 29044 20956 29096
rect 10232 28976 10284 29028
rect 12164 29019 12216 29028
rect 12164 28985 12173 29019
rect 12173 28985 12207 29019
rect 12207 28985 12216 29019
rect 12164 28976 12216 28985
rect 14648 28976 14700 29028
rect 15752 28976 15804 29028
rect 14096 28908 14148 28960
rect 15292 28908 15344 28960
rect 21824 29019 21876 29028
rect 21824 28985 21833 29019
rect 21833 28985 21867 29019
rect 21867 28985 21876 29019
rect 25412 29112 25464 29164
rect 22836 29044 22888 29096
rect 23756 29044 23808 29096
rect 24952 29044 25004 29096
rect 21824 28976 21876 28985
rect 24676 28976 24728 29028
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 10876 28747 10928 28756
rect 10876 28713 10885 28747
rect 10885 28713 10919 28747
rect 10919 28713 10928 28747
rect 10876 28704 10928 28713
rect 11428 28611 11480 28620
rect 11428 28577 11437 28611
rect 11437 28577 11471 28611
rect 11471 28577 11480 28611
rect 11428 28568 11480 28577
rect 11704 28568 11756 28620
rect 12716 28568 12768 28620
rect 13728 28704 13780 28756
rect 14924 28704 14976 28756
rect 18880 28747 18932 28756
rect 18880 28713 18889 28747
rect 18889 28713 18923 28747
rect 18923 28713 18932 28747
rect 18880 28704 18932 28713
rect 23756 28704 23808 28756
rect 14096 28568 14148 28620
rect 16488 28636 16540 28688
rect 15384 28611 15436 28620
rect 15384 28577 15393 28611
rect 15393 28577 15427 28611
rect 15427 28577 15436 28611
rect 15384 28568 15436 28577
rect 18972 28568 19024 28620
rect 20996 28568 21048 28620
rect 21364 28568 21416 28620
rect 22192 28568 22244 28620
rect 24768 28636 24820 28688
rect 23664 28568 23716 28620
rect 24860 28568 24912 28620
rect 26056 28568 26108 28620
rect 15108 28500 15160 28552
rect 19340 28500 19392 28552
rect 20628 28543 20680 28552
rect 20628 28509 20637 28543
rect 20637 28509 20671 28543
rect 20671 28509 20680 28543
rect 20628 28500 20680 28509
rect 22284 28500 22336 28552
rect 22560 28500 22612 28552
rect 24952 28543 25004 28552
rect 24952 28509 24961 28543
rect 24961 28509 24995 28543
rect 24995 28509 25004 28543
rect 24952 28500 25004 28509
rect 9680 28432 9732 28484
rect 11612 28432 11664 28484
rect 11520 28364 11572 28416
rect 16304 28432 16356 28484
rect 18880 28432 18932 28484
rect 20904 28475 20956 28484
rect 20904 28441 20913 28475
rect 20913 28441 20947 28475
rect 20947 28441 20956 28475
rect 20904 28432 20956 28441
rect 14832 28407 14884 28416
rect 14832 28373 14841 28407
rect 14841 28373 14875 28407
rect 14875 28373 14884 28407
rect 14832 28364 14884 28373
rect 16028 28407 16080 28416
rect 16028 28373 16037 28407
rect 16037 28373 16071 28407
rect 16071 28373 16080 28407
rect 16028 28364 16080 28373
rect 16488 28364 16540 28416
rect 18696 28364 18748 28416
rect 19708 28364 19760 28416
rect 21640 28364 21692 28416
rect 21732 28364 21784 28416
rect 25964 28432 26016 28484
rect 23940 28407 23992 28416
rect 23940 28373 23949 28407
rect 23949 28373 23983 28407
rect 23983 28373 23992 28407
rect 23940 28364 23992 28373
rect 24400 28364 24452 28416
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 11612 28160 11664 28212
rect 13728 28203 13780 28212
rect 13728 28169 13737 28203
rect 13737 28169 13771 28203
rect 13771 28169 13780 28203
rect 13728 28160 13780 28169
rect 15568 28203 15620 28212
rect 15568 28169 15577 28203
rect 15577 28169 15611 28203
rect 15611 28169 15620 28203
rect 15568 28160 15620 28169
rect 18880 28160 18932 28212
rect 19708 28203 19760 28212
rect 19708 28169 19717 28203
rect 19717 28169 19751 28203
rect 19751 28169 19760 28203
rect 19708 28160 19760 28169
rect 13452 28092 13504 28144
rect 22192 28160 22244 28212
rect 26240 28160 26292 28212
rect 20628 28092 20680 28144
rect 11060 28024 11112 28076
rect 16304 28024 16356 28076
rect 16672 28024 16724 28076
rect 18788 28024 18840 28076
rect 11704 27999 11756 28008
rect 11704 27965 11713 27999
rect 11713 27965 11747 27999
rect 11747 27965 11756 27999
rect 11704 27956 11756 27965
rect 10784 27888 10836 27940
rect 15384 27888 15436 27940
rect 16764 27956 16816 28008
rect 13820 27820 13872 27872
rect 16304 27863 16356 27872
rect 16304 27829 16313 27863
rect 16313 27829 16347 27863
rect 16347 27829 16356 27863
rect 16304 27820 16356 27829
rect 16856 27863 16908 27872
rect 16856 27829 16865 27863
rect 16865 27829 16899 27863
rect 16899 27829 16908 27863
rect 16856 27820 16908 27829
rect 17408 27999 17460 28008
rect 17408 27965 17417 27999
rect 17417 27965 17451 27999
rect 17451 27965 17460 27999
rect 17408 27956 17460 27965
rect 17960 27956 18012 28008
rect 17684 27888 17736 27940
rect 21824 28024 21876 28076
rect 18512 27863 18564 27872
rect 18512 27829 18521 27863
rect 18521 27829 18555 27863
rect 18555 27829 18564 27863
rect 18512 27820 18564 27829
rect 18788 27863 18840 27872
rect 18788 27829 18797 27863
rect 18797 27829 18831 27863
rect 18831 27829 18840 27863
rect 18788 27820 18840 27829
rect 19156 27820 19208 27872
rect 22100 27888 22152 27940
rect 22836 27956 22888 28008
rect 23480 27999 23532 28008
rect 23480 27965 23489 27999
rect 23489 27965 23523 27999
rect 23523 27965 23532 27999
rect 23480 27956 23532 27965
rect 23940 27956 23992 28008
rect 22376 27820 22428 27872
rect 22560 27820 22612 27872
rect 25228 27863 25280 27872
rect 25228 27829 25237 27863
rect 25237 27829 25271 27863
rect 25271 27829 25280 27863
rect 25228 27820 25280 27829
rect 25412 27863 25464 27872
rect 25412 27829 25421 27863
rect 25421 27829 25455 27863
rect 25455 27829 25464 27863
rect 25412 27820 25464 27829
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 11428 27616 11480 27668
rect 12716 27616 12768 27668
rect 15108 27616 15160 27668
rect 18880 27616 18932 27668
rect 19984 27616 20036 27668
rect 23664 27616 23716 27668
rect 10784 27523 10836 27532
rect 10784 27489 10793 27523
rect 10793 27489 10827 27523
rect 10827 27489 10836 27523
rect 10784 27480 10836 27489
rect 13084 27548 13136 27600
rect 16120 27548 16172 27600
rect 23480 27548 23532 27600
rect 24768 27548 24820 27600
rect 9312 27276 9364 27328
rect 15108 27480 15160 27532
rect 17776 27480 17828 27532
rect 22836 27480 22888 27532
rect 24124 27523 24176 27532
rect 24124 27489 24133 27523
rect 24133 27489 24167 27523
rect 24167 27489 24176 27523
rect 24124 27480 24176 27489
rect 25044 27523 25096 27532
rect 25044 27489 25053 27523
rect 25053 27489 25087 27523
rect 25087 27489 25096 27523
rect 25044 27480 25096 27489
rect 14832 27412 14884 27464
rect 17960 27412 18012 27464
rect 23940 27412 23992 27464
rect 25412 27412 25464 27464
rect 13820 27344 13872 27396
rect 12624 27276 12676 27328
rect 13728 27276 13780 27328
rect 15476 27276 15528 27328
rect 16028 27344 16080 27396
rect 20076 27344 20128 27396
rect 22376 27387 22428 27396
rect 22376 27353 22385 27387
rect 22385 27353 22419 27387
rect 22419 27353 22428 27387
rect 22376 27344 22428 27353
rect 23664 27344 23716 27396
rect 16488 27319 16540 27328
rect 16488 27285 16497 27319
rect 16497 27285 16531 27319
rect 16531 27285 16540 27319
rect 16488 27276 16540 27285
rect 17592 27276 17644 27328
rect 21640 27319 21692 27328
rect 21640 27285 21649 27319
rect 21649 27285 21683 27319
rect 21683 27285 21692 27319
rect 21640 27276 21692 27285
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 9772 27072 9824 27124
rect 10876 27072 10928 27124
rect 11704 27072 11756 27124
rect 11152 27004 11204 27056
rect 12716 27072 12768 27124
rect 13636 27004 13688 27056
rect 15200 27072 15252 27124
rect 16856 27072 16908 27124
rect 15752 27047 15804 27056
rect 15752 27013 15761 27047
rect 15761 27013 15795 27047
rect 15795 27013 15804 27047
rect 15752 27004 15804 27013
rect 19248 27072 19300 27124
rect 19984 27115 20036 27124
rect 19984 27081 19993 27115
rect 19993 27081 20027 27115
rect 20027 27081 20036 27115
rect 19984 27072 20036 27081
rect 22744 27072 22796 27124
rect 24768 27072 24820 27124
rect 11704 26936 11756 26988
rect 12808 26936 12860 26988
rect 13084 26979 13136 26988
rect 13084 26945 13093 26979
rect 13093 26945 13127 26979
rect 13127 26945 13136 26979
rect 13084 26936 13136 26945
rect 14832 26936 14884 26988
rect 16580 26936 16632 26988
rect 18880 27004 18932 27056
rect 22928 27004 22980 27056
rect 25228 27004 25280 27056
rect 26240 27004 26292 27056
rect 22652 26936 22704 26988
rect 23296 26936 23348 26988
rect 11336 26868 11388 26920
rect 9312 26800 9364 26852
rect 13452 26868 13504 26920
rect 22100 26868 22152 26920
rect 23480 26868 23532 26920
rect 25596 26868 25648 26920
rect 3424 26732 3476 26784
rect 11980 26732 12032 26784
rect 14924 26732 14976 26784
rect 18972 26732 19024 26784
rect 21824 26775 21876 26784
rect 21824 26741 21833 26775
rect 21833 26741 21867 26775
rect 21867 26741 21876 26775
rect 21824 26732 21876 26741
rect 22376 26775 22428 26784
rect 22376 26741 22385 26775
rect 22385 26741 22419 26775
rect 22419 26741 22428 26775
rect 22376 26732 22428 26741
rect 24860 26732 24912 26784
rect 25964 26732 26016 26784
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 11152 26571 11204 26580
rect 11152 26537 11161 26571
rect 11161 26537 11195 26571
rect 11195 26537 11204 26571
rect 11152 26528 11204 26537
rect 13636 26528 13688 26580
rect 16028 26528 16080 26580
rect 17040 26528 17092 26580
rect 17592 26528 17644 26580
rect 19892 26528 19944 26580
rect 20076 26528 20128 26580
rect 9772 26392 9824 26444
rect 11060 26392 11112 26444
rect 11612 26460 11664 26512
rect 22100 26528 22152 26580
rect 22284 26571 22336 26580
rect 22284 26537 22293 26571
rect 22293 26537 22327 26571
rect 22327 26537 22336 26571
rect 22284 26528 22336 26537
rect 24952 26528 25004 26580
rect 8576 26256 8628 26308
rect 11796 26256 11848 26308
rect 15016 26392 15068 26444
rect 15200 26392 15252 26444
rect 14556 26324 14608 26376
rect 15108 26324 15160 26376
rect 16580 26392 16632 26444
rect 21088 26460 21140 26512
rect 21824 26460 21876 26512
rect 16948 26324 17000 26376
rect 17408 26392 17460 26444
rect 19432 26435 19484 26444
rect 19432 26401 19441 26435
rect 19441 26401 19475 26435
rect 19475 26401 19484 26435
rect 19432 26392 19484 26401
rect 20996 26392 21048 26444
rect 21640 26392 21692 26444
rect 14832 26256 14884 26308
rect 15568 26256 15620 26308
rect 16028 26299 16080 26308
rect 16028 26265 16037 26299
rect 16037 26265 16071 26299
rect 16071 26265 16080 26299
rect 16028 26256 16080 26265
rect 16304 26256 16356 26308
rect 17224 26324 17276 26376
rect 22560 26460 22612 26512
rect 25044 26460 25096 26512
rect 22284 26392 22336 26444
rect 22744 26324 22796 26376
rect 23388 26324 23440 26376
rect 24032 26367 24084 26376
rect 24032 26333 24041 26367
rect 24041 26333 24075 26367
rect 24075 26333 24084 26367
rect 24032 26324 24084 26333
rect 24860 26324 24912 26376
rect 25136 26392 25188 26444
rect 25228 26435 25280 26444
rect 25228 26401 25237 26435
rect 25237 26401 25271 26435
rect 25271 26401 25280 26435
rect 25228 26392 25280 26401
rect 25412 26392 25464 26444
rect 19984 26256 20036 26308
rect 25136 26256 25188 26308
rect 25872 26324 25924 26376
rect 25596 26256 25648 26308
rect 18328 26188 18380 26240
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 12624 26027 12676 26036
rect 12624 25993 12633 26027
rect 12633 25993 12667 26027
rect 12667 25993 12676 26027
rect 12624 25984 12676 25993
rect 14648 25984 14700 26036
rect 10692 25916 10744 25968
rect 14188 25916 14240 25968
rect 16304 25984 16356 26036
rect 18328 25984 18380 26036
rect 18880 25984 18932 26036
rect 20168 25984 20220 26036
rect 22468 26027 22520 26036
rect 22468 25993 22477 26027
rect 22477 25993 22511 26027
rect 22511 25993 22520 26027
rect 22468 25984 22520 25993
rect 17592 25916 17644 25968
rect 18420 25916 18472 25968
rect 25136 25984 25188 26036
rect 12532 25891 12584 25900
rect 12532 25857 12541 25891
rect 12541 25857 12575 25891
rect 12575 25857 12584 25891
rect 12532 25848 12584 25857
rect 24860 25916 24912 25968
rect 11336 25780 11388 25832
rect 14096 25823 14148 25832
rect 14096 25789 14105 25823
rect 14105 25789 14139 25823
rect 14139 25789 14148 25823
rect 14096 25780 14148 25789
rect 15384 25823 15436 25832
rect 15384 25789 15393 25823
rect 15393 25789 15427 25823
rect 15427 25789 15436 25823
rect 15384 25780 15436 25789
rect 18604 25780 18656 25832
rect 14832 25644 14884 25696
rect 15016 25644 15068 25696
rect 17776 25712 17828 25764
rect 16856 25687 16908 25696
rect 16856 25653 16865 25687
rect 16865 25653 16899 25687
rect 16899 25653 16908 25687
rect 16856 25644 16908 25653
rect 21180 25644 21232 25696
rect 23940 25891 23992 25900
rect 23940 25857 23949 25891
rect 23949 25857 23983 25891
rect 23983 25857 23992 25891
rect 23940 25848 23992 25857
rect 23388 25780 23440 25832
rect 25136 25823 25188 25832
rect 25136 25789 25145 25823
rect 25145 25789 25179 25823
rect 25179 25789 25188 25823
rect 25136 25780 25188 25789
rect 22376 25712 22428 25764
rect 22836 25712 22888 25764
rect 21640 25644 21692 25696
rect 22468 25644 22520 25696
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 11704 25440 11756 25492
rect 16488 25440 16540 25492
rect 18880 25440 18932 25492
rect 20260 25483 20312 25492
rect 20260 25449 20269 25483
rect 20269 25449 20303 25483
rect 20303 25449 20312 25483
rect 20260 25440 20312 25449
rect 23940 25440 23992 25492
rect 24032 25440 24084 25492
rect 12716 25372 12768 25424
rect 10876 25347 10928 25356
rect 10876 25313 10885 25347
rect 10885 25313 10919 25347
rect 10919 25313 10928 25347
rect 10876 25304 10928 25313
rect 14556 25304 14608 25356
rect 14648 25304 14700 25356
rect 14832 25347 14884 25356
rect 14832 25313 14841 25347
rect 14841 25313 14875 25347
rect 14875 25313 14884 25347
rect 14832 25304 14884 25313
rect 12716 25236 12768 25288
rect 13360 25236 13412 25288
rect 16856 25304 16908 25356
rect 15200 25236 15252 25288
rect 17776 25279 17828 25288
rect 17776 25245 17785 25279
rect 17785 25245 17819 25279
rect 17819 25245 17828 25279
rect 17776 25236 17828 25245
rect 18328 25236 18380 25288
rect 20260 25236 20312 25288
rect 24860 25372 24912 25424
rect 22376 25304 22428 25356
rect 10324 25100 10376 25152
rect 15384 25168 15436 25220
rect 16396 25168 16448 25220
rect 12624 25143 12676 25152
rect 12624 25109 12633 25143
rect 12633 25109 12667 25143
rect 12667 25109 12676 25143
rect 12624 25100 12676 25109
rect 15660 25100 15712 25152
rect 15752 25143 15804 25152
rect 15752 25109 15761 25143
rect 15761 25109 15795 25143
rect 15795 25109 15804 25143
rect 15752 25100 15804 25109
rect 16488 25100 16540 25152
rect 19064 25168 19116 25220
rect 19340 25211 19392 25220
rect 19340 25177 19349 25211
rect 19349 25177 19383 25211
rect 19383 25177 19392 25211
rect 19340 25168 19392 25177
rect 20076 25168 20128 25220
rect 25320 25279 25372 25288
rect 25320 25245 25329 25279
rect 25329 25245 25363 25279
rect 25363 25245 25372 25279
rect 25320 25236 25372 25245
rect 18512 25100 18564 25152
rect 19892 25143 19944 25152
rect 19892 25109 19901 25143
rect 19901 25109 19935 25143
rect 19935 25109 19944 25143
rect 19892 25100 19944 25109
rect 23848 25211 23900 25220
rect 23848 25177 23857 25211
rect 23857 25177 23891 25211
rect 23891 25177 23900 25211
rect 23848 25168 23900 25177
rect 26056 25168 26108 25220
rect 25136 25100 25188 25152
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 7564 24896 7616 24948
rect 9404 24828 9456 24880
rect 11152 24896 11204 24948
rect 14832 24896 14884 24948
rect 15660 24896 15712 24948
rect 16396 24896 16448 24948
rect 18328 24896 18380 24948
rect 18788 24896 18840 24948
rect 19340 24896 19392 24948
rect 12716 24828 12768 24880
rect 13544 24828 13596 24880
rect 14648 24828 14700 24880
rect 15936 24828 15988 24880
rect 17040 24828 17092 24880
rect 12164 24803 12216 24812
rect 12164 24769 12173 24803
rect 12173 24769 12207 24803
rect 12207 24769 12216 24803
rect 12164 24760 12216 24769
rect 12808 24760 12860 24812
rect 18880 24828 18932 24880
rect 24124 24828 24176 24880
rect 25136 24828 25188 24880
rect 10876 24692 10928 24744
rect 11060 24692 11112 24744
rect 13912 24692 13964 24744
rect 14556 24692 14608 24744
rect 15016 24692 15068 24744
rect 18328 24760 18380 24812
rect 19432 24760 19484 24812
rect 21088 24760 21140 24812
rect 23296 24760 23348 24812
rect 18144 24692 18196 24744
rect 11060 24556 11112 24608
rect 11152 24599 11204 24608
rect 11152 24565 11161 24599
rect 11161 24565 11195 24599
rect 11195 24565 11204 24599
rect 11152 24556 11204 24565
rect 15200 24624 15252 24676
rect 17040 24624 17092 24676
rect 20444 24692 20496 24744
rect 22284 24692 22336 24744
rect 22652 24735 22704 24744
rect 22652 24701 22661 24735
rect 22661 24701 22695 24735
rect 22695 24701 22704 24735
rect 22652 24692 22704 24701
rect 25136 24692 25188 24744
rect 23572 24624 23624 24676
rect 15108 24556 15160 24608
rect 15568 24556 15620 24608
rect 17868 24556 17920 24608
rect 18144 24556 18196 24608
rect 18696 24556 18748 24608
rect 22100 24599 22152 24608
rect 22100 24565 22109 24599
rect 22109 24565 22143 24599
rect 22143 24565 22152 24599
rect 22100 24556 22152 24565
rect 25228 24556 25280 24608
rect 25412 24556 25464 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 9496 24216 9548 24268
rect 12624 24352 12676 24404
rect 12900 24352 12952 24404
rect 13544 24352 13596 24404
rect 15108 24352 15160 24404
rect 20444 24352 20496 24404
rect 25320 24395 25372 24404
rect 25320 24361 25329 24395
rect 25329 24361 25363 24395
rect 25363 24361 25372 24395
rect 25320 24352 25372 24361
rect 26056 24352 26108 24404
rect 19156 24284 19208 24336
rect 21088 24284 21140 24336
rect 21456 24284 21508 24336
rect 23296 24284 23348 24336
rect 25412 24284 25464 24336
rect 25964 24284 26016 24336
rect 11060 24216 11112 24268
rect 12348 24216 12400 24268
rect 18972 24216 19024 24268
rect 19432 24259 19484 24268
rect 19432 24225 19441 24259
rect 19441 24225 19475 24259
rect 19475 24225 19484 24259
rect 19432 24216 19484 24225
rect 7840 24148 7892 24200
rect 17684 24191 17736 24200
rect 17684 24157 17693 24191
rect 17693 24157 17727 24191
rect 17727 24157 17736 24191
rect 17684 24148 17736 24157
rect 18512 24191 18564 24200
rect 18512 24157 18521 24191
rect 18521 24157 18555 24191
rect 18555 24157 18564 24191
rect 18512 24148 18564 24157
rect 19248 24148 19300 24200
rect 22192 24216 22244 24268
rect 24124 24216 24176 24268
rect 9404 24080 9456 24132
rect 10876 24055 10928 24064
rect 10876 24021 10885 24055
rect 10885 24021 10919 24055
rect 10919 24021 10928 24055
rect 10876 24012 10928 24021
rect 11980 24080 12032 24132
rect 12716 24080 12768 24132
rect 18880 24080 18932 24132
rect 13912 24012 13964 24064
rect 16580 24012 16632 24064
rect 18788 24012 18840 24064
rect 22284 24080 22336 24132
rect 19892 24012 19944 24064
rect 23572 24012 23624 24064
rect 24952 24012 25004 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 9680 23808 9732 23860
rect 7840 23672 7892 23724
rect 9404 23672 9456 23724
rect 10416 23851 10468 23860
rect 10416 23817 10425 23851
rect 10425 23817 10459 23851
rect 10459 23817 10468 23851
rect 10416 23808 10468 23817
rect 14188 23808 14240 23860
rect 14924 23851 14976 23860
rect 14924 23817 14933 23851
rect 14933 23817 14967 23851
rect 14967 23817 14976 23851
rect 14924 23808 14976 23817
rect 16580 23808 16632 23860
rect 17776 23808 17828 23860
rect 13636 23783 13688 23792
rect 13636 23749 13645 23783
rect 13645 23749 13679 23783
rect 13679 23749 13688 23783
rect 13636 23740 13688 23749
rect 13728 23783 13780 23792
rect 13728 23749 13737 23783
rect 13737 23749 13771 23783
rect 13771 23749 13780 23783
rect 13728 23740 13780 23749
rect 15844 23740 15896 23792
rect 18788 23808 18840 23860
rect 18880 23851 18932 23860
rect 18880 23817 18889 23851
rect 18889 23817 18923 23851
rect 18923 23817 18932 23851
rect 18880 23808 18932 23817
rect 19064 23808 19116 23860
rect 25136 23808 25188 23860
rect 25412 23851 25464 23860
rect 25412 23817 25421 23851
rect 25421 23817 25455 23851
rect 25455 23817 25464 23851
rect 25412 23808 25464 23817
rect 14004 23672 14056 23724
rect 10048 23604 10100 23656
rect 10968 23647 11020 23656
rect 10968 23613 10977 23647
rect 10977 23613 11011 23647
rect 11011 23613 11020 23647
rect 10968 23604 11020 23613
rect 10324 23536 10376 23588
rect 12900 23536 12952 23588
rect 13912 23604 13964 23656
rect 15660 23647 15712 23656
rect 15660 23613 15669 23647
rect 15669 23613 15703 23647
rect 15703 23613 15712 23647
rect 15660 23604 15712 23613
rect 19616 23715 19668 23724
rect 19616 23681 19625 23715
rect 19625 23681 19659 23715
rect 19659 23681 19668 23715
rect 19616 23672 19668 23681
rect 19524 23604 19576 23656
rect 20352 23672 20404 23724
rect 20812 23715 20864 23724
rect 20812 23681 20821 23715
rect 20821 23681 20855 23715
rect 20855 23681 20864 23715
rect 20812 23672 20864 23681
rect 21364 23672 21416 23724
rect 21456 23715 21508 23724
rect 21456 23681 21465 23715
rect 21465 23681 21499 23715
rect 21499 23681 21508 23715
rect 21456 23672 21508 23681
rect 22008 23672 22060 23724
rect 19892 23647 19944 23656
rect 19892 23613 19901 23647
rect 19901 23613 19935 23647
rect 19935 23613 19944 23647
rect 19892 23604 19944 23613
rect 20996 23647 21048 23656
rect 20996 23613 21005 23647
rect 21005 23613 21039 23647
rect 21039 23613 21048 23647
rect 20996 23604 21048 23613
rect 23388 23740 23440 23792
rect 26056 23740 26108 23792
rect 23204 23715 23256 23724
rect 23204 23681 23213 23715
rect 23213 23681 23247 23715
rect 23247 23681 23256 23715
rect 23204 23672 23256 23681
rect 24952 23672 25004 23724
rect 23572 23604 23624 23656
rect 22100 23536 22152 23588
rect 22284 23536 22336 23588
rect 9404 23468 9456 23520
rect 10876 23468 10928 23520
rect 12624 23468 12676 23520
rect 12808 23468 12860 23520
rect 17316 23468 17368 23520
rect 17776 23468 17828 23520
rect 19064 23468 19116 23520
rect 19248 23511 19300 23520
rect 19248 23477 19257 23511
rect 19257 23477 19291 23511
rect 19291 23477 19300 23511
rect 19248 23468 19300 23477
rect 19340 23468 19392 23520
rect 23940 23468 23992 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 9220 23264 9272 23316
rect 10140 23264 10192 23316
rect 15200 23264 15252 23316
rect 9404 23196 9456 23248
rect 8668 23128 8720 23180
rect 10324 23128 10376 23180
rect 10600 23128 10652 23180
rect 11704 23171 11756 23180
rect 11704 23137 11713 23171
rect 11713 23137 11747 23171
rect 11747 23137 11756 23171
rect 11704 23128 11756 23137
rect 11796 23171 11848 23180
rect 11796 23137 11805 23171
rect 11805 23137 11839 23171
rect 11839 23137 11848 23171
rect 11796 23128 11848 23137
rect 12716 23196 12768 23248
rect 10784 23060 10836 23112
rect 11612 23103 11664 23112
rect 11612 23069 11621 23103
rect 11621 23069 11655 23103
rect 11655 23069 11664 23103
rect 11612 23060 11664 23069
rect 14188 23060 14240 23112
rect 10416 22992 10468 23044
rect 14096 22992 14148 23044
rect 15660 23060 15712 23112
rect 17132 23264 17184 23316
rect 19524 23264 19576 23316
rect 18880 23196 18932 23248
rect 18420 23171 18472 23180
rect 18420 23137 18429 23171
rect 18429 23137 18463 23171
rect 18463 23137 18472 23171
rect 18420 23128 18472 23137
rect 20444 23128 20496 23180
rect 20812 23128 20864 23180
rect 25872 23196 25924 23248
rect 25320 23128 25372 23180
rect 18328 23060 18380 23112
rect 19248 23060 19300 23112
rect 21640 23060 21692 23112
rect 16856 22992 16908 23044
rect 23756 23060 23808 23112
rect 25412 23060 25464 23112
rect 25872 22992 25924 23044
rect 10508 22924 10560 22976
rect 12164 22924 12216 22976
rect 17776 22924 17828 22976
rect 18696 22924 18748 22976
rect 18972 22924 19024 22976
rect 22100 22924 22152 22976
rect 24584 22967 24636 22976
rect 24584 22933 24593 22967
rect 24593 22933 24627 22967
rect 24627 22933 24636 22967
rect 24584 22924 24636 22933
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 11336 22720 11388 22772
rect 14096 22720 14148 22772
rect 14188 22720 14240 22772
rect 14740 22720 14792 22772
rect 16856 22763 16908 22772
rect 16856 22729 16865 22763
rect 16865 22729 16899 22763
rect 16899 22729 16908 22763
rect 16856 22720 16908 22729
rect 18328 22720 18380 22772
rect 15108 22652 15160 22704
rect 19064 22720 19116 22772
rect 19248 22720 19300 22772
rect 19616 22720 19668 22772
rect 22376 22720 22428 22772
rect 20812 22652 20864 22704
rect 7840 22584 7892 22636
rect 9496 22584 9548 22636
rect 12348 22627 12400 22636
rect 12348 22593 12357 22627
rect 12357 22593 12391 22627
rect 12391 22593 12400 22627
rect 12348 22584 12400 22593
rect 13912 22584 13964 22636
rect 18696 22584 18748 22636
rect 20904 22584 20956 22636
rect 21088 22627 21140 22636
rect 21088 22593 21097 22627
rect 21097 22593 21131 22627
rect 21131 22593 21140 22627
rect 21088 22584 21140 22593
rect 22100 22627 22152 22636
rect 22100 22593 22109 22627
rect 22109 22593 22143 22627
rect 22143 22593 22152 22627
rect 22100 22584 22152 22593
rect 23940 22627 23992 22636
rect 23940 22593 23949 22627
rect 23949 22593 23983 22627
rect 23983 22593 23992 22627
rect 23940 22584 23992 22593
rect 11152 22516 11204 22568
rect 13360 22516 13412 22568
rect 20168 22516 20220 22568
rect 23296 22559 23348 22568
rect 23296 22525 23305 22559
rect 23305 22525 23339 22559
rect 23339 22525 23348 22559
rect 23296 22516 23348 22525
rect 24768 22559 24820 22568
rect 24768 22525 24777 22559
rect 24777 22525 24811 22559
rect 24811 22525 24820 22559
rect 24768 22516 24820 22525
rect 6920 22380 6972 22432
rect 11796 22448 11848 22500
rect 15200 22448 15252 22500
rect 21088 22448 21140 22500
rect 14096 22423 14148 22432
rect 14096 22389 14105 22423
rect 14105 22389 14139 22423
rect 14139 22389 14148 22423
rect 14096 22380 14148 22389
rect 20720 22423 20772 22432
rect 20720 22389 20729 22423
rect 20729 22389 20763 22423
rect 20763 22389 20772 22423
rect 20720 22380 20772 22389
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 13912 22176 13964 22228
rect 22008 22176 22060 22228
rect 11520 22108 11572 22160
rect 9220 21972 9272 22024
rect 12808 22108 12860 22160
rect 12624 22083 12676 22092
rect 12624 22049 12633 22083
rect 12633 22049 12667 22083
rect 12667 22049 12676 22083
rect 12624 22040 12676 22049
rect 15752 22108 15804 22160
rect 8300 21836 8352 21888
rect 9496 21836 9548 21888
rect 10324 21879 10376 21888
rect 10324 21845 10333 21879
rect 10333 21845 10367 21879
rect 10367 21845 10376 21879
rect 10324 21836 10376 21845
rect 10692 21879 10744 21888
rect 10692 21845 10701 21879
rect 10701 21845 10735 21879
rect 10735 21845 10744 21879
rect 10692 21836 10744 21845
rect 11060 21879 11112 21888
rect 11060 21845 11069 21879
rect 11069 21845 11103 21879
rect 11103 21845 11112 21879
rect 11060 21836 11112 21845
rect 14096 21972 14148 22024
rect 16948 22040 17000 22092
rect 20352 22083 20404 22092
rect 20352 22049 20361 22083
rect 20361 22049 20395 22083
rect 20395 22049 20404 22083
rect 20352 22040 20404 22049
rect 22192 22040 22244 22092
rect 23388 22176 23440 22228
rect 23756 22219 23808 22228
rect 23756 22185 23765 22219
rect 23765 22185 23799 22219
rect 23799 22185 23808 22219
rect 23756 22176 23808 22185
rect 25228 22176 25280 22228
rect 23204 22108 23256 22160
rect 25044 22083 25096 22092
rect 25044 22049 25053 22083
rect 25053 22049 25087 22083
rect 25087 22049 25096 22083
rect 25044 22040 25096 22049
rect 14832 21879 14884 21888
rect 14832 21845 14841 21879
rect 14841 21845 14875 21879
rect 14875 21845 14884 21879
rect 14832 21836 14884 21845
rect 15200 21879 15252 21888
rect 15200 21845 15209 21879
rect 15209 21845 15243 21879
rect 15243 21845 15252 21879
rect 15200 21836 15252 21845
rect 16488 21904 16540 21956
rect 16580 21836 16632 21888
rect 16948 21904 17000 21956
rect 17040 21836 17092 21888
rect 17132 21836 17184 21888
rect 21180 21904 21232 21956
rect 22100 21904 22152 21956
rect 22284 21904 22336 21956
rect 20076 21879 20128 21888
rect 20076 21845 20085 21879
rect 20085 21845 20119 21879
rect 20119 21845 20128 21879
rect 20076 21836 20128 21845
rect 20260 21836 20312 21888
rect 23204 21836 23256 21888
rect 23296 21836 23348 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 10232 21632 10284 21684
rect 11060 21632 11112 21684
rect 20260 21632 20312 21684
rect 21456 21632 21508 21684
rect 22284 21632 22336 21684
rect 22560 21632 22612 21684
rect 24216 21632 24268 21684
rect 24952 21632 25004 21684
rect 9036 21564 9088 21616
rect 12072 21564 12124 21616
rect 15108 21564 15160 21616
rect 15384 21564 15436 21616
rect 20076 21564 20128 21616
rect 22192 21564 22244 21616
rect 8300 21496 8352 21548
rect 9956 21496 10008 21548
rect 11152 21496 11204 21548
rect 14832 21496 14884 21548
rect 22008 21496 22060 21548
rect 24124 21564 24176 21616
rect 8484 21428 8536 21480
rect 9312 21428 9364 21480
rect 10968 21471 11020 21480
rect 10968 21437 10977 21471
rect 10977 21437 11011 21471
rect 11011 21437 11020 21471
rect 10968 21428 11020 21437
rect 12440 21428 12492 21480
rect 12716 21428 12768 21480
rect 14096 21428 14148 21480
rect 19064 21428 19116 21480
rect 20168 21471 20220 21480
rect 20168 21437 20177 21471
rect 20177 21437 20211 21471
rect 20211 21437 20220 21471
rect 20168 21428 20220 21437
rect 7748 21292 7800 21344
rect 8300 21292 8352 21344
rect 8668 21335 8720 21344
rect 8668 21301 8677 21335
rect 8677 21301 8711 21335
rect 8711 21301 8720 21335
rect 8668 21292 8720 21301
rect 14556 21360 14608 21412
rect 22468 21360 22520 21412
rect 12532 21292 12584 21344
rect 14372 21292 14424 21344
rect 15016 21292 15068 21344
rect 15108 21335 15160 21344
rect 15108 21301 15117 21335
rect 15117 21301 15151 21335
rect 15151 21301 15160 21335
rect 15108 21292 15160 21301
rect 19064 21292 19116 21344
rect 19524 21335 19576 21344
rect 19524 21301 19533 21335
rect 19533 21301 19567 21335
rect 19567 21301 19576 21335
rect 19524 21292 19576 21301
rect 21732 21292 21784 21344
rect 25320 21428 25372 21480
rect 23572 21292 23624 21344
rect 25044 21335 25096 21344
rect 25044 21301 25053 21335
rect 25053 21301 25087 21335
rect 25087 21301 25096 21335
rect 25044 21292 25096 21301
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 4804 21088 4856 21140
rect 19064 21088 19116 21140
rect 20904 21088 20956 21140
rect 22100 21088 22152 21140
rect 25044 21088 25096 21140
rect 13360 21020 13412 21072
rect 16580 21020 16632 21072
rect 9956 20995 10008 21004
rect 9956 20961 9965 20995
rect 9965 20961 9999 20995
rect 9999 20961 10008 20995
rect 9956 20952 10008 20961
rect 19708 20952 19760 21004
rect 22008 20995 22060 21004
rect 22008 20961 22017 20995
rect 22017 20961 22051 20995
rect 22051 20961 22060 20995
rect 22008 20952 22060 20961
rect 9772 20884 9824 20936
rect 18696 20884 18748 20936
rect 19248 20884 19300 20936
rect 3516 20816 3568 20868
rect 10140 20816 10192 20868
rect 10876 20816 10928 20868
rect 12440 20816 12492 20868
rect 14648 20816 14700 20868
rect 15752 20816 15804 20868
rect 8668 20748 8720 20800
rect 9036 20791 9088 20800
rect 9036 20757 9045 20791
rect 9045 20757 9079 20791
rect 9079 20757 9088 20791
rect 9036 20748 9088 20757
rect 15108 20748 15160 20800
rect 20996 20927 21048 20936
rect 20996 20893 21005 20927
rect 21005 20893 21039 20927
rect 21039 20893 21048 20927
rect 20996 20884 21048 20893
rect 24860 20952 24912 21004
rect 24952 20952 25004 21004
rect 23940 20884 23992 20936
rect 16488 20748 16540 20800
rect 17040 20748 17092 20800
rect 17592 20748 17644 20800
rect 19616 20748 19668 20800
rect 24860 20748 24912 20800
rect 24952 20791 25004 20800
rect 24952 20757 24961 20791
rect 24961 20757 24995 20791
rect 24995 20757 25004 20791
rect 24952 20748 25004 20757
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 10416 20587 10468 20596
rect 10416 20553 10425 20587
rect 10425 20553 10459 20587
rect 10459 20553 10468 20587
rect 10416 20544 10468 20553
rect 12624 20544 12676 20596
rect 13636 20544 13688 20596
rect 15568 20544 15620 20596
rect 8300 20476 8352 20528
rect 9312 20476 9364 20528
rect 14648 20408 14700 20460
rect 19432 20544 19484 20596
rect 20812 20587 20864 20596
rect 20812 20553 20821 20587
rect 20821 20553 20855 20587
rect 20855 20553 20864 20587
rect 20812 20544 20864 20553
rect 20904 20587 20956 20596
rect 20904 20553 20913 20587
rect 20913 20553 20947 20587
rect 20947 20553 20956 20587
rect 20904 20544 20956 20553
rect 25320 20587 25372 20596
rect 25320 20553 25329 20587
rect 25329 20553 25363 20587
rect 25363 20553 25372 20587
rect 25320 20544 25372 20553
rect 17132 20519 17184 20528
rect 17132 20485 17141 20519
rect 17141 20485 17175 20519
rect 17175 20485 17184 20519
rect 17132 20476 17184 20485
rect 17592 20476 17644 20528
rect 22744 20476 22796 20528
rect 23388 20476 23440 20528
rect 24124 20476 24176 20528
rect 18420 20408 18472 20460
rect 18696 20408 18748 20460
rect 18788 20408 18840 20460
rect 19156 20408 19208 20460
rect 19800 20408 19852 20460
rect 21824 20408 21876 20460
rect 22192 20451 22244 20460
rect 22192 20417 22201 20451
rect 22201 20417 22235 20451
rect 22235 20417 22244 20451
rect 22192 20408 22244 20417
rect 22468 20408 22520 20460
rect 7748 20383 7800 20392
rect 7748 20349 7757 20383
rect 7757 20349 7791 20383
rect 7791 20349 7800 20383
rect 7748 20340 7800 20349
rect 8484 20340 8536 20392
rect 9496 20340 9548 20392
rect 9956 20340 10008 20392
rect 10232 20340 10284 20392
rect 12716 20383 12768 20392
rect 12716 20349 12725 20383
rect 12725 20349 12759 20383
rect 12759 20349 12768 20383
rect 12716 20340 12768 20349
rect 13452 20340 13504 20392
rect 14372 20340 14424 20392
rect 8484 20204 8536 20256
rect 9312 20204 9364 20256
rect 10416 20204 10468 20256
rect 13544 20204 13596 20256
rect 15108 20272 15160 20324
rect 20996 20340 21048 20392
rect 22284 20340 22336 20392
rect 23572 20383 23624 20392
rect 23572 20349 23581 20383
rect 23581 20349 23615 20383
rect 23615 20349 23624 20383
rect 23572 20340 23624 20349
rect 25136 20340 25188 20392
rect 19156 20272 19208 20324
rect 23480 20272 23532 20324
rect 18696 20204 18748 20256
rect 19064 20247 19116 20256
rect 19064 20213 19073 20247
rect 19073 20213 19107 20247
rect 19107 20213 19116 20247
rect 19064 20204 19116 20213
rect 19800 20204 19852 20256
rect 20536 20204 20588 20256
rect 22744 20247 22796 20256
rect 22744 20213 22753 20247
rect 22753 20213 22787 20247
rect 22787 20213 22796 20247
rect 22744 20204 22796 20213
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 8484 20043 8536 20052
rect 8484 20009 8493 20043
rect 8493 20009 8527 20043
rect 8527 20009 8536 20043
rect 8484 20000 8536 20009
rect 14004 20000 14056 20052
rect 15752 20000 15804 20052
rect 22192 20000 22244 20052
rect 23940 20000 23992 20052
rect 17132 19932 17184 19984
rect 7748 19864 7800 19916
rect 9772 19864 9824 19916
rect 11980 19907 12032 19916
rect 11980 19873 11989 19907
rect 11989 19873 12023 19907
rect 12023 19873 12032 19907
rect 11980 19864 12032 19873
rect 15844 19864 15896 19916
rect 17868 19864 17920 19916
rect 20260 19864 20312 19916
rect 12716 19796 12768 19848
rect 16672 19839 16724 19848
rect 16672 19805 16681 19839
rect 16681 19805 16715 19839
rect 16715 19805 16724 19839
rect 16672 19796 16724 19805
rect 18604 19796 18656 19848
rect 21456 19796 21508 19848
rect 8484 19728 8536 19780
rect 9404 19771 9456 19780
rect 9404 19737 9413 19771
rect 9413 19737 9447 19771
rect 9447 19737 9456 19771
rect 9404 19728 9456 19737
rect 10416 19728 10468 19780
rect 11060 19728 11112 19780
rect 14648 19728 14700 19780
rect 10876 19703 10928 19712
rect 10876 19669 10885 19703
rect 10885 19669 10919 19703
rect 10919 19669 10928 19703
rect 10876 19660 10928 19669
rect 11704 19703 11756 19712
rect 11704 19669 11713 19703
rect 11713 19669 11747 19703
rect 11747 19669 11756 19703
rect 11704 19660 11756 19669
rect 15844 19728 15896 19780
rect 17040 19660 17092 19712
rect 18420 19660 18472 19712
rect 20168 19771 20220 19780
rect 20168 19737 20177 19771
rect 20177 19737 20211 19771
rect 20211 19737 20220 19771
rect 20168 19728 20220 19737
rect 21456 19660 21508 19712
rect 21640 19703 21692 19712
rect 21640 19669 21649 19703
rect 21649 19669 21683 19703
rect 21683 19669 21692 19703
rect 24124 19771 24176 19780
rect 24124 19737 24133 19771
rect 24133 19737 24167 19771
rect 24167 19737 24176 19771
rect 25412 19771 25464 19780
rect 24124 19728 24176 19737
rect 25412 19737 25421 19771
rect 25421 19737 25455 19771
rect 25455 19737 25464 19771
rect 25412 19728 25464 19737
rect 21640 19660 21692 19669
rect 23388 19660 23440 19712
rect 24952 19660 25004 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 8760 19499 8812 19508
rect 8760 19465 8769 19499
rect 8769 19465 8803 19499
rect 8803 19465 8812 19499
rect 8760 19456 8812 19465
rect 11704 19499 11756 19508
rect 11704 19465 11713 19499
rect 11713 19465 11747 19499
rect 11747 19465 11756 19499
rect 11704 19456 11756 19465
rect 11796 19456 11848 19508
rect 8392 19388 8444 19440
rect 9036 19320 9088 19372
rect 10140 19320 10192 19372
rect 10416 19320 10468 19372
rect 17316 19499 17368 19508
rect 17316 19465 17325 19499
rect 17325 19465 17359 19499
rect 17359 19465 17368 19499
rect 17316 19456 17368 19465
rect 19524 19456 19576 19508
rect 20720 19456 20772 19508
rect 24584 19456 24636 19508
rect 25136 19499 25188 19508
rect 25136 19465 25145 19499
rect 25145 19465 25179 19499
rect 25179 19465 25188 19499
rect 25136 19456 25188 19465
rect 25412 19499 25464 19508
rect 25412 19465 25421 19499
rect 25421 19465 25455 19499
rect 25455 19465 25464 19499
rect 25412 19456 25464 19465
rect 6552 19295 6604 19304
rect 6552 19261 6561 19295
rect 6561 19261 6595 19295
rect 6595 19261 6604 19295
rect 6552 19252 6604 19261
rect 6920 19252 6972 19304
rect 9312 19295 9364 19304
rect 9312 19261 9321 19295
rect 9321 19261 9355 19295
rect 9355 19261 9364 19295
rect 9312 19252 9364 19261
rect 10968 19252 11020 19304
rect 12440 19252 12492 19304
rect 8300 19159 8352 19168
rect 8300 19125 8309 19159
rect 8309 19125 8343 19159
rect 8343 19125 8352 19159
rect 8300 19116 8352 19125
rect 9128 19116 9180 19168
rect 13544 19252 13596 19304
rect 16120 19363 16172 19372
rect 16120 19329 16129 19363
rect 16129 19329 16163 19363
rect 16163 19329 16172 19363
rect 16120 19320 16172 19329
rect 16212 19320 16264 19372
rect 22192 19388 22244 19440
rect 15752 19252 15804 19304
rect 19156 19363 19208 19372
rect 19156 19329 19165 19363
rect 19165 19329 19199 19363
rect 19199 19329 19208 19363
rect 19156 19320 19208 19329
rect 19248 19320 19300 19372
rect 23572 19388 23624 19440
rect 23940 19388 23992 19440
rect 24124 19388 24176 19440
rect 19340 19252 19392 19304
rect 14832 19184 14884 19236
rect 21640 19252 21692 19304
rect 22100 19252 22152 19304
rect 21548 19184 21600 19236
rect 21824 19227 21876 19236
rect 21824 19193 21833 19227
rect 21833 19193 21867 19227
rect 21867 19193 21876 19227
rect 21824 19184 21876 19193
rect 21916 19184 21968 19236
rect 12808 19116 12860 19168
rect 14372 19116 14424 19168
rect 14648 19159 14700 19168
rect 14648 19125 14657 19159
rect 14657 19125 14691 19159
rect 14691 19125 14700 19159
rect 14648 19116 14700 19125
rect 15108 19116 15160 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 10048 18955 10100 18964
rect 10048 18921 10057 18955
rect 10057 18921 10091 18955
rect 10091 18921 10100 18955
rect 10048 18912 10100 18921
rect 10784 18912 10836 18964
rect 7932 18844 7984 18896
rect 11060 18844 11112 18896
rect 16672 18844 16724 18896
rect 8300 18776 8352 18828
rect 10600 18819 10652 18828
rect 10600 18785 10609 18819
rect 10609 18785 10643 18819
rect 10643 18785 10652 18819
rect 10600 18776 10652 18785
rect 10876 18776 10928 18828
rect 6644 18751 6696 18760
rect 6644 18717 6653 18751
rect 6653 18717 6687 18751
rect 6687 18717 6696 18751
rect 6644 18708 6696 18717
rect 8668 18708 8720 18760
rect 11704 18708 11756 18760
rect 12164 18708 12216 18760
rect 8300 18640 8352 18692
rect 9496 18640 9548 18692
rect 17500 18819 17552 18828
rect 17500 18785 17509 18819
rect 17509 18785 17543 18819
rect 17543 18785 17552 18819
rect 17500 18776 17552 18785
rect 17316 18708 17368 18760
rect 17776 18708 17828 18760
rect 24400 18844 24452 18896
rect 23848 18819 23900 18828
rect 23848 18785 23857 18819
rect 23857 18785 23891 18819
rect 23891 18785 23900 18819
rect 23848 18776 23900 18785
rect 22192 18751 22244 18760
rect 22192 18717 22201 18751
rect 22201 18717 22235 18751
rect 22235 18717 22244 18751
rect 22192 18708 22244 18717
rect 22744 18751 22796 18760
rect 22744 18717 22753 18751
rect 22753 18717 22787 18751
rect 22787 18717 22796 18751
rect 22744 18708 22796 18717
rect 25596 18912 25648 18964
rect 12348 18640 12400 18692
rect 23388 18640 23440 18692
rect 25228 18640 25280 18692
rect 8484 18572 8536 18624
rect 10876 18572 10928 18624
rect 11060 18572 11112 18624
rect 12624 18572 12676 18624
rect 13452 18572 13504 18624
rect 13820 18615 13872 18624
rect 13820 18581 13829 18615
rect 13829 18581 13863 18615
rect 13863 18581 13872 18615
rect 13820 18572 13872 18581
rect 14280 18615 14332 18624
rect 14280 18581 14289 18615
rect 14289 18581 14323 18615
rect 14323 18581 14332 18615
rect 14280 18572 14332 18581
rect 17040 18572 17092 18624
rect 17132 18572 17184 18624
rect 17592 18572 17644 18624
rect 20536 18572 20588 18624
rect 22100 18572 22152 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 9496 18411 9548 18420
rect 9496 18377 9505 18411
rect 9505 18377 9539 18411
rect 9539 18377 9548 18411
rect 9496 18368 9548 18377
rect 8300 18300 8352 18352
rect 10508 18368 10560 18420
rect 10784 18368 10836 18420
rect 12348 18368 12400 18420
rect 13820 18368 13872 18420
rect 11796 18300 11848 18352
rect 16672 18368 16724 18420
rect 10416 18232 10468 18284
rect 6644 18164 6696 18216
rect 11336 18232 11388 18284
rect 12440 18275 12492 18284
rect 12440 18241 12449 18275
rect 12449 18241 12483 18275
rect 12483 18241 12492 18275
rect 12440 18232 12492 18241
rect 16580 18232 16632 18284
rect 22652 18300 22704 18352
rect 24860 18300 24912 18352
rect 9772 18096 9824 18148
rect 9128 18028 9180 18080
rect 12808 18164 12860 18216
rect 14188 18164 14240 18216
rect 16672 18164 16724 18216
rect 18696 18164 18748 18216
rect 10876 18096 10928 18148
rect 22100 18275 22152 18284
rect 22100 18241 22109 18275
rect 22109 18241 22143 18275
rect 22143 18241 22152 18275
rect 22100 18232 22152 18241
rect 23480 18232 23532 18284
rect 24676 18207 24728 18216
rect 24676 18173 24685 18207
rect 24685 18173 24719 18207
rect 24719 18173 24728 18207
rect 24676 18164 24728 18173
rect 20812 18096 20864 18148
rect 11060 18071 11112 18080
rect 11060 18037 11069 18071
rect 11069 18037 11103 18071
rect 11103 18037 11112 18071
rect 11060 18028 11112 18037
rect 18328 18028 18380 18080
rect 21088 18071 21140 18080
rect 21088 18037 21097 18071
rect 21097 18037 21131 18071
rect 21131 18037 21140 18071
rect 21088 18028 21140 18037
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 7656 17824 7708 17876
rect 15200 17824 15252 17876
rect 20720 17824 20772 17876
rect 24032 17824 24084 17876
rect 7840 17688 7892 17740
rect 11704 17688 11756 17740
rect 11980 17688 12032 17740
rect 13820 17756 13872 17808
rect 13360 17688 13412 17740
rect 16304 17756 16356 17808
rect 17224 17756 17276 17808
rect 17868 17756 17920 17808
rect 18328 17756 18380 17808
rect 17592 17688 17644 17740
rect 18880 17688 18932 17740
rect 21548 17756 21600 17808
rect 9772 17663 9824 17672
rect 9772 17629 9781 17663
rect 9781 17629 9815 17663
rect 9815 17629 9824 17663
rect 9772 17620 9824 17629
rect 14280 17620 14332 17672
rect 15752 17620 15804 17672
rect 16948 17620 17000 17672
rect 19340 17620 19392 17672
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 25688 17756 25740 17808
rect 24860 17688 24912 17740
rect 24952 17688 25004 17740
rect 25136 17731 25188 17740
rect 25136 17697 25145 17731
rect 25145 17697 25179 17731
rect 25179 17697 25188 17731
rect 25136 17688 25188 17697
rect 22836 17663 22888 17672
rect 22836 17629 22845 17663
rect 22845 17629 22879 17663
rect 22879 17629 22888 17663
rect 22836 17620 22888 17629
rect 8852 17552 8904 17604
rect 9956 17552 10008 17604
rect 11060 17552 11112 17604
rect 13728 17552 13780 17604
rect 16856 17552 16908 17604
rect 17684 17552 17736 17604
rect 17776 17595 17828 17604
rect 17776 17561 17785 17595
rect 17785 17561 17819 17595
rect 17819 17561 17828 17595
rect 17776 17552 17828 17561
rect 7196 17527 7248 17536
rect 7196 17493 7205 17527
rect 7205 17493 7239 17527
rect 7239 17493 7248 17527
rect 7196 17484 7248 17493
rect 7656 17484 7708 17536
rect 9404 17484 9456 17536
rect 13176 17484 13228 17536
rect 15476 17527 15528 17536
rect 15476 17493 15485 17527
rect 15485 17493 15519 17527
rect 15519 17493 15528 17527
rect 15476 17484 15528 17493
rect 17408 17527 17460 17536
rect 17408 17493 17417 17527
rect 17417 17493 17451 17527
rect 17451 17493 17460 17527
rect 17408 17484 17460 17493
rect 17868 17527 17920 17536
rect 17868 17493 17877 17527
rect 17877 17493 17911 17527
rect 17911 17493 17920 17527
rect 18696 17527 18748 17536
rect 17868 17484 17920 17493
rect 18696 17493 18705 17527
rect 18705 17493 18739 17527
rect 18739 17493 18748 17527
rect 18696 17484 18748 17493
rect 19892 17484 19944 17536
rect 22008 17595 22060 17604
rect 22008 17561 22017 17595
rect 22017 17561 22051 17595
rect 22051 17561 22060 17595
rect 22008 17552 22060 17561
rect 22192 17595 22244 17604
rect 22192 17561 22201 17595
rect 22201 17561 22235 17595
rect 22235 17561 22244 17595
rect 22192 17552 22244 17561
rect 21088 17484 21140 17536
rect 25044 17552 25096 17604
rect 23756 17484 23808 17536
rect 24676 17484 24728 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 7196 17280 7248 17332
rect 9220 17280 9272 17332
rect 9404 17323 9456 17332
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 11520 17280 11572 17332
rect 12440 17280 12492 17332
rect 13728 17280 13780 17332
rect 9772 17212 9824 17264
rect 13176 17255 13228 17264
rect 13176 17221 13185 17255
rect 13185 17221 13219 17255
rect 13219 17221 13228 17255
rect 13176 17212 13228 17221
rect 16396 17280 16448 17332
rect 16580 17280 16632 17332
rect 17592 17280 17644 17332
rect 20168 17280 20220 17332
rect 22008 17323 22060 17332
rect 22008 17289 22017 17323
rect 22017 17289 22051 17323
rect 22051 17289 22060 17323
rect 22008 17280 22060 17289
rect 24492 17280 24544 17332
rect 11520 17144 11572 17196
rect 16948 17255 17000 17264
rect 16948 17221 16957 17255
rect 16957 17221 16991 17255
rect 16991 17221 17000 17255
rect 16948 17212 17000 17221
rect 18972 17212 19024 17264
rect 20812 17212 20864 17264
rect 21824 17212 21876 17264
rect 23664 17212 23716 17264
rect 23480 17187 23532 17196
rect 23480 17153 23489 17187
rect 23489 17153 23523 17187
rect 23523 17153 23532 17187
rect 23480 17144 23532 17153
rect 24860 17144 24912 17196
rect 7564 17008 7616 17060
rect 3332 16940 3384 16992
rect 8576 17076 8628 17128
rect 9404 17076 9456 17128
rect 9588 17119 9640 17128
rect 9588 17085 9597 17119
rect 9597 17085 9631 17119
rect 9631 17085 9640 17119
rect 9588 17076 9640 17085
rect 11060 17076 11112 17128
rect 11520 16983 11572 16992
rect 11520 16949 11529 16983
rect 11529 16949 11563 16983
rect 11563 16949 11572 16983
rect 11520 16940 11572 16949
rect 11980 16940 12032 16992
rect 12716 17076 12768 17128
rect 13544 17076 13596 17128
rect 15568 17076 15620 17128
rect 16120 17076 16172 17128
rect 16948 17076 17000 17128
rect 17868 17076 17920 17128
rect 18880 17119 18932 17128
rect 18880 17085 18889 17119
rect 18889 17085 18923 17119
rect 18923 17085 18932 17119
rect 18880 17076 18932 17085
rect 22560 17076 22612 17128
rect 13636 17008 13688 17060
rect 15936 17008 15988 17060
rect 16028 17008 16080 17060
rect 20904 17008 20956 17060
rect 13820 16940 13872 16992
rect 16672 16940 16724 16992
rect 18696 16940 18748 16992
rect 18972 16940 19024 16992
rect 20352 16940 20404 16992
rect 22100 16940 22152 16992
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 8576 16779 8628 16788
rect 8576 16745 8585 16779
rect 8585 16745 8619 16779
rect 8619 16745 8628 16779
rect 8576 16736 8628 16745
rect 11336 16779 11388 16788
rect 11336 16745 11345 16779
rect 11345 16745 11379 16779
rect 11379 16745 11388 16779
rect 11336 16736 11388 16745
rect 11888 16736 11940 16788
rect 11612 16668 11664 16720
rect 11336 16600 11388 16652
rect 12808 16600 12860 16652
rect 13820 16668 13872 16720
rect 14648 16736 14700 16788
rect 13544 16600 13596 16652
rect 16488 16668 16540 16720
rect 21824 16736 21876 16788
rect 16948 16668 17000 16720
rect 17776 16668 17828 16720
rect 19800 16668 19852 16720
rect 13636 16532 13688 16584
rect 10324 16464 10376 16516
rect 9864 16439 9916 16448
rect 9864 16405 9873 16439
rect 9873 16405 9907 16439
rect 9907 16405 9916 16439
rect 9864 16396 9916 16405
rect 10232 16439 10284 16448
rect 10232 16405 10241 16439
rect 10241 16405 10275 16439
rect 10275 16405 10284 16439
rect 10232 16396 10284 16405
rect 14372 16464 14424 16516
rect 13544 16439 13596 16448
rect 13544 16405 13553 16439
rect 13553 16405 13587 16439
rect 13587 16405 13596 16439
rect 13544 16396 13596 16405
rect 14280 16439 14332 16448
rect 14280 16405 14289 16439
rect 14289 16405 14323 16439
rect 14323 16405 14332 16439
rect 14280 16396 14332 16405
rect 15476 16532 15528 16584
rect 16396 16600 16448 16652
rect 17868 16600 17920 16652
rect 20260 16643 20312 16652
rect 20260 16609 20269 16643
rect 20269 16609 20303 16643
rect 20303 16609 20312 16643
rect 20260 16600 20312 16609
rect 15660 16464 15712 16516
rect 16856 16464 16908 16516
rect 15016 16439 15068 16448
rect 15016 16405 15025 16439
rect 15025 16405 15059 16439
rect 15059 16405 15068 16439
rect 15016 16396 15068 16405
rect 15844 16396 15896 16448
rect 16212 16439 16264 16448
rect 16212 16405 16221 16439
rect 16221 16405 16255 16439
rect 16255 16405 16264 16439
rect 16212 16396 16264 16405
rect 18696 16439 18748 16448
rect 18696 16405 18705 16439
rect 18705 16405 18739 16439
rect 18739 16405 18748 16439
rect 18696 16396 18748 16405
rect 19432 16396 19484 16448
rect 19524 16396 19576 16448
rect 20444 16464 20496 16516
rect 21824 16464 21876 16516
rect 22376 16532 22428 16584
rect 22652 16575 22704 16584
rect 22652 16541 22661 16575
rect 22661 16541 22695 16575
rect 22695 16541 22704 16575
rect 22652 16532 22704 16541
rect 23388 16532 23440 16584
rect 24768 16575 24820 16584
rect 24768 16541 24777 16575
rect 24777 16541 24811 16575
rect 24811 16541 24820 16575
rect 24768 16532 24820 16541
rect 22284 16464 22336 16516
rect 23848 16464 23900 16516
rect 24216 16464 24268 16516
rect 24860 16464 24912 16516
rect 22100 16396 22152 16448
rect 22376 16396 22428 16448
rect 22836 16396 22888 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 8300 16235 8352 16244
rect 8300 16201 8309 16235
rect 8309 16201 8343 16235
rect 8343 16201 8352 16235
rect 8300 16192 8352 16201
rect 9312 16192 9364 16244
rect 11612 16192 11664 16244
rect 15016 16192 15068 16244
rect 15660 16192 15712 16244
rect 16212 16235 16264 16244
rect 16212 16201 16221 16235
rect 16221 16201 16255 16235
rect 16255 16201 16264 16235
rect 16212 16192 16264 16201
rect 16856 16235 16908 16244
rect 16856 16201 16865 16235
rect 16865 16201 16899 16235
rect 16899 16201 16908 16235
rect 16856 16192 16908 16201
rect 18696 16192 18748 16244
rect 24768 16192 24820 16244
rect 8392 16124 8444 16176
rect 8668 16124 8720 16176
rect 11704 16124 11756 16176
rect 6552 16099 6604 16108
rect 6552 16065 6561 16099
rect 6561 16065 6595 16099
rect 6595 16065 6604 16099
rect 6552 16056 6604 16065
rect 8392 15988 8444 16040
rect 9588 15988 9640 16040
rect 12716 16124 12768 16176
rect 14372 16124 14424 16176
rect 12440 16056 12492 16108
rect 12256 15988 12308 16040
rect 12072 15920 12124 15972
rect 5172 15852 5224 15904
rect 11980 15852 12032 15904
rect 14280 16056 14332 16108
rect 14740 16056 14792 16108
rect 14372 15988 14424 16040
rect 15016 16031 15068 16040
rect 15016 15997 15025 16031
rect 15025 15997 15059 16031
rect 15059 15997 15068 16031
rect 15016 15988 15068 15997
rect 17224 16167 17276 16176
rect 17224 16133 17233 16167
rect 17233 16133 17267 16167
rect 17267 16133 17276 16167
rect 17224 16124 17276 16133
rect 19340 16124 19392 16176
rect 20260 16124 20312 16176
rect 19432 16056 19484 16108
rect 19800 16056 19852 16108
rect 21824 16124 21876 16176
rect 18788 15988 18840 16040
rect 21180 16031 21232 16040
rect 21180 15997 21189 16031
rect 21189 15997 21223 16031
rect 21223 15997 21232 16031
rect 21180 15988 21232 15997
rect 21364 16031 21416 16040
rect 21364 15997 21373 16031
rect 21373 15997 21407 16031
rect 21407 15997 21416 16031
rect 21364 15988 21416 15997
rect 14280 15920 14332 15972
rect 18696 15920 18748 15972
rect 19156 15920 19208 15972
rect 20812 15920 20864 15972
rect 14004 15852 14056 15904
rect 17316 15895 17368 15904
rect 17316 15861 17325 15895
rect 17325 15861 17359 15895
rect 17359 15861 17368 15895
rect 17316 15852 17368 15861
rect 17684 15852 17736 15904
rect 18604 15852 18656 15904
rect 21456 15852 21508 15904
rect 23572 16056 23624 16108
rect 22376 15988 22428 16040
rect 24584 15988 24636 16040
rect 22284 15852 22336 15904
rect 23388 15852 23440 15904
rect 23756 15895 23808 15904
rect 23756 15861 23765 15895
rect 23765 15861 23799 15895
rect 23799 15861 23808 15895
rect 23756 15852 23808 15861
rect 24216 15852 24268 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 9036 15648 9088 15700
rect 11152 15648 11204 15700
rect 15016 15648 15068 15700
rect 17132 15648 17184 15700
rect 18236 15648 18288 15700
rect 5448 15580 5500 15632
rect 12716 15580 12768 15632
rect 9588 15512 9640 15564
rect 12256 15555 12308 15564
rect 12256 15521 12265 15555
rect 12265 15521 12299 15555
rect 12299 15521 12308 15555
rect 12256 15512 12308 15521
rect 16396 15555 16448 15564
rect 16396 15521 16405 15555
rect 16405 15521 16439 15555
rect 16439 15521 16448 15555
rect 16396 15512 16448 15521
rect 18328 15512 18380 15564
rect 8668 15444 8720 15496
rect 13360 15444 13412 15496
rect 19156 15648 19208 15700
rect 20444 15648 20496 15700
rect 23020 15648 23072 15700
rect 21364 15580 21416 15632
rect 20260 15512 20312 15564
rect 22284 15555 22336 15564
rect 22284 15521 22293 15555
rect 22293 15521 22327 15555
rect 22327 15521 22336 15555
rect 22284 15512 22336 15521
rect 23756 15512 23808 15564
rect 20812 15444 20864 15496
rect 9220 15376 9272 15428
rect 12532 15376 12584 15428
rect 16396 15376 16448 15428
rect 16948 15376 17000 15428
rect 19708 15419 19760 15428
rect 19708 15385 19717 15419
rect 19717 15385 19751 15419
rect 19751 15385 19760 15419
rect 19708 15376 19760 15385
rect 21088 15444 21140 15496
rect 21364 15376 21416 15428
rect 23020 15376 23072 15428
rect 23940 15512 23992 15564
rect 24676 15512 24728 15564
rect 10048 15308 10100 15360
rect 12440 15308 12492 15360
rect 14188 15308 14240 15360
rect 14280 15351 14332 15360
rect 14280 15317 14289 15351
rect 14289 15317 14323 15351
rect 14323 15317 14332 15351
rect 14280 15308 14332 15317
rect 14740 15351 14792 15360
rect 14740 15317 14749 15351
rect 14749 15317 14783 15351
rect 14783 15317 14792 15351
rect 14740 15308 14792 15317
rect 15752 15351 15804 15360
rect 15752 15317 15761 15351
rect 15761 15317 15795 15351
rect 15795 15317 15804 15351
rect 15752 15308 15804 15317
rect 16764 15308 16816 15360
rect 17500 15308 17552 15360
rect 19524 15308 19576 15360
rect 20352 15308 20404 15360
rect 23940 15308 23992 15360
rect 24216 15308 24268 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 10140 15147 10192 15156
rect 10140 15113 10149 15147
rect 10149 15113 10183 15147
rect 10183 15113 10192 15147
rect 10140 15104 10192 15113
rect 8668 15036 8720 15088
rect 11428 15036 11480 15088
rect 14280 15104 14332 15156
rect 15752 15104 15804 15156
rect 17224 15104 17276 15156
rect 19616 15104 19668 15156
rect 21088 15104 21140 15156
rect 21916 15104 21968 15156
rect 16120 15036 16172 15088
rect 19248 15036 19300 15088
rect 9588 14968 9640 15020
rect 8300 14900 8352 14952
rect 9036 14832 9088 14884
rect 11244 14900 11296 14952
rect 15936 14968 15988 15020
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 23204 15036 23256 15088
rect 23296 15079 23348 15088
rect 23296 15045 23305 15079
rect 23305 15045 23339 15079
rect 23339 15045 23348 15079
rect 23296 15036 23348 15045
rect 25136 15079 25188 15088
rect 25136 15045 25145 15079
rect 25145 15045 25179 15079
rect 25179 15045 25188 15079
rect 25136 15036 25188 15045
rect 21364 15011 21416 15020
rect 21364 14977 21373 15011
rect 21373 14977 21407 15011
rect 21407 14977 21416 15011
rect 21364 14968 21416 14977
rect 22008 14968 22060 15020
rect 24124 15011 24176 15020
rect 24124 14977 24133 15011
rect 24133 14977 24167 15011
rect 24167 14977 24176 15011
rect 24124 14968 24176 14977
rect 11612 14832 11664 14884
rect 11980 14832 12032 14884
rect 13636 14832 13688 14884
rect 16580 14900 16632 14952
rect 19892 14900 19944 14952
rect 20444 14900 20496 14952
rect 22744 14900 22796 14952
rect 8300 14764 8352 14816
rect 11520 14764 11572 14816
rect 12348 14764 12400 14816
rect 12808 14764 12860 14816
rect 15476 14764 15528 14816
rect 15844 14764 15896 14816
rect 22284 14764 22336 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 7840 14560 7892 14612
rect 8668 14560 8720 14612
rect 9036 14560 9088 14612
rect 6460 14467 6512 14476
rect 6460 14433 6469 14467
rect 6469 14433 6503 14467
rect 6503 14433 6512 14467
rect 6460 14424 6512 14433
rect 8300 14424 8352 14476
rect 9312 14288 9364 14340
rect 12624 14560 12676 14612
rect 14648 14560 14700 14612
rect 20168 14560 20220 14612
rect 24032 14560 24084 14612
rect 10232 14467 10284 14476
rect 10232 14433 10241 14467
rect 10241 14433 10275 14467
rect 10275 14433 10284 14467
rect 10232 14424 10284 14433
rect 11888 14424 11940 14476
rect 12256 14424 12308 14476
rect 16856 14492 16908 14544
rect 15384 14424 15436 14476
rect 19524 14492 19576 14544
rect 22468 14492 22520 14544
rect 17132 14467 17184 14476
rect 17132 14433 17141 14467
rect 17141 14433 17175 14467
rect 17175 14433 17184 14467
rect 17132 14424 17184 14433
rect 20628 14424 20680 14476
rect 23296 14424 23348 14476
rect 24860 14424 24912 14476
rect 9588 14356 9640 14408
rect 13084 14356 13136 14408
rect 13636 14288 13688 14340
rect 14740 14331 14792 14340
rect 14740 14297 14749 14331
rect 14749 14297 14783 14331
rect 14783 14297 14792 14331
rect 14740 14288 14792 14297
rect 16120 14356 16172 14408
rect 19616 14356 19668 14408
rect 21640 14356 21692 14408
rect 24492 14356 24544 14408
rect 25044 14399 25096 14408
rect 25044 14365 25053 14399
rect 25053 14365 25087 14399
rect 25087 14365 25096 14399
rect 25044 14356 25096 14365
rect 12716 14220 12768 14272
rect 13912 14263 13964 14272
rect 13912 14229 13921 14263
rect 13921 14229 13955 14263
rect 13955 14229 13964 14263
rect 13912 14220 13964 14229
rect 14280 14263 14332 14272
rect 14280 14229 14289 14263
rect 14289 14229 14323 14263
rect 14323 14229 14332 14263
rect 14280 14220 14332 14229
rect 14648 14263 14700 14272
rect 14648 14229 14657 14263
rect 14657 14229 14691 14263
rect 14691 14229 14700 14263
rect 14648 14220 14700 14229
rect 16488 14263 16540 14272
rect 16488 14229 16497 14263
rect 16497 14229 16531 14263
rect 16531 14229 16540 14263
rect 16488 14220 16540 14229
rect 21272 14288 21324 14340
rect 19340 14220 19392 14272
rect 19892 14220 19944 14272
rect 21824 14263 21876 14272
rect 21824 14229 21833 14263
rect 21833 14229 21867 14263
rect 21867 14229 21876 14263
rect 21824 14220 21876 14229
rect 24860 14263 24912 14272
rect 24860 14229 24869 14263
rect 24869 14229 24903 14263
rect 24903 14229 24912 14263
rect 24860 14220 24912 14229
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 8300 14016 8352 14068
rect 9588 14016 9640 14068
rect 12256 14059 12308 14068
rect 12256 14025 12265 14059
rect 12265 14025 12299 14059
rect 12299 14025 12308 14059
rect 12256 14016 12308 14025
rect 13084 14016 13136 14068
rect 15568 14059 15620 14068
rect 15568 14025 15577 14059
rect 15577 14025 15611 14059
rect 15611 14025 15620 14059
rect 15568 14016 15620 14025
rect 16488 14016 16540 14068
rect 7932 13948 7984 14000
rect 8668 13948 8720 14000
rect 12348 13948 12400 14000
rect 17132 13948 17184 14000
rect 19156 13991 19208 14000
rect 19156 13957 19165 13991
rect 19165 13957 19199 13991
rect 19199 13957 19208 13991
rect 19156 13948 19208 13957
rect 19524 13991 19576 14000
rect 19524 13957 19533 13991
rect 19533 13957 19567 13991
rect 19567 13957 19576 13991
rect 19524 13948 19576 13957
rect 19616 13948 19668 14000
rect 9588 13880 9640 13932
rect 10232 13812 10284 13864
rect 11060 13812 11112 13864
rect 12256 13812 12308 13864
rect 12808 13744 12860 13796
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 13820 13812 13872 13821
rect 16488 13812 16540 13864
rect 16856 13855 16908 13864
rect 16856 13821 16865 13855
rect 16865 13821 16899 13855
rect 16899 13821 16908 13855
rect 16856 13812 16908 13821
rect 17592 13812 17644 13864
rect 17868 13812 17920 13864
rect 21088 13923 21140 13932
rect 21088 13889 21097 13923
rect 21097 13889 21131 13923
rect 21131 13889 21140 13923
rect 21088 13880 21140 13889
rect 18880 13812 18932 13864
rect 23388 14016 23440 14068
rect 21548 13948 21600 14000
rect 21272 13880 21324 13932
rect 24216 13880 24268 13932
rect 15568 13744 15620 13796
rect 22652 13812 22704 13864
rect 22836 13855 22888 13864
rect 22836 13821 22845 13855
rect 22845 13821 22879 13855
rect 22879 13821 22888 13855
rect 22836 13812 22888 13821
rect 12624 13719 12676 13728
rect 12624 13685 12633 13719
rect 12633 13685 12667 13719
rect 12667 13685 12676 13719
rect 12624 13676 12676 13685
rect 14096 13719 14148 13728
rect 14096 13685 14126 13719
rect 14126 13685 14148 13719
rect 14096 13676 14148 13685
rect 18328 13676 18380 13728
rect 20628 13676 20680 13728
rect 20904 13719 20956 13728
rect 20904 13685 20913 13719
rect 20913 13685 20947 13719
rect 20947 13685 20956 13719
rect 20904 13676 20956 13685
rect 20996 13676 21048 13728
rect 23204 13812 23256 13864
rect 23848 13676 23900 13728
rect 25044 13719 25096 13728
rect 25044 13685 25053 13719
rect 25053 13685 25087 13719
rect 25087 13685 25096 13719
rect 25044 13676 25096 13685
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 8392 13472 8444 13524
rect 8668 13515 8720 13524
rect 8668 13481 8677 13515
rect 8677 13481 8711 13515
rect 8711 13481 8720 13515
rect 8668 13472 8720 13481
rect 8852 13472 8904 13524
rect 13544 13472 13596 13524
rect 14740 13472 14792 13524
rect 21088 13515 21140 13524
rect 21088 13481 21097 13515
rect 21097 13481 21131 13515
rect 21131 13481 21140 13515
rect 21088 13472 21140 13481
rect 24492 13472 24544 13524
rect 9312 13404 9364 13456
rect 6460 13336 6512 13388
rect 9680 13336 9732 13388
rect 11796 13404 11848 13456
rect 14556 13404 14608 13456
rect 17132 13404 17184 13456
rect 24216 13404 24268 13456
rect 11704 13336 11756 13388
rect 13820 13336 13872 13388
rect 15384 13336 15436 13388
rect 15752 13379 15804 13388
rect 15752 13345 15761 13379
rect 15761 13345 15795 13379
rect 15795 13345 15804 13379
rect 15752 13336 15804 13345
rect 12440 13268 12492 13320
rect 8668 13200 8720 13252
rect 9680 13175 9732 13184
rect 9680 13141 9689 13175
rect 9689 13141 9723 13175
rect 9723 13141 9732 13175
rect 9680 13132 9732 13141
rect 11980 13200 12032 13252
rect 12072 13132 12124 13184
rect 12164 13175 12216 13184
rect 12164 13141 12173 13175
rect 12173 13141 12207 13175
rect 12207 13141 12216 13175
rect 12164 13132 12216 13141
rect 12992 13268 13044 13320
rect 13360 13268 13412 13320
rect 14372 13268 14424 13320
rect 14556 13268 14608 13320
rect 14924 13311 14976 13320
rect 14924 13277 14933 13311
rect 14933 13277 14967 13311
rect 14967 13277 14976 13311
rect 14924 13268 14976 13277
rect 16212 13268 16264 13320
rect 20076 13336 20128 13388
rect 20444 13336 20496 13388
rect 22836 13336 22888 13388
rect 23756 13379 23808 13388
rect 23756 13345 23765 13379
rect 23765 13345 23799 13379
rect 23799 13345 23808 13379
rect 23756 13336 23808 13345
rect 17500 13311 17552 13320
rect 17500 13277 17509 13311
rect 17509 13277 17543 13311
rect 17543 13277 17552 13311
rect 17500 13268 17552 13277
rect 18696 13268 18748 13320
rect 18328 13200 18380 13252
rect 18420 13200 18472 13252
rect 19432 13311 19484 13320
rect 19432 13277 19441 13311
rect 19441 13277 19475 13311
rect 19475 13277 19484 13311
rect 19432 13268 19484 13277
rect 20720 13243 20772 13252
rect 20720 13209 20729 13243
rect 20729 13209 20763 13243
rect 20763 13209 20772 13243
rect 20720 13200 20772 13209
rect 13912 13175 13964 13184
rect 13912 13141 13921 13175
rect 13921 13141 13955 13175
rect 13955 13141 13964 13175
rect 13912 13132 13964 13141
rect 14648 13175 14700 13184
rect 14648 13141 14657 13175
rect 14657 13141 14691 13175
rect 14691 13141 14700 13175
rect 14648 13132 14700 13141
rect 15292 13132 15344 13184
rect 15384 13132 15436 13184
rect 15844 13132 15896 13184
rect 21548 13268 21600 13320
rect 25044 13336 25096 13388
rect 23388 13200 23440 13252
rect 21640 13132 21692 13184
rect 24308 13132 24360 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 7748 12928 7800 12980
rect 9220 12928 9272 12980
rect 9404 12971 9456 12980
rect 9404 12937 9413 12971
rect 9413 12937 9447 12971
rect 9447 12937 9456 12971
rect 9404 12928 9456 12937
rect 10048 12928 10100 12980
rect 11060 12928 11112 12980
rect 11796 12928 11848 12980
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 11980 12928 12032 12980
rect 12256 12971 12308 12980
rect 12256 12937 12265 12971
rect 12265 12937 12299 12971
rect 12299 12937 12308 12971
rect 12256 12928 12308 12937
rect 12440 12928 12492 12980
rect 12624 12860 12676 12912
rect 13084 12903 13136 12912
rect 13084 12869 13093 12903
rect 13093 12869 13127 12903
rect 13127 12869 13136 12903
rect 13084 12860 13136 12869
rect 13452 12860 13504 12912
rect 14372 12928 14424 12980
rect 16948 12928 17000 12980
rect 17408 12928 17460 12980
rect 19432 12928 19484 12980
rect 21272 12928 21324 12980
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 7288 12792 7340 12844
rect 8208 12835 8260 12844
rect 8208 12801 8217 12835
rect 8217 12801 8251 12835
rect 8251 12801 8260 12835
rect 8208 12792 8260 12801
rect 11796 12792 11848 12844
rect 6920 12724 6972 12776
rect 7840 12724 7892 12776
rect 8484 12767 8536 12776
rect 8484 12733 8493 12767
rect 8493 12733 8527 12767
rect 8527 12733 8536 12767
rect 8484 12724 8536 12733
rect 9772 12724 9824 12776
rect 9956 12724 10008 12776
rect 10968 12767 11020 12776
rect 10968 12733 10977 12767
rect 10977 12733 11011 12767
rect 11011 12733 11020 12767
rect 10968 12724 11020 12733
rect 12808 12792 12860 12844
rect 10416 12656 10468 12708
rect 8852 12588 8904 12640
rect 11888 12656 11940 12708
rect 12992 12588 13044 12640
rect 15108 12792 15160 12844
rect 13820 12724 13872 12776
rect 14096 12724 14148 12776
rect 13544 12588 13596 12640
rect 14372 12588 14424 12640
rect 15016 12631 15068 12640
rect 15016 12597 15025 12631
rect 15025 12597 15059 12631
rect 15059 12597 15068 12631
rect 15016 12588 15068 12597
rect 15476 12835 15528 12844
rect 15476 12801 15485 12835
rect 15485 12801 15519 12835
rect 15519 12801 15528 12835
rect 15476 12792 15528 12801
rect 17224 12835 17276 12844
rect 17224 12801 17233 12835
rect 17233 12801 17267 12835
rect 17267 12801 17276 12835
rect 17224 12792 17276 12801
rect 20628 12860 20680 12912
rect 23296 12860 23348 12912
rect 24308 12928 24360 12980
rect 18788 12792 18840 12844
rect 20812 12792 20864 12844
rect 21088 12835 21140 12844
rect 21088 12801 21097 12835
rect 21097 12801 21131 12835
rect 21131 12801 21140 12835
rect 21088 12792 21140 12801
rect 15568 12767 15620 12776
rect 15568 12733 15577 12767
rect 15577 12733 15611 12767
rect 15611 12733 15620 12767
rect 15568 12724 15620 12733
rect 15844 12724 15896 12776
rect 18880 12724 18932 12776
rect 19248 12767 19300 12776
rect 19248 12733 19257 12767
rect 19257 12733 19291 12767
rect 19291 12733 19300 12767
rect 19248 12724 19300 12733
rect 22100 12792 22152 12844
rect 22192 12835 22244 12844
rect 22192 12801 22201 12835
rect 22201 12801 22235 12835
rect 22235 12801 22244 12835
rect 22192 12792 22244 12801
rect 22468 12792 22520 12844
rect 22836 12792 22888 12844
rect 17132 12656 17184 12708
rect 21180 12656 21232 12708
rect 22008 12699 22060 12708
rect 22008 12665 22017 12699
rect 22017 12665 22051 12699
rect 22051 12665 22060 12699
rect 22008 12656 22060 12665
rect 22560 12656 22612 12708
rect 19432 12588 19484 12640
rect 21916 12588 21968 12640
rect 22100 12588 22152 12640
rect 22468 12588 22520 12640
rect 22836 12588 22888 12640
rect 23388 12588 23440 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 7564 12384 7616 12436
rect 11428 12427 11480 12436
rect 11428 12393 11437 12427
rect 11437 12393 11471 12427
rect 11471 12393 11480 12427
rect 11428 12384 11480 12393
rect 12532 12384 12584 12436
rect 13912 12384 13964 12436
rect 17316 12384 17368 12436
rect 18512 12384 18564 12436
rect 18880 12384 18932 12436
rect 21732 12384 21784 12436
rect 24124 12384 24176 12436
rect 12440 12316 12492 12368
rect 14096 12316 14148 12368
rect 14188 12316 14240 12368
rect 15200 12316 15252 12368
rect 18604 12316 18656 12368
rect 18972 12316 19024 12368
rect 22468 12316 22520 12368
rect 22836 12316 22888 12368
rect 7012 12248 7064 12300
rect 8208 12291 8260 12300
rect 8208 12257 8217 12291
rect 8217 12257 8251 12291
rect 8251 12257 8260 12291
rect 8208 12248 8260 12257
rect 9312 12248 9364 12300
rect 11060 12248 11112 12300
rect 11980 12291 12032 12300
rect 11980 12257 11989 12291
rect 11989 12257 12023 12291
rect 12023 12257 12032 12291
rect 11980 12248 12032 12257
rect 12532 12112 12584 12164
rect 13728 12248 13780 12300
rect 15844 12248 15896 12300
rect 16856 12248 16908 12300
rect 12808 12180 12860 12232
rect 13452 12180 13504 12232
rect 14648 12180 14700 12232
rect 17316 12223 17368 12232
rect 17316 12189 17325 12223
rect 17325 12189 17359 12223
rect 17359 12189 17368 12223
rect 17316 12180 17368 12189
rect 18788 12248 18840 12300
rect 20444 12291 20496 12300
rect 20444 12257 20453 12291
rect 20453 12257 20487 12291
rect 20487 12257 20496 12291
rect 20444 12248 20496 12257
rect 21272 12248 21324 12300
rect 19248 12180 19300 12232
rect 20168 12180 20220 12232
rect 8484 12044 8536 12096
rect 9404 12044 9456 12096
rect 10600 12087 10652 12096
rect 10600 12053 10609 12087
rect 10609 12053 10643 12087
rect 10643 12053 10652 12087
rect 10600 12044 10652 12053
rect 12440 12044 12492 12096
rect 13268 12044 13320 12096
rect 15016 12112 15068 12164
rect 16948 12112 17000 12164
rect 19708 12112 19760 12164
rect 15568 12044 15620 12096
rect 16028 12044 16080 12096
rect 18420 12044 18472 12096
rect 18972 12044 19024 12096
rect 22008 12112 22060 12164
rect 24492 12180 24544 12232
rect 23572 12112 23624 12164
rect 24952 12112 25004 12164
rect 21732 12044 21784 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 3700 11840 3752 11892
rect 9312 11840 9364 11892
rect 9680 11840 9732 11892
rect 10876 11840 10928 11892
rect 12716 11840 12768 11892
rect 13360 11840 13412 11892
rect 13452 11883 13504 11892
rect 13452 11849 13461 11883
rect 13461 11849 13495 11883
rect 13495 11849 13504 11883
rect 13452 11840 13504 11849
rect 13912 11840 13964 11892
rect 14004 11840 14056 11892
rect 14832 11840 14884 11892
rect 15200 11840 15252 11892
rect 16764 11840 16816 11892
rect 17040 11840 17092 11892
rect 14188 11772 14240 11824
rect 15016 11772 15068 11824
rect 18420 11883 18472 11892
rect 18420 11849 18429 11883
rect 18429 11849 18463 11883
rect 18463 11849 18472 11883
rect 18420 11840 18472 11849
rect 19524 11840 19576 11892
rect 8668 11704 8720 11756
rect 9404 11704 9456 11756
rect 9496 11704 9548 11756
rect 11244 11747 11296 11756
rect 11244 11713 11253 11747
rect 11253 11713 11287 11747
rect 11287 11713 11296 11747
rect 11244 11704 11296 11713
rect 14004 11704 14056 11756
rect 15108 11704 15160 11756
rect 15384 11747 15436 11756
rect 15384 11713 15393 11747
rect 15393 11713 15427 11747
rect 15427 11713 15436 11747
rect 15384 11704 15436 11713
rect 15660 11704 15712 11756
rect 16120 11704 16172 11756
rect 16580 11704 16632 11756
rect 19984 11772 20036 11824
rect 20168 11840 20220 11892
rect 24400 11840 24452 11892
rect 24860 11772 24912 11824
rect 19524 11704 19576 11756
rect 20076 11747 20128 11756
rect 20076 11713 20085 11747
rect 20085 11713 20119 11747
rect 20119 11713 20128 11747
rect 20076 11704 20128 11713
rect 12440 11679 12492 11688
rect 12440 11645 12449 11679
rect 12449 11645 12483 11679
rect 12483 11645 12492 11679
rect 12440 11636 12492 11645
rect 13728 11679 13780 11688
rect 13728 11645 13737 11679
rect 13737 11645 13771 11679
rect 13771 11645 13780 11679
rect 13728 11636 13780 11645
rect 16672 11636 16724 11688
rect 17868 11636 17920 11688
rect 19708 11636 19760 11688
rect 19984 11636 20036 11688
rect 23756 11704 23808 11756
rect 24952 11704 25004 11756
rect 11060 11568 11112 11620
rect 8300 11500 8352 11552
rect 8944 11500 8996 11552
rect 9404 11543 9456 11552
rect 9404 11509 9413 11543
rect 9413 11509 9447 11543
rect 9447 11509 9456 11543
rect 9404 11500 9456 11509
rect 10416 11500 10468 11552
rect 11796 11500 11848 11552
rect 21732 11568 21784 11620
rect 24768 11679 24820 11688
rect 24768 11645 24777 11679
rect 24777 11645 24811 11679
rect 24811 11645 24820 11679
rect 24768 11636 24820 11645
rect 25780 11568 25832 11620
rect 17224 11500 17276 11552
rect 18512 11500 18564 11552
rect 19156 11500 19208 11552
rect 19432 11543 19484 11552
rect 19432 11509 19441 11543
rect 19441 11509 19475 11543
rect 19475 11509 19484 11543
rect 19432 11500 19484 11509
rect 21364 11500 21416 11552
rect 22284 11500 22336 11552
rect 23296 11500 23348 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 10600 11296 10652 11348
rect 12808 11228 12860 11280
rect 12900 11228 12952 11280
rect 12164 11160 12216 11212
rect 9036 11092 9088 11144
rect 11060 11092 11112 11144
rect 12532 11092 12584 11144
rect 12900 11092 12952 11144
rect 15292 11296 15344 11348
rect 15384 11296 15436 11348
rect 16304 11296 16356 11348
rect 17224 11339 17276 11348
rect 17224 11305 17233 11339
rect 17233 11305 17267 11339
rect 17267 11305 17276 11339
rect 17224 11296 17276 11305
rect 21824 11296 21876 11348
rect 13084 11228 13136 11280
rect 13360 11228 13412 11280
rect 13544 11160 13596 11212
rect 14004 11228 14056 11280
rect 14188 11228 14240 11280
rect 14740 11228 14792 11280
rect 16672 11271 16724 11280
rect 16672 11237 16681 11271
rect 16681 11237 16715 11271
rect 16715 11237 16724 11271
rect 16672 11228 16724 11237
rect 17868 11271 17920 11280
rect 17868 11237 17877 11271
rect 17877 11237 17911 11271
rect 17911 11237 17920 11271
rect 17868 11228 17920 11237
rect 20628 11228 20680 11280
rect 22560 11228 22612 11280
rect 23572 11296 23624 11348
rect 16948 11160 17000 11212
rect 18604 11203 18656 11212
rect 18604 11169 18613 11203
rect 18613 11169 18647 11203
rect 18647 11169 18656 11203
rect 18604 11160 18656 11169
rect 10416 11024 10468 11076
rect 9680 10956 9732 11008
rect 10876 10999 10928 11008
rect 10876 10965 10885 10999
rect 10885 10965 10919 10999
rect 10919 10965 10928 10999
rect 10876 10956 10928 10965
rect 11244 10956 11296 11008
rect 12256 11024 12308 11076
rect 13728 11024 13780 11076
rect 14004 11024 14056 11076
rect 16212 11092 16264 11144
rect 17500 11092 17552 11144
rect 19984 11135 20036 11144
rect 19984 11101 19993 11135
rect 19993 11101 20027 11135
rect 20027 11101 20036 11135
rect 19984 11092 20036 11101
rect 20996 11160 21048 11212
rect 25504 11228 25556 11280
rect 20720 11092 20772 11144
rect 21180 11092 21232 11144
rect 23296 11203 23348 11212
rect 23296 11169 23305 11203
rect 23305 11169 23339 11203
rect 23339 11169 23348 11203
rect 23296 11160 23348 11169
rect 21732 11135 21784 11144
rect 21732 11101 21741 11135
rect 21741 11101 21775 11135
rect 21775 11101 21784 11135
rect 21732 11092 21784 11101
rect 21824 11092 21876 11144
rect 22284 11092 22336 11144
rect 14280 10999 14332 11008
rect 14280 10965 14289 10999
rect 14289 10965 14323 10999
rect 14323 10965 14332 10999
rect 14280 10956 14332 10965
rect 15200 11067 15252 11076
rect 15200 11033 15209 11067
rect 15209 11033 15243 11067
rect 15243 11033 15252 11067
rect 15200 11024 15252 11033
rect 15292 11024 15344 11076
rect 15476 10956 15528 11008
rect 17408 11024 17460 11076
rect 19340 10956 19392 11008
rect 20812 11024 20864 11076
rect 20996 11024 21048 11076
rect 23940 11092 23992 11144
rect 25044 11024 25096 11076
rect 19800 10956 19852 11008
rect 20168 10956 20220 11008
rect 24492 10956 24544 11008
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 9956 10795 10008 10804
rect 9956 10761 9965 10795
rect 9965 10761 9999 10795
rect 9999 10761 10008 10795
rect 9956 10752 10008 10761
rect 12348 10795 12400 10804
rect 12348 10761 12357 10795
rect 12357 10761 12391 10795
rect 12391 10761 12400 10795
rect 12348 10752 12400 10761
rect 12716 10795 12768 10804
rect 12716 10761 12725 10795
rect 12725 10761 12759 10795
rect 12759 10761 12768 10795
rect 12716 10752 12768 10761
rect 7104 10412 7156 10464
rect 10416 10684 10468 10736
rect 10876 10616 10928 10668
rect 12808 10659 12860 10668
rect 12808 10625 12817 10659
rect 12817 10625 12851 10659
rect 12851 10625 12860 10659
rect 12808 10616 12860 10625
rect 12716 10548 12768 10600
rect 13452 10684 13504 10736
rect 15384 10684 15436 10736
rect 17224 10752 17276 10804
rect 17684 10752 17736 10804
rect 18420 10752 18472 10804
rect 18880 10752 18932 10804
rect 20168 10752 20220 10804
rect 17776 10684 17828 10736
rect 18328 10684 18380 10736
rect 18604 10684 18656 10736
rect 21272 10752 21324 10804
rect 22008 10752 22060 10804
rect 10416 10523 10468 10532
rect 10416 10489 10425 10523
rect 10425 10489 10459 10523
rect 10459 10489 10468 10523
rect 10416 10480 10468 10489
rect 9036 10412 9088 10464
rect 11244 10455 11296 10464
rect 11244 10421 11253 10455
rect 11253 10421 11287 10455
rect 11287 10421 11296 10455
rect 11244 10412 11296 10421
rect 12256 10480 12308 10532
rect 14004 10548 14056 10600
rect 14464 10591 14516 10600
rect 14464 10557 14473 10591
rect 14473 10557 14507 10591
rect 14507 10557 14516 10591
rect 14464 10548 14516 10557
rect 16856 10616 16908 10668
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 18788 10616 18840 10668
rect 19984 10659 20036 10668
rect 19984 10625 19993 10659
rect 19993 10625 20027 10659
rect 20027 10625 20036 10659
rect 19984 10616 20036 10625
rect 21088 10659 21140 10668
rect 21088 10625 21097 10659
rect 21097 10625 21131 10659
rect 21131 10625 21140 10659
rect 21088 10616 21140 10625
rect 16488 10548 16540 10600
rect 13636 10480 13688 10532
rect 15384 10480 15436 10532
rect 20076 10548 20128 10600
rect 20628 10548 20680 10600
rect 21272 10591 21324 10600
rect 21272 10557 21281 10591
rect 21281 10557 21315 10591
rect 21315 10557 21324 10591
rect 21272 10548 21324 10557
rect 23664 10752 23716 10804
rect 23388 10727 23440 10736
rect 23388 10693 23397 10727
rect 23397 10693 23431 10727
rect 23431 10693 23440 10727
rect 23388 10684 23440 10693
rect 22652 10616 22704 10668
rect 22468 10548 22520 10600
rect 11888 10412 11940 10464
rect 17684 10455 17736 10464
rect 17684 10421 17693 10455
rect 17693 10421 17727 10455
rect 17727 10421 17736 10455
rect 17684 10412 17736 10421
rect 18052 10412 18104 10464
rect 19524 10455 19576 10464
rect 19524 10421 19533 10455
rect 19533 10421 19567 10455
rect 19567 10421 19576 10455
rect 19524 10412 19576 10421
rect 22192 10480 22244 10532
rect 24400 10480 24452 10532
rect 21824 10412 21876 10464
rect 22100 10412 22152 10464
rect 23388 10412 23440 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 11060 10251 11112 10260
rect 11060 10217 11069 10251
rect 11069 10217 11103 10251
rect 11103 10217 11112 10251
rect 11060 10208 11112 10217
rect 11612 10251 11664 10260
rect 11612 10217 11621 10251
rect 11621 10217 11655 10251
rect 11655 10217 11664 10251
rect 11612 10208 11664 10217
rect 12072 10208 12124 10260
rect 13636 10208 13688 10260
rect 13912 10208 13964 10260
rect 14096 10208 14148 10260
rect 15660 10251 15712 10260
rect 15660 10217 15669 10251
rect 15669 10217 15703 10251
rect 15703 10217 15712 10251
rect 15660 10208 15712 10217
rect 19340 10208 19392 10260
rect 19524 10208 19576 10260
rect 9128 10072 9180 10124
rect 9956 10072 10008 10124
rect 12532 10140 12584 10192
rect 14832 10140 14884 10192
rect 17592 10140 17644 10192
rect 18328 10140 18380 10192
rect 11980 10072 12032 10124
rect 13544 10072 13596 10124
rect 15016 10115 15068 10124
rect 9036 10004 9088 10056
rect 12716 10004 12768 10056
rect 10324 9936 10376 9988
rect 12348 9936 12400 9988
rect 12532 9936 12584 9988
rect 15016 10081 15025 10115
rect 15025 10081 15059 10115
rect 15059 10081 15068 10115
rect 15016 10072 15068 10081
rect 14556 10004 14608 10056
rect 15844 10072 15896 10124
rect 20352 10140 20404 10192
rect 22008 10208 22060 10260
rect 24584 10251 24636 10260
rect 24584 10217 24593 10251
rect 24593 10217 24627 10251
rect 24627 10217 24636 10251
rect 24584 10208 24636 10217
rect 24492 10140 24544 10192
rect 15660 9936 15712 9988
rect 7104 9868 7156 9920
rect 11888 9868 11940 9920
rect 12808 9868 12860 9920
rect 14740 9868 14792 9920
rect 15476 9868 15528 9920
rect 15844 9911 15896 9920
rect 15844 9877 15853 9911
rect 15853 9877 15887 9911
rect 15887 9877 15896 9911
rect 15844 9868 15896 9877
rect 19248 10072 19300 10124
rect 19340 10072 19392 10124
rect 20260 10072 20312 10124
rect 22008 10072 22060 10124
rect 23388 10115 23440 10124
rect 23388 10081 23397 10115
rect 23397 10081 23431 10115
rect 23431 10081 23440 10115
rect 23388 10072 23440 10081
rect 16948 10004 17000 10056
rect 22100 10004 22152 10056
rect 22744 10004 22796 10056
rect 19064 9936 19116 9988
rect 20444 9936 20496 9988
rect 20720 9936 20772 9988
rect 20904 9936 20956 9988
rect 16764 9868 16816 9920
rect 17592 9868 17644 9920
rect 18512 9868 18564 9920
rect 19708 9868 19760 9920
rect 19800 9868 19852 9920
rect 20168 9911 20220 9920
rect 20168 9877 20177 9911
rect 20177 9877 20211 9911
rect 20211 9877 20220 9911
rect 20168 9868 20220 9877
rect 20628 9868 20680 9920
rect 24676 9868 24728 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 10968 9664 11020 9716
rect 12716 9664 12768 9716
rect 14556 9664 14608 9716
rect 15844 9664 15896 9716
rect 20168 9664 20220 9716
rect 20260 9664 20312 9716
rect 10508 9596 10560 9648
rect 12256 9596 12308 9648
rect 12440 9596 12492 9648
rect 11704 9571 11756 9580
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 15384 9528 15436 9580
rect 12348 9460 12400 9512
rect 13820 9392 13872 9444
rect 14096 9460 14148 9512
rect 14556 9503 14608 9512
rect 14556 9469 14565 9503
rect 14565 9469 14599 9503
rect 14599 9469 14608 9503
rect 14556 9460 14608 9469
rect 15568 9503 15620 9512
rect 15568 9469 15577 9503
rect 15577 9469 15611 9503
rect 15611 9469 15620 9503
rect 15568 9460 15620 9469
rect 15752 9503 15804 9512
rect 15752 9469 15761 9503
rect 15761 9469 15795 9503
rect 15795 9469 15804 9503
rect 15752 9460 15804 9469
rect 14648 9392 14700 9444
rect 17500 9596 17552 9648
rect 18052 9596 18104 9648
rect 19064 9596 19116 9648
rect 20628 9596 20680 9648
rect 20260 9571 20312 9580
rect 20260 9537 20269 9571
rect 20269 9537 20303 9571
rect 20303 9537 20312 9571
rect 20260 9528 20312 9537
rect 21088 9664 21140 9716
rect 21456 9596 21508 9648
rect 16948 9460 17000 9512
rect 18880 9460 18932 9512
rect 21088 9460 21140 9512
rect 21180 9503 21232 9512
rect 21180 9469 21189 9503
rect 21189 9469 21223 9503
rect 21223 9469 21232 9503
rect 21180 9460 21232 9469
rect 22100 9528 22152 9580
rect 22652 9571 22704 9580
rect 22652 9537 22661 9571
rect 22661 9537 22695 9571
rect 22695 9537 22704 9571
rect 22652 9528 22704 9537
rect 24032 9528 24084 9580
rect 23388 9460 23440 9512
rect 24400 9460 24452 9512
rect 22652 9392 22704 9444
rect 12348 9324 12400 9376
rect 13728 9324 13780 9376
rect 15660 9324 15712 9376
rect 15936 9324 15988 9376
rect 16856 9367 16908 9376
rect 16856 9333 16865 9367
rect 16865 9333 16899 9367
rect 16899 9333 16908 9367
rect 16856 9324 16908 9333
rect 17132 9324 17184 9376
rect 17592 9367 17644 9376
rect 17592 9333 17622 9367
rect 17622 9333 17644 9367
rect 17592 9324 17644 9333
rect 17960 9324 18012 9376
rect 18880 9324 18932 9376
rect 19800 9324 19852 9376
rect 22468 9324 22520 9376
rect 24860 9367 24912 9376
rect 24860 9333 24869 9367
rect 24869 9333 24903 9367
rect 24903 9333 24912 9367
rect 24860 9324 24912 9333
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 10968 9120 11020 9172
rect 11888 9120 11940 9172
rect 12808 9120 12860 9172
rect 14648 9120 14700 9172
rect 15108 9120 15160 9172
rect 15292 9120 15344 9172
rect 17408 9120 17460 9172
rect 17500 9120 17552 9172
rect 20076 9120 20128 9172
rect 20904 9120 20956 9172
rect 13360 9052 13412 9104
rect 11704 8984 11756 9036
rect 11888 8984 11940 9036
rect 15568 9052 15620 9104
rect 15752 9052 15804 9104
rect 13544 9027 13596 9036
rect 13544 8993 13553 9027
rect 13553 8993 13587 9027
rect 13587 8993 13596 9027
rect 13544 8984 13596 8993
rect 14556 8984 14608 9036
rect 16488 9027 16540 9036
rect 16488 8993 16497 9027
rect 16497 8993 16531 9027
rect 16531 8993 16540 9027
rect 16488 8984 16540 8993
rect 2780 8916 2832 8968
rect 4804 8916 4856 8968
rect 10968 8916 11020 8968
rect 12440 8916 12492 8968
rect 15844 8916 15896 8968
rect 15936 8916 15988 8968
rect 17132 8916 17184 8968
rect 19616 9052 19668 9104
rect 17960 8984 18012 9036
rect 24860 9052 24912 9104
rect 19616 8959 19668 8968
rect 19616 8925 19625 8959
rect 19625 8925 19659 8959
rect 19659 8925 19668 8959
rect 19616 8916 19668 8925
rect 9680 8848 9732 8900
rect 2412 8780 2464 8832
rect 8576 8780 8628 8832
rect 10968 8780 11020 8832
rect 14648 8823 14700 8832
rect 14648 8789 14657 8823
rect 14657 8789 14691 8823
rect 14691 8789 14700 8823
rect 14648 8780 14700 8789
rect 14832 8780 14884 8832
rect 15016 8780 15068 8832
rect 15384 8823 15436 8832
rect 15384 8789 15393 8823
rect 15393 8789 15427 8823
rect 15427 8789 15436 8823
rect 15384 8780 15436 8789
rect 15660 8780 15712 8832
rect 16856 8780 16908 8832
rect 17500 8891 17552 8900
rect 17500 8857 17509 8891
rect 17509 8857 17543 8891
rect 17543 8857 17552 8891
rect 17500 8848 17552 8857
rect 18696 8891 18748 8900
rect 18696 8857 18705 8891
rect 18705 8857 18739 8891
rect 18739 8857 18748 8891
rect 18696 8848 18748 8857
rect 19340 8848 19392 8900
rect 19800 8848 19852 8900
rect 17776 8780 17828 8832
rect 21456 8780 21508 8832
rect 22652 8959 22704 8968
rect 22652 8925 22661 8959
rect 22661 8925 22695 8959
rect 22695 8925 22704 8959
rect 22652 8916 22704 8925
rect 24216 8916 24268 8968
rect 24952 8848 25004 8900
rect 24032 8780 24084 8832
rect 24584 8823 24636 8832
rect 24584 8789 24593 8823
rect 24593 8789 24627 8823
rect 24627 8789 24636 8823
rect 24584 8780 24636 8789
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 9680 8576 9732 8628
rect 9956 8576 10008 8628
rect 12624 8576 12676 8628
rect 12532 8508 12584 8560
rect 13728 8508 13780 8560
rect 14556 8576 14608 8628
rect 14096 8551 14148 8560
rect 14096 8517 14105 8551
rect 14105 8517 14139 8551
rect 14139 8517 14148 8551
rect 14096 8508 14148 8517
rect 16856 8508 16908 8560
rect 14648 8440 14700 8492
rect 15108 8440 15160 8492
rect 17224 8483 17276 8492
rect 17224 8449 17233 8483
rect 17233 8449 17267 8483
rect 17267 8449 17276 8483
rect 17224 8440 17276 8449
rect 11428 8372 11480 8424
rect 13360 8372 13412 8424
rect 18236 8440 18288 8492
rect 18420 8483 18472 8492
rect 18420 8449 18429 8483
rect 18429 8449 18463 8483
rect 18463 8449 18472 8483
rect 18420 8440 18472 8449
rect 12808 8304 12860 8356
rect 17408 8415 17460 8424
rect 17408 8381 17417 8415
rect 17417 8381 17451 8415
rect 17451 8381 17460 8415
rect 17408 8372 17460 8381
rect 17776 8304 17828 8356
rect 18880 8372 18932 8424
rect 11980 8236 12032 8288
rect 18236 8304 18288 8356
rect 18512 8304 18564 8356
rect 23664 8508 23716 8560
rect 22192 8483 22244 8492
rect 22192 8449 22201 8483
rect 22201 8449 22235 8483
rect 22235 8449 22244 8483
rect 22192 8440 22244 8449
rect 20536 8372 20588 8424
rect 22284 8372 22336 8424
rect 22468 8372 22520 8424
rect 24768 8415 24820 8424
rect 24768 8381 24777 8415
rect 24777 8381 24811 8415
rect 24811 8381 24820 8415
rect 24768 8372 24820 8381
rect 20812 8304 20864 8356
rect 17960 8236 18012 8288
rect 22560 8236 22612 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 11796 8032 11848 8084
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 16120 8032 16172 8084
rect 16396 8032 16448 8084
rect 17776 8032 17828 8084
rect 19064 8032 19116 8084
rect 8392 7896 8444 7948
rect 11428 7871 11480 7880
rect 11428 7837 11437 7871
rect 11437 7837 11471 7871
rect 11471 7837 11480 7871
rect 11428 7828 11480 7837
rect 10324 7760 10376 7812
rect 11980 7896 12032 7948
rect 14004 7896 14056 7948
rect 14832 7939 14884 7948
rect 14832 7905 14841 7939
rect 14841 7905 14875 7939
rect 14875 7905 14884 7939
rect 14832 7896 14884 7905
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 13728 7828 13780 7880
rect 14464 7828 14516 7880
rect 14648 7871 14700 7880
rect 14648 7837 14657 7871
rect 14657 7837 14691 7871
rect 14691 7837 14700 7871
rect 14648 7828 14700 7837
rect 18788 7964 18840 8016
rect 19616 7964 19668 8016
rect 21824 7964 21876 8016
rect 15752 7896 15804 7948
rect 25320 8032 25372 8084
rect 25044 7964 25096 8016
rect 22376 7939 22428 7948
rect 22376 7905 22385 7939
rect 22385 7905 22419 7939
rect 22419 7905 22428 7939
rect 22376 7896 22428 7905
rect 16580 7828 16632 7880
rect 17960 7828 18012 7880
rect 12624 7692 12676 7744
rect 13360 7692 13412 7744
rect 15292 7760 15344 7812
rect 15844 7760 15896 7812
rect 20720 7760 20772 7812
rect 14004 7692 14056 7744
rect 15200 7692 15252 7744
rect 15660 7692 15712 7744
rect 18788 7692 18840 7744
rect 19892 7735 19944 7744
rect 19892 7701 19901 7735
rect 19901 7701 19935 7735
rect 19935 7701 19944 7735
rect 19892 7692 19944 7701
rect 21824 7828 21876 7880
rect 22100 7871 22152 7880
rect 22100 7837 22109 7871
rect 22109 7837 22143 7871
rect 22143 7837 22152 7871
rect 22100 7828 22152 7837
rect 24032 7828 24084 7880
rect 24216 7828 24268 7880
rect 21640 7760 21692 7812
rect 22376 7692 22428 7744
rect 23388 7692 23440 7744
rect 23848 7735 23900 7744
rect 23848 7701 23857 7735
rect 23857 7701 23891 7735
rect 23891 7701 23900 7735
rect 23848 7692 23900 7701
rect 24216 7735 24268 7744
rect 24216 7701 24225 7735
rect 24225 7701 24259 7735
rect 24259 7701 24268 7735
rect 24216 7692 24268 7701
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 11980 7531 12032 7540
rect 11980 7497 11989 7531
rect 11989 7497 12023 7531
rect 12023 7497 12032 7531
rect 11980 7488 12032 7497
rect 12624 7531 12676 7540
rect 12624 7497 12633 7531
rect 12633 7497 12667 7531
rect 12667 7497 12676 7531
rect 12624 7488 12676 7497
rect 13636 7488 13688 7540
rect 18328 7488 18380 7540
rect 19064 7488 19116 7540
rect 23480 7488 23532 7540
rect 11520 7420 11572 7472
rect 12072 7420 12124 7472
rect 14280 7420 14332 7472
rect 14464 7420 14516 7472
rect 16304 7420 16356 7472
rect 18880 7420 18932 7472
rect 20352 7420 20404 7472
rect 19892 7352 19944 7404
rect 20720 7352 20772 7404
rect 21916 7352 21968 7404
rect 25136 7463 25188 7472
rect 25136 7429 25145 7463
rect 25145 7429 25179 7463
rect 25179 7429 25188 7463
rect 25136 7420 25188 7429
rect 9036 7327 9088 7336
rect 9036 7293 9045 7327
rect 9045 7293 9079 7327
rect 9079 7293 9088 7327
rect 9036 7284 9088 7293
rect 10968 7284 11020 7336
rect 11152 7284 11204 7336
rect 10784 7259 10836 7268
rect 10784 7225 10793 7259
rect 10793 7225 10827 7259
rect 10827 7225 10836 7259
rect 10784 7216 10836 7225
rect 13452 7148 13504 7200
rect 16672 7284 16724 7336
rect 17592 7284 17644 7336
rect 17776 7216 17828 7268
rect 15108 7148 15160 7200
rect 16672 7191 16724 7200
rect 16672 7157 16681 7191
rect 16681 7157 16715 7191
rect 16715 7157 16724 7191
rect 16672 7148 16724 7157
rect 17040 7148 17092 7200
rect 18512 7327 18564 7336
rect 18512 7293 18521 7327
rect 18521 7293 18555 7327
rect 18555 7293 18564 7327
rect 18512 7284 18564 7293
rect 19248 7284 19300 7336
rect 19800 7284 19852 7336
rect 23480 7352 23532 7404
rect 24860 7284 24912 7336
rect 23572 7216 23624 7268
rect 22836 7148 22888 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 12348 6944 12400 6996
rect 14832 6944 14884 6996
rect 11704 6808 11756 6860
rect 14188 6851 14240 6860
rect 14188 6817 14197 6851
rect 14197 6817 14231 6851
rect 14231 6817 14240 6851
rect 14648 6876 14700 6928
rect 14188 6808 14240 6817
rect 17408 6851 17460 6860
rect 17408 6817 17417 6851
rect 17417 6817 17451 6851
rect 17451 6817 17460 6851
rect 17408 6808 17460 6817
rect 17868 6808 17920 6860
rect 19892 6944 19944 6996
rect 20168 6944 20220 6996
rect 18512 6876 18564 6928
rect 19616 6876 19668 6928
rect 19800 6876 19852 6928
rect 23848 6876 23900 6928
rect 19892 6851 19944 6860
rect 19892 6817 19901 6851
rect 19901 6817 19935 6851
rect 19935 6817 19944 6851
rect 19892 6808 19944 6817
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 13728 6740 13780 6749
rect 15476 6783 15528 6792
rect 15476 6749 15485 6783
rect 15485 6749 15519 6783
rect 15519 6749 15528 6783
rect 15476 6740 15528 6749
rect 16948 6740 17000 6792
rect 11060 6715 11112 6724
rect 11060 6681 11069 6715
rect 11069 6681 11103 6715
rect 11103 6681 11112 6715
rect 11060 6672 11112 6681
rect 11520 6672 11572 6724
rect 14648 6715 14700 6724
rect 14648 6681 14657 6715
rect 14657 6681 14691 6715
rect 14691 6681 14700 6715
rect 14648 6672 14700 6681
rect 12440 6604 12492 6656
rect 13544 6647 13596 6656
rect 13544 6613 13553 6647
rect 13553 6613 13587 6647
rect 13587 6613 13596 6647
rect 13544 6604 13596 6613
rect 14280 6604 14332 6656
rect 16672 6672 16724 6724
rect 17868 6672 17920 6724
rect 19524 6740 19576 6792
rect 20444 6808 20496 6860
rect 20260 6740 20312 6792
rect 21548 6740 21600 6792
rect 21732 6740 21784 6792
rect 21916 6740 21968 6792
rect 23296 6808 23348 6860
rect 24032 6808 24084 6860
rect 24492 6808 24544 6860
rect 19524 6604 19576 6656
rect 19800 6647 19852 6656
rect 19800 6613 19809 6647
rect 19809 6613 19843 6647
rect 19843 6613 19852 6647
rect 19800 6604 19852 6613
rect 25136 6672 25188 6724
rect 23296 6604 23348 6656
rect 23388 6604 23440 6656
rect 24860 6604 24912 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 11152 6400 11204 6452
rect 12808 6443 12860 6452
rect 12808 6409 12817 6443
rect 12817 6409 12851 6443
rect 12851 6409 12860 6443
rect 12808 6400 12860 6409
rect 17868 6400 17920 6452
rect 18328 6400 18380 6452
rect 6368 6264 6420 6316
rect 11152 6264 11204 6316
rect 10968 6239 11020 6248
rect 10968 6205 10977 6239
rect 10977 6205 11011 6239
rect 11011 6205 11020 6239
rect 10968 6196 11020 6205
rect 12256 6239 12308 6248
rect 12256 6205 12265 6239
rect 12265 6205 12299 6239
rect 12299 6205 12308 6239
rect 12256 6196 12308 6205
rect 14004 6332 14056 6384
rect 19524 6400 19576 6452
rect 20352 6400 20404 6452
rect 12716 6264 12768 6316
rect 14188 6264 14240 6316
rect 2688 6128 2740 6180
rect 10324 6128 10376 6180
rect 13360 6128 13412 6180
rect 13636 6196 13688 6248
rect 16120 6239 16172 6248
rect 16120 6205 16129 6239
rect 16129 6205 16163 6239
rect 16163 6205 16172 6239
rect 16120 6196 16172 6205
rect 13728 6128 13780 6180
rect 17224 6307 17276 6316
rect 17224 6273 17233 6307
rect 17233 6273 17267 6307
rect 17267 6273 17276 6307
rect 17224 6264 17276 6273
rect 20444 6332 20496 6384
rect 22652 6400 22704 6452
rect 23756 6400 23808 6452
rect 17316 6196 17368 6248
rect 22560 6332 22612 6384
rect 22008 6307 22060 6316
rect 22008 6273 22017 6307
rect 22017 6273 22051 6307
rect 22051 6273 22060 6307
rect 22008 6264 22060 6273
rect 21732 6196 21784 6248
rect 23848 6196 23900 6248
rect 22008 6128 22060 6180
rect 24124 6264 24176 6316
rect 15200 6060 15252 6112
rect 15660 6060 15712 6112
rect 19616 6060 19668 6112
rect 19800 6060 19852 6112
rect 20260 6060 20312 6112
rect 23848 6060 23900 6112
rect 24124 6060 24176 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 11060 5856 11112 5908
rect 12256 5856 12308 5908
rect 14004 5856 14056 5908
rect 14372 5856 14424 5908
rect 11336 5788 11388 5840
rect 15936 5788 15988 5840
rect 10784 5720 10836 5772
rect 12164 5720 12216 5772
rect 9036 5652 9088 5704
rect 9588 5652 9640 5704
rect 11612 5652 11664 5704
rect 12532 5695 12584 5704
rect 12532 5661 12541 5695
rect 12541 5661 12575 5695
rect 12575 5661 12584 5695
rect 12532 5652 12584 5661
rect 15200 5763 15252 5772
rect 15200 5729 15209 5763
rect 15209 5729 15243 5763
rect 15243 5729 15252 5763
rect 15200 5720 15252 5729
rect 15384 5763 15436 5772
rect 15384 5729 15393 5763
rect 15393 5729 15427 5763
rect 15427 5729 15436 5763
rect 15384 5720 15436 5729
rect 15108 5652 15160 5704
rect 16948 5720 17000 5772
rect 17408 5856 17460 5908
rect 19984 5856 20036 5908
rect 21548 5856 21600 5908
rect 21916 5856 21968 5908
rect 25228 5899 25280 5908
rect 25228 5865 25237 5899
rect 25237 5865 25271 5899
rect 25271 5865 25280 5899
rect 25228 5856 25280 5865
rect 18788 5652 18840 5704
rect 11060 5584 11112 5636
rect 13452 5584 13504 5636
rect 16672 5584 16724 5636
rect 16856 5516 16908 5568
rect 19892 5763 19944 5772
rect 19892 5729 19901 5763
rect 19901 5729 19935 5763
rect 19935 5729 19944 5763
rect 19892 5720 19944 5729
rect 22008 5788 22060 5840
rect 20628 5652 20680 5704
rect 21456 5695 21508 5704
rect 21456 5661 21465 5695
rect 21465 5661 21499 5695
rect 21499 5661 21508 5695
rect 21456 5652 21508 5661
rect 22744 5652 22796 5704
rect 23848 5652 23900 5704
rect 23940 5652 23992 5704
rect 24584 5652 24636 5704
rect 20904 5516 20956 5568
rect 23756 5584 23808 5636
rect 25136 5584 25188 5636
rect 24584 5516 24636 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 3424 5312 3476 5364
rect 10692 5312 10744 5364
rect 11612 5312 11664 5364
rect 11060 5244 11112 5296
rect 11520 5287 11572 5296
rect 11520 5253 11529 5287
rect 11529 5253 11563 5287
rect 11563 5253 11572 5287
rect 11520 5244 11572 5253
rect 11704 5244 11756 5296
rect 13636 5312 13688 5364
rect 14188 5312 14240 5364
rect 17316 5312 17368 5364
rect 11428 5176 11480 5228
rect 14464 5244 14516 5296
rect 17868 5287 17920 5296
rect 17868 5253 17877 5287
rect 17877 5253 17911 5287
rect 17911 5253 17920 5287
rect 17868 5244 17920 5253
rect 11888 5151 11940 5160
rect 11888 5117 11897 5151
rect 11897 5117 11931 5151
rect 11931 5117 11940 5151
rect 11888 5108 11940 5117
rect 12072 5108 12124 5160
rect 18512 5176 18564 5228
rect 20168 5176 20220 5228
rect 20444 5312 20496 5364
rect 21916 5312 21968 5364
rect 20812 5244 20864 5296
rect 21088 5219 21140 5228
rect 21088 5185 21097 5219
rect 21097 5185 21131 5219
rect 21131 5185 21140 5219
rect 21088 5176 21140 5185
rect 21548 5287 21600 5296
rect 21548 5253 21557 5287
rect 21557 5253 21591 5287
rect 21591 5253 21600 5287
rect 21548 5244 21600 5253
rect 22008 5176 22060 5228
rect 22100 5219 22152 5228
rect 22100 5185 22109 5219
rect 22109 5185 22143 5219
rect 22143 5185 22152 5219
rect 22100 5176 22152 5185
rect 23756 5176 23808 5228
rect 15200 5108 15252 5160
rect 15752 5151 15804 5160
rect 15752 5117 15761 5151
rect 15761 5117 15795 5151
rect 15795 5117 15804 5151
rect 15752 5108 15804 5117
rect 21272 5108 21324 5160
rect 21548 5108 21600 5160
rect 23480 5108 23532 5160
rect 14924 5040 14976 5092
rect 18420 5040 18472 5092
rect 20168 5040 20220 5092
rect 24216 5040 24268 5092
rect 13912 4972 13964 5024
rect 15476 4972 15528 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 10140 4811 10192 4820
rect 10140 4777 10149 4811
rect 10149 4777 10183 4811
rect 10183 4777 10192 4811
rect 10140 4768 10192 4777
rect 11244 4768 11296 4820
rect 11428 4768 11480 4820
rect 11888 4768 11940 4820
rect 20168 4768 20220 4820
rect 21272 4811 21324 4820
rect 21272 4777 21281 4811
rect 21281 4777 21315 4811
rect 21315 4777 21324 4811
rect 21272 4768 21324 4777
rect 22376 4768 22428 4820
rect 1492 4632 1544 4684
rect 9588 4632 9640 4684
rect 1768 4607 1820 4616
rect 1768 4573 1777 4607
rect 1777 4573 1811 4607
rect 1811 4573 1820 4607
rect 1768 4564 1820 4573
rect 7104 4607 7156 4616
rect 7104 4573 7113 4607
rect 7113 4573 7147 4607
rect 7147 4573 7156 4607
rect 7104 4564 7156 4573
rect 11244 4632 11296 4684
rect 14924 4632 14976 4684
rect 15108 4675 15160 4684
rect 15108 4641 15117 4675
rect 15117 4641 15151 4675
rect 15151 4641 15160 4675
rect 15108 4632 15160 4641
rect 16856 4743 16908 4752
rect 16856 4709 16865 4743
rect 16865 4709 16899 4743
rect 16899 4709 16908 4743
rect 16856 4700 16908 4709
rect 15476 4632 15528 4684
rect 15844 4632 15896 4684
rect 18512 4632 18564 4684
rect 10692 4496 10744 4548
rect 14280 4564 14332 4616
rect 14740 4564 14792 4616
rect 11060 4428 11112 4480
rect 14924 4496 14976 4548
rect 15384 4539 15436 4548
rect 15384 4505 15393 4539
rect 15393 4505 15427 4539
rect 15427 4505 15436 4539
rect 15384 4496 15436 4505
rect 13452 4428 13504 4480
rect 14464 4428 14516 4480
rect 14556 4428 14608 4480
rect 15844 4496 15896 4548
rect 18328 4539 18380 4548
rect 18328 4505 18337 4539
rect 18337 4505 18371 4539
rect 18371 4505 18380 4539
rect 18328 4496 18380 4505
rect 21824 4607 21876 4616
rect 21824 4573 21833 4607
rect 21833 4573 21867 4607
rect 21867 4573 21876 4607
rect 21824 4564 21876 4573
rect 22008 4564 22060 4616
rect 24032 4700 24084 4752
rect 19708 4496 19760 4548
rect 19800 4539 19852 4548
rect 19800 4505 19809 4539
rect 19809 4505 19843 4539
rect 19843 4505 19852 4539
rect 19800 4496 19852 4505
rect 20260 4496 20312 4548
rect 16672 4428 16724 4480
rect 19984 4428 20036 4480
rect 23756 4471 23808 4480
rect 23756 4437 23765 4471
rect 23765 4437 23799 4471
rect 23799 4437 23808 4471
rect 23756 4428 23808 4437
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 1768 4224 1820 4276
rect 14556 4224 14608 4276
rect 15476 4224 15528 4276
rect 17224 4224 17276 4276
rect 20260 4224 20312 4276
rect 24676 4267 24728 4276
rect 24676 4233 24685 4267
rect 24685 4233 24719 4267
rect 24719 4233 24728 4267
rect 24676 4224 24728 4233
rect 1492 4088 1544 4140
rect 1860 4088 1912 4140
rect 4068 4088 4120 4140
rect 9220 4088 9272 4140
rect 2688 3995 2740 4004
rect 2688 3961 2697 3995
rect 2697 3961 2731 3995
rect 2731 3961 2740 3995
rect 2688 3952 2740 3961
rect 7288 3952 7340 4004
rect 10324 4063 10376 4072
rect 10324 4029 10333 4063
rect 10333 4029 10367 4063
rect 10367 4029 10376 4063
rect 10324 4020 10376 4029
rect 10600 4131 10652 4140
rect 10600 4097 10609 4131
rect 10609 4097 10643 4131
rect 10643 4097 10652 4131
rect 10600 4088 10652 4097
rect 12256 4131 12308 4140
rect 12256 4097 12265 4131
rect 12265 4097 12299 4131
rect 12299 4097 12308 4131
rect 12256 4088 12308 4097
rect 14188 4199 14240 4208
rect 14188 4165 14197 4199
rect 14197 4165 14231 4199
rect 14231 4165 14240 4199
rect 14188 4156 14240 4165
rect 15568 4156 15620 4208
rect 13360 4088 13412 4140
rect 13912 4131 13964 4140
rect 13912 4097 13921 4131
rect 13921 4097 13955 4131
rect 13955 4097 13964 4131
rect 13912 4088 13964 4097
rect 12624 4020 12676 4072
rect 11704 3952 11756 4004
rect 4068 3884 4120 3936
rect 4804 3927 4856 3936
rect 4804 3893 4813 3927
rect 4813 3893 4847 3927
rect 4847 3893 4856 3927
rect 4804 3884 4856 3893
rect 5264 3884 5316 3936
rect 7012 3927 7064 3936
rect 7012 3893 7021 3927
rect 7021 3893 7055 3927
rect 7055 3893 7064 3927
rect 7012 3884 7064 3893
rect 9220 3884 9272 3936
rect 10048 3927 10100 3936
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 12164 3884 12216 3936
rect 16212 4020 16264 4072
rect 17776 4088 17828 4140
rect 20904 4131 20956 4140
rect 20904 4097 20913 4131
rect 20913 4097 20947 4131
rect 20947 4097 20956 4131
rect 20904 4088 20956 4097
rect 20996 4131 21048 4140
rect 20996 4097 21005 4131
rect 21005 4097 21039 4131
rect 21039 4097 21048 4131
rect 20996 4088 21048 4097
rect 21824 4131 21876 4140
rect 21824 4097 21833 4131
rect 21833 4097 21867 4131
rect 21867 4097 21876 4131
rect 21824 4088 21876 4097
rect 22008 4088 22060 4140
rect 18420 4020 18472 4072
rect 21272 4020 21324 4072
rect 21916 4020 21968 4072
rect 24124 4063 24176 4072
rect 24124 4029 24133 4063
rect 24133 4029 24167 4063
rect 24167 4029 24176 4063
rect 24124 4020 24176 4029
rect 19064 3952 19116 4004
rect 22560 3952 22612 4004
rect 17500 3884 17552 3936
rect 19156 3884 19208 3936
rect 19892 3884 19944 3936
rect 21456 3884 21508 3936
rect 21916 3884 21968 3936
rect 22100 3884 22152 3936
rect 23756 3884 23808 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 3332 3680 3384 3732
rect 7840 3680 7892 3732
rect 8392 3723 8444 3732
rect 8392 3689 8401 3723
rect 8401 3689 8435 3723
rect 8435 3689 8444 3723
rect 8392 3680 8444 3689
rect 10508 3680 10560 3732
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 6368 3655 6420 3664
rect 6368 3621 6377 3655
rect 6377 3621 6411 3655
rect 6411 3621 6420 3655
rect 6368 3612 6420 3621
rect 8852 3612 8904 3664
rect 13820 3680 13872 3732
rect 14924 3680 14976 3732
rect 18512 3680 18564 3732
rect 20260 3680 20312 3732
rect 21548 3680 21600 3732
rect 22652 3680 22704 3732
rect 8392 3544 8444 3596
rect 10048 3544 10100 3596
rect 12532 3544 12584 3596
rect 12808 3587 12860 3596
rect 12808 3553 12817 3587
rect 12817 3553 12851 3587
rect 12851 3553 12860 3587
rect 12808 3544 12860 3553
rect 2228 3476 2280 3528
rect 4436 3519 4488 3528
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 4804 3476 4856 3528
rect 7012 3476 7064 3528
rect 8484 3476 8536 3528
rect 7380 3408 7432 3460
rect 10692 3476 10744 3528
rect 14372 3612 14424 3664
rect 17408 3612 17460 3664
rect 18328 3612 18380 3664
rect 18788 3612 18840 3664
rect 14004 3544 14056 3596
rect 15476 3544 15528 3596
rect 17684 3544 17736 3596
rect 18696 3544 18748 3596
rect 16028 3476 16080 3528
rect 19524 3544 19576 3596
rect 19340 3476 19392 3528
rect 15016 3408 15068 3460
rect 3332 3383 3384 3392
rect 3332 3349 3341 3383
rect 3341 3349 3375 3383
rect 3375 3349 3384 3383
rect 3332 3340 3384 3349
rect 3792 3383 3844 3392
rect 3792 3349 3801 3383
rect 3801 3349 3835 3383
rect 3835 3349 3844 3383
rect 3792 3340 3844 3349
rect 6276 3340 6328 3392
rect 7748 3383 7800 3392
rect 7748 3349 7757 3383
rect 7757 3349 7791 3383
rect 7791 3349 7800 3383
rect 7748 3340 7800 3349
rect 9312 3340 9364 3392
rect 9588 3340 9640 3392
rect 10324 3340 10376 3392
rect 17132 3408 17184 3460
rect 17684 3408 17736 3460
rect 20076 3544 20128 3596
rect 21364 3519 21416 3528
rect 21364 3485 21373 3519
rect 21373 3485 21407 3519
rect 21407 3485 21416 3519
rect 21364 3476 21416 3485
rect 22744 3544 22796 3596
rect 24032 3519 24084 3528
rect 24032 3485 24041 3519
rect 24041 3485 24075 3519
rect 24075 3485 24084 3519
rect 24032 3476 24084 3485
rect 24308 3476 24360 3528
rect 24584 3519 24636 3528
rect 24584 3485 24593 3519
rect 24593 3485 24627 3519
rect 24627 3485 24636 3519
rect 24584 3476 24636 3485
rect 21640 3408 21692 3460
rect 22836 3408 22888 3460
rect 23020 3408 23072 3460
rect 23756 3408 23808 3460
rect 16396 3340 16448 3392
rect 20444 3340 20496 3392
rect 20536 3340 20588 3392
rect 23112 3340 23164 3392
rect 24584 3340 24636 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 9128 3136 9180 3188
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 10324 3179 10376 3188
rect 10324 3145 10333 3179
rect 10333 3145 10367 3179
rect 10367 3145 10376 3179
rect 10324 3136 10376 3145
rect 11336 3136 11388 3188
rect 13912 3136 13964 3188
rect 14188 3136 14240 3188
rect 16488 3136 16540 3188
rect 17868 3136 17920 3188
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 3700 3043 3752 3052
rect 3700 3009 3709 3043
rect 3709 3009 3743 3043
rect 3743 3009 3752 3043
rect 3700 3000 3752 3009
rect 5448 3043 5500 3052
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 5448 3000 5500 3009
rect 6644 3000 6696 3052
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 10324 3000 10376 3052
rect 2596 2932 2648 2984
rect 3332 2932 3384 2984
rect 5172 2975 5224 2984
rect 5172 2941 5181 2975
rect 5181 2941 5215 2975
rect 5215 2941 5224 2975
rect 5172 2932 5224 2941
rect 7748 2932 7800 2984
rect 11060 3000 11112 3052
rect 11796 3000 11848 3052
rect 16580 3068 16632 3120
rect 14096 3000 14148 3052
rect 18604 3000 18656 3052
rect 18972 3000 19024 3052
rect 11428 2932 11480 2984
rect 11704 2975 11756 2984
rect 11704 2941 11713 2975
rect 11713 2941 11747 2975
rect 11747 2941 11756 2975
rect 11704 2932 11756 2941
rect 13636 2975 13688 2984
rect 13636 2941 13645 2975
rect 13645 2941 13679 2975
rect 13679 2941 13688 2975
rect 13636 2932 13688 2941
rect 14740 2932 14792 2984
rect 15844 2932 15896 2984
rect 20536 3068 20588 3120
rect 20904 3136 20956 3188
rect 22192 3179 22244 3188
rect 22192 3145 22201 3179
rect 22201 3145 22235 3179
rect 22235 3145 22244 3179
rect 22192 3136 22244 3145
rect 22560 3136 22612 3188
rect 23664 3179 23716 3188
rect 23664 3145 23673 3179
rect 23673 3145 23707 3179
rect 23707 3145 23716 3179
rect 23664 3136 23716 3145
rect 24216 3179 24268 3188
rect 24216 3145 24225 3179
rect 24225 3145 24259 3179
rect 24259 3145 24268 3179
rect 24216 3136 24268 3145
rect 21916 3068 21968 3120
rect 22100 3111 22152 3120
rect 22100 3077 22109 3111
rect 22109 3077 22143 3111
rect 22143 3077 22152 3111
rect 22100 3068 22152 3077
rect 23020 3068 23072 3120
rect 23572 3111 23624 3120
rect 23572 3077 23581 3111
rect 23581 3077 23615 3111
rect 23615 3077 23624 3111
rect 23572 3068 23624 3077
rect 23756 3068 23808 3120
rect 21824 3000 21876 3052
rect 22928 3000 22980 3052
rect 25136 3043 25188 3052
rect 25136 3009 25145 3043
rect 25145 3009 25179 3043
rect 25179 3009 25188 3043
rect 25136 3000 25188 3009
rect 21364 2932 21416 2984
rect 23480 2932 23532 2984
rect 11152 2864 11204 2916
rect 15108 2864 15160 2916
rect 17224 2864 17276 2916
rect 19524 2864 19576 2916
rect 22100 2864 22152 2916
rect 24952 2907 25004 2916
rect 24952 2873 24961 2907
rect 24961 2873 24995 2907
rect 24995 2873 25004 2907
rect 24952 2864 25004 2873
rect 4436 2796 4488 2848
rect 4896 2839 4948 2848
rect 4896 2805 4905 2839
rect 4905 2805 4939 2839
rect 4939 2805 4948 2839
rect 4896 2796 4948 2805
rect 14832 2796 14884 2848
rect 16948 2796 17000 2848
rect 19892 2796 19944 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 8576 2592 8628 2644
rect 9772 2524 9824 2576
rect 5448 2499 5500 2508
rect 5448 2465 5457 2499
rect 5457 2465 5491 2499
rect 5491 2465 5500 2499
rect 5448 2456 5500 2465
rect 2964 2388 3016 2440
rect 4896 2388 4948 2440
rect 5540 2388 5592 2440
rect 5908 2320 5960 2372
rect 7840 2388 7892 2440
rect 8300 2388 8352 2440
rect 9312 2431 9364 2440
rect 9312 2397 9321 2431
rect 9321 2397 9355 2431
rect 9355 2397 9364 2431
rect 9312 2388 9364 2397
rect 15752 2592 15804 2644
rect 16028 2592 16080 2644
rect 13452 2524 13504 2576
rect 18696 2635 18748 2644
rect 18696 2601 18705 2635
rect 18705 2601 18739 2635
rect 18739 2601 18748 2635
rect 18696 2592 18748 2601
rect 22284 2592 22336 2644
rect 23204 2592 23256 2644
rect 12164 2388 12216 2440
rect 12440 2431 12492 2440
rect 12440 2397 12449 2431
rect 12449 2397 12483 2431
rect 12483 2397 12492 2431
rect 12440 2388 12492 2397
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 8852 2320 8904 2372
rect 9956 2320 10008 2372
rect 2596 2252 2648 2304
rect 4528 2295 4580 2304
rect 4528 2261 4537 2295
rect 4537 2261 4571 2295
rect 4571 2261 4580 2295
rect 4528 2252 4580 2261
rect 6644 2252 6696 2304
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 8392 2252 8444 2304
rect 11980 2320 12032 2372
rect 13268 2363 13320 2372
rect 13268 2329 13277 2363
rect 13277 2329 13311 2363
rect 13311 2329 13320 2363
rect 13268 2320 13320 2329
rect 14372 2456 14424 2508
rect 16028 2456 16080 2508
rect 14464 2431 14516 2440
rect 14464 2397 14473 2431
rect 14473 2397 14507 2431
rect 14507 2397 14516 2431
rect 14464 2388 14516 2397
rect 16120 2388 16172 2440
rect 17316 2499 17368 2508
rect 17316 2465 17325 2499
rect 17325 2465 17359 2499
rect 17359 2465 17368 2499
rect 17316 2456 17368 2465
rect 16764 2388 16816 2440
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 19892 2499 19944 2508
rect 19892 2465 19901 2499
rect 19901 2465 19935 2499
rect 19935 2465 19944 2499
rect 19892 2456 19944 2465
rect 22192 2524 22244 2576
rect 22100 2456 22152 2508
rect 24860 2456 24912 2508
rect 21456 2431 21508 2440
rect 21456 2397 21465 2431
rect 21465 2397 21499 2431
rect 21499 2397 21508 2431
rect 21456 2388 21508 2397
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 15660 2252 15712 2304
rect 21180 2252 21232 2304
rect 25136 2320 25188 2372
rect 23296 2252 23348 2304
rect 25228 2295 25280 2304
rect 25228 2261 25237 2295
rect 25237 2261 25271 2295
rect 25271 2261 25280 2295
rect 25228 2252 25280 2261
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 4528 2048 4580 2100
rect 8392 2048 8444 2100
rect 15200 2048 15252 2100
rect 11336 1980 11388 2032
rect 7840 1912 7892 1964
rect 17040 1912 17092 1964
rect 7104 1844 7156 1896
rect 12716 1844 12768 1896
rect 11244 1776 11296 1828
rect 25228 1776 25280 1828
<< metal2 >>
rect 1030 56200 1086 57000
rect 2410 56200 2466 57000
rect 3790 56200 3846 57000
rect 5170 56200 5226 57000
rect 6550 56200 6606 57000
rect 7930 56200 7986 57000
rect 9310 56200 9366 57000
rect 10690 56200 10746 57000
rect 12070 56200 12126 57000
rect 12176 56222 12388 56250
rect 1044 53650 1072 56200
rect 2424 54126 2452 56200
rect 2412 54120 2464 54126
rect 2412 54062 2464 54068
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 3804 53650 3832 56200
rect 4068 54188 4120 54194
rect 4068 54130 4120 54136
rect 4804 54188 4856 54194
rect 4804 54130 4856 54136
rect 1032 53644 1084 53650
rect 1032 53586 1084 53592
rect 3792 53644 3844 53650
rect 3792 53586 3844 53592
rect 4080 53242 4108 54130
rect 4160 53576 4212 53582
rect 4160 53518 4212 53524
rect 4068 53236 4120 53242
rect 4068 53178 4120 53184
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 4172 52698 4200 53518
rect 4160 52692 4212 52698
rect 4160 52634 4212 52640
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 4816 51406 4844 54130
rect 5184 54126 5212 56200
rect 5172 54120 5224 54126
rect 5172 54062 5224 54068
rect 6564 53650 6592 56200
rect 7944 55214 7972 56200
rect 7852 55186 7972 55214
rect 7380 54188 7432 54194
rect 7380 54130 7432 54136
rect 6552 53644 6604 53650
rect 6552 53586 6604 53592
rect 5540 53508 5592 53514
rect 5540 53450 5592 53456
rect 4804 51400 4856 51406
rect 4804 51342 4856 51348
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 5552 50522 5580 53450
rect 7392 51610 7420 54130
rect 7852 54126 7880 55186
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 9324 54126 9352 56200
rect 9588 54188 9640 54194
rect 9588 54130 9640 54136
rect 7840 54120 7892 54126
rect 7840 54062 7892 54068
rect 9312 54120 9364 54126
rect 9312 54062 9364 54068
rect 8576 54052 8628 54058
rect 8576 53994 8628 54000
rect 7840 53576 7892 53582
rect 7840 53518 7892 53524
rect 7748 53100 7800 53106
rect 7748 53042 7800 53048
rect 7380 51604 7432 51610
rect 7380 51546 7432 51552
rect 5540 50516 5592 50522
rect 5540 50458 5592 50464
rect 7760 50454 7788 53042
rect 7852 51542 7880 53518
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 7840 51536 7892 51542
rect 7840 51478 7892 51484
rect 8484 51400 8536 51406
rect 8484 51342 8536 51348
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 8392 50516 8444 50522
rect 8392 50458 8444 50464
rect 7748 50448 7800 50454
rect 7748 50390 7800 50396
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 7760 48142 7788 50390
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 8404 48686 8432 50458
rect 8300 48680 8352 48686
rect 8300 48622 8352 48628
rect 8392 48680 8444 48686
rect 8392 48622 8444 48628
rect 7748 48136 7800 48142
rect 7748 48078 7800 48084
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 7760 46034 7788 48078
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 8312 47462 8340 48622
rect 8300 47456 8352 47462
rect 8300 47398 8352 47404
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 8496 46170 8524 51342
rect 8588 50386 8616 53994
rect 9496 52488 9548 52494
rect 9496 52430 9548 52436
rect 8576 50380 8628 50386
rect 8576 50322 8628 50328
rect 8588 47734 8616 50322
rect 9128 48884 9180 48890
rect 9128 48826 9180 48832
rect 9140 48550 9168 48826
rect 9128 48544 9180 48550
rect 9128 48486 9180 48492
rect 8576 47728 8628 47734
rect 8576 47670 8628 47676
rect 8484 46164 8536 46170
rect 8484 46106 8536 46112
rect 7748 46028 7800 46034
rect 7748 45970 7800 45976
rect 7840 45960 7892 45966
rect 7840 45902 7892 45908
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 7852 38010 7880 45902
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 9140 44878 9168 48486
rect 9508 47802 9536 52430
rect 9600 50522 9628 54130
rect 10704 53718 10732 56200
rect 12084 56114 12112 56200
rect 12176 56114 12204 56222
rect 12084 56086 12204 56114
rect 11704 54188 11756 54194
rect 11704 54130 11756 54136
rect 10692 53712 10744 53718
rect 10692 53654 10744 53660
rect 10692 53576 10744 53582
rect 10692 53518 10744 53524
rect 10508 51400 10560 51406
rect 10508 51342 10560 51348
rect 9588 50516 9640 50522
rect 9588 50458 9640 50464
rect 9588 50244 9640 50250
rect 9588 50186 9640 50192
rect 9220 47796 9272 47802
rect 9220 47738 9272 47744
rect 9496 47796 9548 47802
rect 9496 47738 9548 47744
rect 9232 47054 9260 47738
rect 9496 47456 9548 47462
rect 9496 47398 9548 47404
rect 9220 47048 9272 47054
rect 9220 46990 9272 46996
rect 9128 44872 9180 44878
rect 9128 44814 9180 44820
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 9036 44328 9088 44334
rect 9036 44270 9088 44276
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 8944 42696 8996 42702
rect 8944 42638 8996 42644
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 7840 38004 7892 38010
rect 7840 37946 7892 37952
rect 8852 37868 8904 37874
rect 8852 37810 8904 37816
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2950 34235 3258 34244
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 8760 30728 8812 30734
rect 8760 30670 8812 30676
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 7656 30252 7708 30258
rect 7656 30194 7708 30200
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 3424 26784 3476 26790
rect 3424 26726 3476 26732
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2412 8832 2464 8838
rect 2792 8809 2820 8910
rect 2412 8774 2464 8780
rect 2778 8800 2834 8809
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 1504 4146 1532 4626
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1780 4282 1808 4558
rect 1768 4276 1820 4282
rect 1768 4218 1820 4224
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1504 800 1532 4082
rect 1872 800 1900 4082
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2240 800 2268 3470
rect 2424 3058 2452 8774
rect 2778 8735 2834 8744
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 2688 6180 2740 6186
rect 2688 6122 2740 6128
rect 2700 4010 2728 6122
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 2688 4004 2740 4010
rect 2688 3946 2740 3952
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 3344 3738 3372 16934
rect 3436 6497 3464 26726
rect 7564 24948 7616 24954
rect 7564 24890 7616 24896
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 4804 21140 4856 21146
rect 4804 21082 4856 21088
rect 3516 20868 3568 20874
rect 3516 20810 3568 20816
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3436 4185 3464 5306
rect 3422 4176 3478 4185
rect 3422 4111 3478 4120
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 3344 2990 3372 3334
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 2608 2310 2636 2926
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2596 2304 2648 2310
rect 2596 2246 2648 2252
rect 2608 800 2636 2246
rect 2976 800 3004 2382
rect 3344 800 3372 2926
rect 3528 1873 3556 20810
rect 3700 11892 3752 11898
rect 3700 11834 3752 11840
rect 3712 3058 3740 11834
rect 4816 8974 4844 21082
rect 6932 19310 6960 22374
rect 6552 19304 6604 19310
rect 6920 19304 6972 19310
rect 6604 19264 6684 19292
rect 6552 19246 6604 19252
rect 6656 18766 6684 19264
rect 6920 19246 6972 19252
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 6656 18222 6684 18702
rect 6644 18216 6696 18222
rect 6644 18158 6696 18164
rect 6552 16108 6604 16114
rect 6656 16096 6684 18158
rect 6604 16068 6684 16096
rect 6552 16050 6604 16056
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4080 3942 4108 4082
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3804 2938 3832 3334
rect 3712 2910 3832 2938
rect 3514 1864 3570 1873
rect 3514 1799 3570 1808
rect 3712 800 3740 2910
rect 4080 800 4108 3878
rect 4816 3534 4844 3878
rect 5184 3602 5212 15846
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4804 3528 4856 3534
rect 5276 3482 5304 3878
rect 4804 3470 4856 3476
rect 4448 2854 4476 3470
rect 4436 2848 4488 2854
rect 4436 2790 4488 2796
rect 4448 800 4476 2790
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 4540 2106 4568 2246
rect 4528 2100 4580 2106
rect 4528 2042 4580 2048
rect 4816 800 4844 3470
rect 5184 3454 5304 3482
rect 5184 2990 5212 3454
rect 5460 3058 5488 15574
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6472 13394 6500 14418
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6932 12782 6960 19246
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7208 17338 7236 17478
rect 7196 17332 7248 17338
rect 7196 17274 7248 17280
rect 7576 17066 7604 24890
rect 7668 17882 7696 30194
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 8576 26308 8628 26314
rect 8576 26250 8628 26256
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 7840 24200 7892 24206
rect 7840 24142 7892 24148
rect 7852 23730 7880 24142
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7840 23724 7892 23730
rect 7840 23666 7892 23672
rect 7852 22642 7880 23666
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7748 21344 7800 21350
rect 7852 21332 7880 22578
rect 8300 21888 8352 21894
rect 8300 21830 8352 21836
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8312 21554 8340 21830
rect 8300 21548 8352 21554
rect 8300 21490 8352 21496
rect 8312 21434 8340 21490
rect 8484 21480 8536 21486
rect 8312 21406 8432 21434
rect 8484 21422 8536 21428
rect 7800 21304 7880 21332
rect 8300 21344 8352 21350
rect 7748 21286 7800 21292
rect 8300 21286 8352 21292
rect 7760 20398 7788 21286
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8312 20534 8340 21286
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 7760 19922 7788 20334
rect 8404 19938 8432 21406
rect 8496 20398 8524 21422
rect 8484 20392 8536 20398
rect 8484 20334 8536 20340
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8496 20058 8524 20198
rect 8484 20052 8536 20058
rect 8484 19994 8536 20000
rect 8496 19938 8524 19994
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 8404 19910 8524 19938
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8404 19446 8432 19910
rect 8484 19780 8536 19786
rect 8484 19722 8536 19728
rect 8392 19440 8444 19446
rect 8392 19382 8444 19388
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 7932 18896 7984 18902
rect 7932 18838 7984 18844
rect 7944 18612 7972 18838
rect 8312 18834 8340 19110
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 7760 18584 7972 18612
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 7024 12306 7052 12786
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7116 9926 7144 10406
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6380 3670 6408 6258
rect 7116 4622 7144 9862
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7300 4010 7328 12786
rect 7564 12436 7616 12442
rect 7668 12434 7696 17478
rect 7760 12986 7788 18584
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8312 18358 8340 18634
rect 8496 18630 8524 19722
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 7840 17740 7892 17746
rect 7840 17682 7892 17688
rect 7852 14618 7880 17682
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8312 16402 8340 18294
rect 8312 16374 8432 16402
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 8312 14958 8340 16186
rect 8404 16182 8432 16374
rect 8392 16176 8444 16182
rect 8392 16118 8444 16124
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7852 13954 7880 14554
rect 8312 14482 8340 14758
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 8312 14074 8340 14418
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 7932 14000 7984 14006
rect 7852 13948 7932 13954
rect 7852 13942 7984 13948
rect 7852 13926 7972 13942
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7616 12406 7696 12434
rect 7564 12378 7616 12384
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 7024 3534 7052 3878
rect 7852 3738 7880 12718
rect 8220 12306 8248 12786
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 8312 11558 8340 14010
rect 8404 13530 8432 15982
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 8496 12782 8524 18566
rect 8588 17134 8616 26250
rect 8668 23180 8720 23186
rect 8668 23122 8720 23128
rect 8680 21350 8708 23122
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8668 20800 8720 20806
rect 8668 20742 8720 20748
rect 8680 18766 8708 20742
rect 8772 19514 8800 30670
rect 8864 29306 8892 37810
rect 8956 30122 8984 42638
rect 9048 34202 9076 44270
rect 9140 42158 9168 44814
rect 9232 44402 9260 46990
rect 9508 45082 9536 47398
rect 9496 45076 9548 45082
rect 9496 45018 9548 45024
rect 9600 44538 9628 50186
rect 10232 49156 10284 49162
rect 10232 49098 10284 49104
rect 9956 48612 10008 48618
rect 9956 48554 10008 48560
rect 9968 44946 9996 48554
rect 9956 44940 10008 44946
rect 9956 44882 10008 44888
rect 9680 44804 9732 44810
rect 9680 44746 9732 44752
rect 9588 44532 9640 44538
rect 9588 44474 9640 44480
rect 9220 44396 9272 44402
rect 9220 44338 9272 44344
rect 9692 42362 9720 44746
rect 10244 42770 10272 49098
rect 10416 46368 10468 46374
rect 10416 46310 10468 46316
rect 10428 44742 10456 46310
rect 10520 45558 10548 51342
rect 10704 49366 10732 53518
rect 10784 51332 10836 51338
rect 10784 51274 10836 51280
rect 10692 49360 10744 49366
rect 10692 49302 10744 49308
rect 10796 46714 10824 51274
rect 11716 49366 11744 54130
rect 12360 54126 12388 56222
rect 13450 56200 13506 57000
rect 13556 56222 13768 56250
rect 13464 56114 13492 56200
rect 13556 56114 13584 56222
rect 13464 56086 13584 56114
rect 13740 55214 13768 56222
rect 14830 56200 14886 57000
rect 16210 56200 16266 57000
rect 16316 56222 16528 56250
rect 13740 55186 13860 55214
rect 13832 54330 13860 55186
rect 13820 54324 13872 54330
rect 13820 54266 13872 54272
rect 14844 54194 14872 56200
rect 16224 56114 16252 56200
rect 16316 56114 16344 56222
rect 16224 56086 16344 56114
rect 14832 54188 14884 54194
rect 16500 54176 16528 56222
rect 17590 56200 17646 57000
rect 18970 56200 19026 57000
rect 20350 56200 20406 57000
rect 20456 56222 20668 56250
rect 17604 54194 17632 56200
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 18984 54330 19012 56200
rect 20364 56114 20392 56200
rect 20456 56114 20484 56222
rect 20364 56086 20484 56114
rect 18972 54324 19024 54330
rect 18972 54266 19024 54272
rect 16580 54188 16632 54194
rect 16500 54148 16580 54176
rect 14832 54130 14884 54136
rect 16580 54130 16632 54136
rect 17592 54188 17644 54194
rect 20640 54176 20668 56222
rect 21730 56200 21786 57000
rect 23110 56200 23166 57000
rect 24490 56200 24546 57000
rect 25870 56200 25926 57000
rect 21744 54194 21772 56200
rect 23124 54194 23152 56200
rect 23386 56128 23442 56137
rect 23386 56063 23442 56072
rect 20720 54188 20772 54194
rect 20640 54148 20720 54176
rect 17592 54130 17644 54136
rect 20720 54130 20772 54136
rect 21732 54188 21784 54194
rect 21732 54130 21784 54136
rect 23112 54188 23164 54194
rect 23112 54130 23164 54136
rect 12348 54120 12400 54126
rect 12348 54062 12400 54068
rect 13912 54052 13964 54058
rect 13912 53994 13964 54000
rect 15660 54052 15712 54058
rect 15660 53994 15712 54000
rect 20168 54052 20220 54058
rect 20168 53994 20220 54000
rect 12716 53984 12768 53990
rect 12716 53926 12768 53932
rect 11704 49360 11756 49366
rect 11704 49302 11756 49308
rect 10876 49156 10928 49162
rect 10876 49098 10928 49104
rect 10784 46708 10836 46714
rect 10784 46650 10836 46656
rect 10796 46594 10824 46650
rect 10612 46578 10824 46594
rect 10612 46572 10836 46578
rect 10612 46566 10784 46572
rect 10508 45552 10560 45558
rect 10508 45494 10560 45500
rect 10416 44736 10468 44742
rect 10416 44678 10468 44684
rect 10520 44266 10548 45494
rect 10508 44260 10560 44266
rect 10508 44202 10560 44208
rect 10232 42764 10284 42770
rect 10232 42706 10284 42712
rect 10612 42702 10640 46566
rect 10784 46514 10836 46520
rect 10784 46436 10836 46442
rect 10784 46378 10836 46384
rect 10796 44402 10824 46378
rect 10784 44396 10836 44402
rect 10784 44338 10836 44344
rect 10692 44192 10744 44198
rect 10692 44134 10744 44140
rect 10600 42696 10652 42702
rect 10600 42638 10652 42644
rect 9680 42356 9732 42362
rect 9680 42298 9732 42304
rect 10704 42158 10732 44134
rect 9128 42152 9180 42158
rect 9128 42094 9180 42100
rect 9772 42152 9824 42158
rect 9772 42094 9824 42100
rect 10692 42152 10744 42158
rect 10692 42094 10744 42100
rect 9784 35630 9812 42094
rect 10888 41818 10916 49098
rect 12624 48000 12676 48006
rect 12624 47942 12676 47948
rect 10968 47728 11020 47734
rect 10968 47670 11020 47676
rect 10980 46714 11008 47670
rect 10968 46708 11020 46714
rect 10968 46650 11020 46656
rect 12532 45960 12584 45966
rect 12532 45902 12584 45908
rect 12544 45558 12572 45902
rect 12636 45558 12664 47942
rect 12532 45552 12584 45558
rect 12532 45494 12584 45500
rect 12624 45552 12676 45558
rect 12624 45494 12676 45500
rect 12728 45490 12756 53926
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 13728 46980 13780 46986
rect 13728 46922 13780 46928
rect 13740 46646 13768 46922
rect 13728 46640 13780 46646
rect 13728 46582 13780 46588
rect 13924 46578 13952 53994
rect 15568 53984 15620 53990
rect 15568 53926 15620 53932
rect 13912 46572 13964 46578
rect 13912 46514 13964 46520
rect 15016 46368 15068 46374
rect 15016 46310 15068 46316
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 15028 46034 15056 46310
rect 15580 46102 15608 53926
rect 15568 46096 15620 46102
rect 15568 46038 15620 46044
rect 15016 46028 15068 46034
rect 15016 45970 15068 45976
rect 15108 45824 15160 45830
rect 15108 45766 15160 45772
rect 12716 45484 12768 45490
rect 12716 45426 12768 45432
rect 14556 45416 14608 45422
rect 14556 45358 14608 45364
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 11520 44804 11572 44810
rect 11520 44746 11572 44752
rect 10968 44192 11020 44198
rect 10968 44134 11020 44140
rect 10876 41812 10928 41818
rect 10876 41754 10928 41760
rect 10980 41682 11008 44134
rect 11532 42294 11560 44746
rect 11704 44736 11756 44742
rect 11704 44678 11756 44684
rect 11520 42288 11572 42294
rect 11520 42230 11572 42236
rect 11532 42022 11560 42230
rect 11716 42022 11744 44678
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 11520 42016 11572 42022
rect 11520 41958 11572 41964
rect 11704 42016 11756 42022
rect 11704 41958 11756 41964
rect 10968 41676 11020 41682
rect 10968 41618 11020 41624
rect 10232 41608 10284 41614
rect 10232 41550 10284 41556
rect 9680 35624 9732 35630
rect 9680 35566 9732 35572
rect 9772 35624 9824 35630
rect 9772 35566 9824 35572
rect 9036 34196 9088 34202
rect 9036 34138 9088 34144
rect 9220 33992 9272 33998
rect 9220 33934 9272 33940
rect 8944 30116 8996 30122
rect 8944 30058 8996 30064
rect 8852 29300 8904 29306
rect 8852 29242 8904 29248
rect 9232 23322 9260 33934
rect 9692 29238 9720 35566
rect 10244 30938 10272 41550
rect 11532 35766 11560 41958
rect 11716 35894 11744 41958
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 11716 35866 11836 35894
rect 11716 35834 11744 35866
rect 11704 35828 11756 35834
rect 11704 35770 11756 35776
rect 11520 35760 11572 35766
rect 11520 35702 11572 35708
rect 11808 35494 11836 35866
rect 12164 35760 12216 35766
rect 12164 35702 12216 35708
rect 11796 35488 11848 35494
rect 11796 35430 11848 35436
rect 11808 34066 11836 35430
rect 11796 34060 11848 34066
rect 11796 34002 11848 34008
rect 10232 30932 10284 30938
rect 10232 30874 10284 30880
rect 12176 30190 12204 35702
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 12624 32768 12676 32774
rect 12624 32710 12676 32716
rect 12532 31952 12584 31958
rect 12532 31894 12584 31900
rect 12544 31754 12572 31894
rect 12452 31726 12572 31754
rect 12072 30184 12124 30190
rect 12072 30126 12124 30132
rect 12164 30184 12216 30190
rect 12164 30126 12216 30132
rect 11520 30048 11572 30054
rect 11520 29990 11572 29996
rect 11428 29708 11480 29714
rect 11428 29650 11480 29656
rect 11336 29572 11388 29578
rect 11336 29514 11388 29520
rect 10416 29300 10468 29306
rect 10416 29242 10468 29248
rect 9680 29232 9732 29238
rect 9680 29174 9732 29180
rect 10232 29028 10284 29034
rect 10232 28970 10284 28976
rect 9680 28484 9732 28490
rect 9680 28426 9732 28432
rect 9312 27328 9364 27334
rect 9312 27270 9364 27276
rect 9324 26858 9352 27270
rect 9312 26852 9364 26858
rect 9312 26794 9364 26800
rect 9220 23316 9272 23322
rect 9220 23258 9272 23264
rect 9220 22024 9272 22030
rect 9220 21966 9272 21972
rect 9036 21616 9088 21622
rect 9036 21558 9088 21564
rect 9048 20806 9076 21558
rect 9036 20800 9088 20806
rect 9036 20742 9088 20748
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 9036 19372 9088 19378
rect 9036 19314 9088 19320
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8588 16794 8616 17070
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8680 16674 8708 18702
rect 8852 17604 8904 17610
rect 8852 17546 8904 17552
rect 8588 16646 8708 16674
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 8404 3738 8432 7890
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8496 3618 8524 12038
rect 8588 8838 8616 16646
rect 8668 16176 8720 16182
rect 8668 16118 8720 16124
rect 8680 15502 8708 16118
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8680 15094 8708 15438
rect 8668 15088 8720 15094
rect 8668 15030 8720 15036
rect 8680 14618 8708 15030
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8680 14006 8708 14554
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 8680 13530 8708 13942
rect 8864 13530 8892 17546
rect 9048 15706 9076 19314
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 9140 18086 9168 19110
rect 9128 18080 9180 18086
rect 9128 18022 9180 18028
rect 9232 17338 9260 21966
rect 9324 21486 9352 26794
rect 9404 24880 9456 24886
rect 9404 24822 9456 24828
rect 9416 24138 9444 24822
rect 9496 24268 9548 24274
rect 9496 24210 9548 24216
rect 9404 24132 9456 24138
rect 9404 24074 9456 24080
rect 9416 23730 9444 24074
rect 9404 23724 9456 23730
rect 9404 23666 9456 23672
rect 9416 23526 9444 23666
rect 9404 23520 9456 23526
rect 9508 23508 9536 24210
rect 9692 23866 9720 28426
rect 9772 27124 9824 27130
rect 9772 27066 9824 27072
rect 9784 26450 9812 27066
rect 9772 26444 9824 26450
rect 9772 26386 9824 26392
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 10048 23656 10100 23662
rect 10048 23598 10100 23604
rect 9508 23480 9628 23508
rect 9404 23462 9456 23468
rect 9416 23338 9444 23462
rect 9416 23310 9536 23338
rect 9404 23248 9456 23254
rect 9404 23190 9456 23196
rect 9312 21480 9364 21486
rect 9312 21422 9364 21428
rect 9312 20528 9364 20534
rect 9312 20470 9364 20476
rect 9324 20262 9352 20470
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9416 19786 9444 23190
rect 9508 22642 9536 23310
rect 9496 22636 9548 22642
rect 9496 22578 9548 22584
rect 9508 21894 9536 22578
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 9496 20392 9548 20398
rect 9496 20334 9548 20340
rect 9404 19780 9456 19786
rect 9404 19722 9456 19728
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9324 16250 9352 19246
rect 9508 18698 9536 20334
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 9508 18426 9536 18634
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9416 17338 9444 17478
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9600 17134 9628 23480
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9968 21010 9996 21490
rect 9956 21004 10008 21010
rect 9956 20946 10008 20952
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 9784 19922 9812 20878
rect 9956 20392 10008 20398
rect 9956 20334 10008 20340
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 9784 18154 9812 19858
rect 9968 18193 9996 20334
rect 10060 18970 10088 23598
rect 10140 23316 10192 23322
rect 10140 23258 10192 23264
rect 10152 20874 10180 23258
rect 10244 21690 10272 28970
rect 10324 25152 10376 25158
rect 10324 25094 10376 25100
rect 10336 23594 10364 25094
rect 10428 23866 10456 29242
rect 10876 29096 10928 29102
rect 10876 29038 10928 29044
rect 10888 28762 10916 29038
rect 10876 28756 10928 28762
rect 10876 28698 10928 28704
rect 11060 28076 11112 28082
rect 11060 28018 11112 28024
rect 10784 27940 10836 27946
rect 10784 27882 10836 27888
rect 10796 27538 10824 27882
rect 10784 27532 10836 27538
rect 10784 27474 10836 27480
rect 10876 27124 10928 27130
rect 10876 27066 10928 27072
rect 10692 25968 10744 25974
rect 10692 25910 10744 25916
rect 10416 23860 10468 23866
rect 10416 23802 10468 23808
rect 10324 23588 10376 23594
rect 10324 23530 10376 23536
rect 10336 23186 10364 23530
rect 10324 23180 10376 23186
rect 10324 23122 10376 23128
rect 10600 23180 10652 23186
rect 10600 23122 10652 23128
rect 10416 23044 10468 23050
rect 10416 22986 10468 22992
rect 10324 21888 10376 21894
rect 10324 21830 10376 21836
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 10140 20868 10192 20874
rect 10140 20810 10192 20816
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 10140 19372 10192 19378
rect 10140 19314 10192 19320
rect 10048 18964 10100 18970
rect 10048 18906 10100 18912
rect 9954 18184 10010 18193
rect 9772 18148 9824 18154
rect 9954 18119 10010 18128
rect 9772 18090 9824 18096
rect 9784 17678 9812 18090
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 9784 17270 9812 17614
rect 9968 17610 9996 18119
rect 9956 17604 10008 17610
rect 9956 17546 10008 17552
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9588 17128 9640 17134
rect 9588 17070 9640 17076
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 9036 14884 9088 14890
rect 9036 14826 9088 14832
rect 9048 14618 9076 14826
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8680 13258 8708 13466
rect 8668 13252 8720 13258
rect 8668 13194 8720 13200
rect 8680 11762 8708 13194
rect 8758 12880 8814 12889
rect 8758 12815 8814 12824
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8772 6914 8800 12815
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8404 3602 8524 3618
rect 8392 3596 8524 3602
rect 8444 3590 8524 3596
rect 8588 6886 8800 6914
rect 8392 3538 8444 3544
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 4908 2446 4936 2790
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5184 800 5212 2926
rect 5446 2544 5502 2553
rect 5446 2479 5448 2488
rect 5500 2479 5502 2488
rect 5448 2450 5500 2456
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5552 800 5580 2382
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 5920 800 5948 2314
rect 6288 800 6316 3334
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6656 2310 6684 2994
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 6656 800 6684 2246
rect 7024 800 7052 3470
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7392 3058 7420 3402
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 1902 7144 2246
rect 7104 1896 7156 1902
rect 7104 1838 7156 1844
rect 7392 800 7420 2994
rect 7760 2990 7788 3334
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7760 800 7788 2926
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 7852 1970 7880 2382
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 8312 1986 8340 2382
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 8404 2106 8432 2246
rect 8392 2100 8444 2106
rect 8392 2042 8444 2048
rect 7840 1964 7892 1970
rect 7840 1906 7892 1912
rect 8128 1958 8340 1986
rect 8128 800 8156 1958
rect 8496 800 8524 3470
rect 8588 2650 8616 6886
rect 8864 3670 8892 12582
rect 9048 12434 9076 14554
rect 9232 12986 9260 15370
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 9324 13462 9352 14282
rect 9312 13456 9364 13462
rect 9312 13398 9364 13404
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9048 12406 9168 12434
rect 8944 11552 8996 11558
rect 8996 11500 9076 11506
rect 8944 11494 9076 11500
rect 8956 11478 9076 11494
rect 9048 11150 9076 11478
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 9048 10470 9076 11086
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 9048 10062 9076 10406
rect 9140 10130 9168 12406
rect 9324 12306 9352 13398
rect 9416 12986 9444 17070
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9600 15570 9628 15982
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9600 15026 9628 15506
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9600 14074 9628 14350
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9600 13938 9628 14010
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9692 13274 9720 13330
rect 9692 13246 9812 13274
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9324 11898 9352 12242
rect 9416 12102 9444 12922
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9692 11898 9720 13126
rect 9784 12782 9812 13246
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9876 12434 9904 16390
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 10060 12986 10088 15302
rect 10152 15162 10180 19314
rect 10244 16454 10272 20334
rect 10336 16522 10364 21830
rect 10428 20602 10456 22986
rect 10508 22976 10560 22982
rect 10508 22918 10560 22924
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 10428 19786 10456 20198
rect 10416 19780 10468 19786
rect 10416 19722 10468 19728
rect 10428 19378 10456 19722
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 10520 18426 10548 22918
rect 10612 18834 10640 23122
rect 10704 21894 10732 25910
rect 10888 25362 10916 27066
rect 11072 26450 11100 28018
rect 11152 27056 11204 27062
rect 11152 26998 11204 27004
rect 11164 26586 11192 26998
rect 11348 26926 11376 29514
rect 11440 28626 11468 29650
rect 11428 28620 11480 28626
rect 11428 28562 11480 28568
rect 11440 27674 11468 28562
rect 11532 28422 11560 29990
rect 12084 29850 12112 30126
rect 12072 29844 12124 29850
rect 12072 29786 12124 29792
rect 12452 29306 12480 31726
rect 12636 29306 12664 32710
rect 13360 32360 13412 32366
rect 13360 32302 13412 32308
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 13372 31278 13400 32302
rect 13360 31272 13412 31278
rect 13360 31214 13412 31220
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 13372 30394 13400 31214
rect 13820 31136 13872 31142
rect 13820 31078 13872 31084
rect 13360 30388 13412 30394
rect 13360 30330 13412 30336
rect 12716 30320 12768 30326
rect 12716 30262 12768 30268
rect 12728 30190 12756 30262
rect 12716 30184 12768 30190
rect 12716 30126 12768 30132
rect 13360 30184 13412 30190
rect 13360 30126 13412 30132
rect 12728 29578 12756 30126
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 13372 29714 13400 30126
rect 13636 30048 13688 30054
rect 13636 29990 13688 29996
rect 13360 29708 13412 29714
rect 13360 29650 13412 29656
rect 12716 29572 12768 29578
rect 12716 29514 12768 29520
rect 12440 29300 12492 29306
rect 12440 29242 12492 29248
rect 12624 29300 12676 29306
rect 12624 29242 12676 29248
rect 13372 29170 13400 29650
rect 13360 29164 13412 29170
rect 13360 29106 13412 29112
rect 13648 29102 13676 29990
rect 13832 29850 13860 31078
rect 14096 30728 14148 30734
rect 14096 30670 14148 30676
rect 14108 30326 14136 30670
rect 14568 30326 14596 45358
rect 15120 44810 15148 45766
rect 15672 44946 15700 53994
rect 16948 53984 17000 53990
rect 16948 53926 17000 53932
rect 15752 46504 15804 46510
rect 15752 46446 15804 46452
rect 15660 44940 15712 44946
rect 15660 44882 15712 44888
rect 15108 44804 15160 44810
rect 15108 44746 15160 44752
rect 15568 42084 15620 42090
rect 15568 42026 15620 42032
rect 15384 33924 15436 33930
rect 15384 33866 15436 33872
rect 15396 32502 15424 33866
rect 15384 32496 15436 32502
rect 15384 32438 15436 32444
rect 14924 31408 14976 31414
rect 14924 31350 14976 31356
rect 14096 30320 14148 30326
rect 14096 30262 14148 30268
rect 14556 30320 14608 30326
rect 14556 30262 14608 30268
rect 13820 29844 13872 29850
rect 13820 29786 13872 29792
rect 13832 29306 13860 29786
rect 14936 29510 14964 31350
rect 15396 30938 15424 32438
rect 15384 30932 15436 30938
rect 15384 30874 15436 30880
rect 15396 30734 15424 30874
rect 15384 30728 15436 30734
rect 15384 30670 15436 30676
rect 15108 30660 15160 30666
rect 15108 30602 15160 30608
rect 14924 29504 14976 29510
rect 14924 29446 14976 29452
rect 13820 29300 13872 29306
rect 13820 29242 13872 29248
rect 13912 29300 13964 29306
rect 13912 29242 13964 29248
rect 13924 29186 13952 29242
rect 14936 29238 14964 29446
rect 13740 29158 13952 29186
rect 14924 29232 14976 29238
rect 14924 29174 14976 29180
rect 11796 29096 11848 29102
rect 11796 29038 11848 29044
rect 13636 29096 13688 29102
rect 13636 29038 13688 29044
rect 11704 28620 11756 28626
rect 11624 28580 11704 28608
rect 11624 28490 11652 28580
rect 11704 28562 11756 28568
rect 11612 28484 11664 28490
rect 11612 28426 11664 28432
rect 11520 28416 11572 28422
rect 11520 28358 11572 28364
rect 11428 27668 11480 27674
rect 11428 27610 11480 27616
rect 11336 26920 11388 26926
rect 11336 26862 11388 26868
rect 11152 26580 11204 26586
rect 11152 26522 11204 26528
rect 11060 26444 11112 26450
rect 11060 26386 11112 26392
rect 10876 25356 10928 25362
rect 10876 25298 10928 25304
rect 11072 24750 11100 26386
rect 11348 25838 11376 26862
rect 11336 25832 11388 25838
rect 11336 25774 11388 25780
rect 11152 24948 11204 24954
rect 11152 24890 11204 24896
rect 10876 24744 10928 24750
rect 10876 24686 10928 24692
rect 11060 24744 11112 24750
rect 11060 24686 11112 24692
rect 10888 24070 10916 24686
rect 11164 24614 11192 24890
rect 11060 24608 11112 24614
rect 11060 24550 11112 24556
rect 11152 24608 11204 24614
rect 11152 24550 11204 24556
rect 11072 24274 11100 24550
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 10876 24064 10928 24070
rect 10876 24006 10928 24012
rect 10888 23526 10916 24006
rect 10968 23656 11020 23662
rect 10968 23598 11020 23604
rect 10876 23520 10928 23526
rect 10876 23462 10928 23468
rect 10784 23112 10836 23118
rect 10784 23054 10836 23060
rect 10692 21888 10744 21894
rect 10692 21830 10744 21836
rect 10796 18970 10824 23054
rect 10980 21486 11008 23598
rect 11164 22574 11192 24550
rect 11336 22772 11388 22778
rect 11336 22714 11388 22720
rect 11152 22568 11204 22574
rect 11152 22510 11204 22516
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 11072 21690 11100 21830
rect 11060 21684 11112 21690
rect 11060 21626 11112 21632
rect 11152 21548 11204 21554
rect 11152 21490 11204 21496
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 10876 20868 10928 20874
rect 10876 20810 10928 20816
rect 10888 19718 10916 20810
rect 11060 19780 11112 19786
rect 11060 19722 11112 19728
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 10888 18834 10916 19654
rect 10968 19304 11020 19310
rect 11072 19292 11100 19722
rect 11020 19264 11100 19292
rect 10968 19246 11020 19252
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10416 18284 10468 18290
rect 10416 18226 10468 18232
rect 10324 16516 10376 16522
rect 10324 16458 10376 16464
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10230 14512 10286 14521
rect 10230 14447 10232 14456
rect 10284 14447 10286 14456
rect 10232 14418 10284 14424
rect 10244 13870 10272 14418
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 9784 12406 9904 12434
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9416 11558 9444 11698
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 9048 7342 9076 9998
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9048 5710 9076 7278
rect 9508 6914 9536 11698
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9692 8906 9720 10950
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9140 6886 9536 6914
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 8852 3664 8904 3670
rect 8852 3606 8904 3612
rect 9140 3194 9168 6886
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9600 4690 9628 5646
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9232 3942 9260 4082
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8852 2372 8904 2378
rect 8852 2314 8904 2320
rect 8864 800 8892 2314
rect 9232 800 9260 3878
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9324 2446 9352 3334
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 9600 800 9628 3334
rect 9692 3194 9720 8570
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9784 2582 9812 12406
rect 9968 10810 9996 12718
rect 10428 12714 10456 18226
rect 10416 12708 10468 12714
rect 10416 12650 10468 12656
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10428 11082 10456 11494
rect 10612 11354 10640 12038
rect 10796 11744 10824 18362
rect 10888 18154 10916 18566
rect 10876 18148 10928 18154
rect 10876 18090 10928 18096
rect 10980 17898 11008 19246
rect 11060 18896 11112 18902
rect 11060 18838 11112 18844
rect 11072 18630 11100 18838
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 10888 17870 11008 17898
rect 10888 11898 10916 17870
rect 11072 17610 11100 18022
rect 11060 17604 11112 17610
rect 11060 17546 11112 17552
rect 11072 17134 11100 17546
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 11164 15706 11192 21490
rect 11348 18290 11376 22714
rect 11532 22166 11560 28358
rect 11624 28218 11652 28426
rect 11612 28212 11664 28218
rect 11612 28154 11664 28160
rect 11704 28008 11756 28014
rect 11704 27950 11756 27956
rect 11716 27130 11744 27950
rect 11704 27124 11756 27130
rect 11704 27066 11756 27072
rect 11716 26994 11744 27066
rect 11704 26988 11756 26994
rect 11704 26930 11756 26936
rect 11612 26512 11664 26518
rect 11612 26454 11664 26460
rect 11624 23118 11652 26454
rect 11808 26314 11836 29038
rect 12164 29028 12216 29034
rect 12164 28970 12216 28976
rect 11980 26784 12032 26790
rect 11980 26726 12032 26732
rect 11796 26308 11848 26314
rect 11796 26250 11848 26256
rect 11704 25492 11756 25498
rect 11704 25434 11756 25440
rect 11716 23186 11744 25434
rect 11992 24138 12020 26726
rect 12176 24818 12204 28970
rect 13740 28914 13768 29158
rect 14648 29028 14700 29034
rect 14648 28970 14700 28976
rect 13648 28886 13768 28914
rect 14096 28960 14148 28966
rect 14096 28902 14148 28908
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 12716 28620 12768 28626
rect 12716 28562 12768 28568
rect 12728 27674 12756 28562
rect 13452 28144 13504 28150
rect 13452 28086 13504 28092
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 12716 27668 12768 27674
rect 12716 27610 12768 27616
rect 12624 27328 12676 27334
rect 12624 27270 12676 27276
rect 12636 26042 12664 27270
rect 12728 27130 12756 27610
rect 13084 27600 13136 27606
rect 13084 27542 13136 27548
rect 12716 27124 12768 27130
rect 12716 27066 12768 27072
rect 12624 26036 12676 26042
rect 12624 25978 12676 25984
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12164 24812 12216 24818
rect 12164 24754 12216 24760
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 11980 24132 12032 24138
rect 11980 24074 12032 24080
rect 11704 23180 11756 23186
rect 11704 23122 11756 23128
rect 11796 23180 11848 23186
rect 11796 23122 11848 23128
rect 11612 23112 11664 23118
rect 11612 23054 11664 23060
rect 11808 22506 11836 23122
rect 11796 22500 11848 22506
rect 11796 22442 11848 22448
rect 11520 22160 11572 22166
rect 11520 22102 11572 22108
rect 11992 19922 12020 24074
rect 12164 22976 12216 22982
rect 12164 22918 12216 22924
rect 12072 21616 12124 21622
rect 12072 21558 12124 21564
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 11716 19514 11744 19654
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11348 16794 11376 18226
rect 11716 17746 11744 18702
rect 11808 18358 11836 19450
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11532 17202 11560 17274
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11532 16998 11560 17138
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11348 16658 11376 16730
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11428 15088 11480 15094
rect 11428 15030 11480 15036
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11072 12986 11100 13806
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10980 12288 11008 12718
rect 11060 12300 11112 12306
rect 10980 12260 11060 12288
rect 11060 12242 11112 12248
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 11256 11762 11284 14894
rect 11440 12442 11468 15030
rect 11532 14822 11560 16934
rect 11612 16720 11664 16726
rect 11612 16662 11664 16668
rect 11624 16250 11652 16662
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11716 16182 11744 17682
rect 11992 16998 12020 17682
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11704 16176 11756 16182
rect 11704 16118 11756 16124
rect 11612 14884 11664 14890
rect 11612 14826 11664 14832
rect 11520 14816 11572 14822
rect 11520 14758 11572 14764
rect 11428 12436 11480 12442
rect 11428 12378 11480 12384
rect 10704 11716 10824 11744
rect 11244 11756 11296 11762
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10416 11076 10468 11082
rect 10416 11018 10468 11024
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 10428 10742 10456 11018
rect 10416 10736 10468 10742
rect 10416 10678 10468 10684
rect 10428 10538 10456 10678
rect 10416 10532 10468 10538
rect 10416 10474 10468 10480
rect 10428 10418 10456 10474
rect 10336 10390 10456 10418
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9968 8634 9996 10066
rect 10336 9994 10364 10390
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 10508 9648 10560 9654
rect 10508 9590 10560 9596
rect 10138 8936 10194 8945
rect 10138 8871 10194 8880
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 10152 4826 10180 8871
rect 10324 7812 10376 7818
rect 10324 7754 10376 7760
rect 10336 6186 10364 7754
rect 10324 6180 10376 6186
rect 10324 6122 10376 6128
rect 10140 4820 10192 4826
rect 10192 4780 10272 4808
rect 10140 4762 10192 4768
rect 10244 4060 10272 4780
rect 10324 4072 10376 4078
rect 10244 4032 10324 4060
rect 10324 4014 10376 4020
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10060 3602 10088 3878
rect 10520 3738 10548 9590
rect 10704 5370 10732 11716
rect 11244 11698 11296 11704
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 11072 11150 11100 11562
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 10888 10674 10916 10950
rect 10876 10668 10928 10674
rect 10876 10610 10928 10616
rect 11072 10266 11100 11086
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11256 10470 11284 10950
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 10980 9178 11008 9658
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10980 8974 11008 9114
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10980 7342 11008 8774
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 10784 7268 10836 7274
rect 10784 7210 10836 7216
rect 10796 5778 10824 7210
rect 10980 6254 11008 7278
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 11072 5914 11100 6666
rect 11164 6458 11192 7278
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 11072 5302 11100 5578
rect 11060 5296 11112 5302
rect 10598 5264 10654 5273
rect 11060 5238 11112 5244
rect 10598 5199 10654 5208
rect 10612 4146 10640 5199
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 10704 3534 10732 4490
rect 11072 4486 11100 5238
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 10336 3194 10364 3334
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 9956 2372 10008 2378
rect 9956 2314 10008 2320
rect 9968 800 9996 2314
rect 10336 800 10364 2994
rect 10704 800 10732 3470
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11072 800 11100 2994
rect 11164 2922 11192 6258
rect 11256 4826 11284 10406
rect 11624 10266 11652 14826
rect 11900 14482 11928 16730
rect 11992 15910 12020 16934
rect 12084 15978 12112 21558
rect 12176 18766 12204 22918
rect 12360 22642 12388 24210
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 12360 22114 12388 22578
rect 12360 22086 12480 22114
rect 12452 21486 12480 22086
rect 12440 21480 12492 21486
rect 12440 21422 12492 21428
rect 12544 21350 12572 25842
rect 12728 25430 12756 27066
rect 13096 26994 13124 27542
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 13084 26988 13136 26994
rect 13084 26930 13136 26936
rect 12716 25424 12768 25430
rect 12716 25366 12768 25372
rect 12728 25294 12756 25366
rect 12716 25288 12768 25294
rect 12716 25230 12768 25236
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12636 24410 12664 25094
rect 12728 24886 12756 25230
rect 12716 24880 12768 24886
rect 12716 24822 12768 24828
rect 12624 24404 12676 24410
rect 12624 24346 12676 24352
rect 12728 24138 12756 24822
rect 12820 24818 12848 26930
rect 13464 26926 13492 28086
rect 13648 27062 13676 28886
rect 13728 28756 13780 28762
rect 13728 28698 13780 28704
rect 13740 28218 13768 28698
rect 14108 28626 14136 28902
rect 14096 28620 14148 28626
rect 14096 28562 14148 28568
rect 13728 28212 13780 28218
rect 13728 28154 13780 28160
rect 13820 27872 13872 27878
rect 13820 27814 13872 27820
rect 13832 27402 13860 27814
rect 13820 27396 13872 27402
rect 13820 27338 13872 27344
rect 13728 27328 13780 27334
rect 13728 27270 13780 27276
rect 13636 27056 13688 27062
rect 13636 26998 13688 27004
rect 13452 26920 13504 26926
rect 13452 26862 13504 26868
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 13636 26580 13688 26586
rect 13636 26522 13688 26528
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 13360 25288 13412 25294
rect 13360 25230 13412 25236
rect 12808 24812 12860 24818
rect 12808 24754 12860 24760
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12900 24404 12952 24410
rect 12900 24346 12952 24352
rect 12716 24132 12768 24138
rect 12716 24074 12768 24080
rect 12912 23594 12940 24346
rect 12900 23588 12952 23594
rect 12900 23530 12952 23536
rect 12624 23520 12676 23526
rect 12624 23462 12676 23468
rect 12808 23520 12860 23526
rect 12808 23462 12860 23468
rect 12636 22098 12664 23462
rect 12716 23248 12768 23254
rect 12716 23190 12768 23196
rect 12624 22092 12676 22098
rect 12624 22034 12676 22040
rect 12728 21570 12756 23190
rect 12820 22166 12848 23462
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13372 22574 13400 25230
rect 13544 24880 13596 24886
rect 13544 24822 13596 24828
rect 13556 24410 13584 24822
rect 13544 24404 13596 24410
rect 13544 24346 13596 24352
rect 13648 23798 13676 26522
rect 13740 23798 13768 27270
rect 14108 25838 14136 28562
rect 14556 26376 14608 26382
rect 14556 26318 14608 26324
rect 14188 25968 14240 25974
rect 14188 25910 14240 25916
rect 14096 25832 14148 25838
rect 14096 25774 14148 25780
rect 13912 24744 13964 24750
rect 13912 24686 13964 24692
rect 13924 24070 13952 24686
rect 13912 24064 13964 24070
rect 13912 24006 13964 24012
rect 13636 23792 13688 23798
rect 13636 23734 13688 23740
rect 13728 23792 13780 23798
rect 13728 23734 13780 23740
rect 13924 23662 13952 24006
rect 14200 23866 14228 25910
rect 14568 25362 14596 26318
rect 14660 26042 14688 28970
rect 14936 28762 14964 29174
rect 14924 28756 14976 28762
rect 14924 28698 14976 28704
rect 15120 28558 15148 30602
rect 15200 29504 15252 29510
rect 15200 29446 15252 29452
rect 15212 29306 15240 29446
rect 15200 29300 15252 29306
rect 15200 29242 15252 29248
rect 15292 28960 15344 28966
rect 15292 28902 15344 28908
rect 15108 28552 15160 28558
rect 15108 28494 15160 28500
rect 14832 28416 14884 28422
rect 14832 28358 14884 28364
rect 14844 27470 14872 28358
rect 15120 27674 15148 28494
rect 15108 27668 15160 27674
rect 15108 27610 15160 27616
rect 15108 27532 15160 27538
rect 15108 27474 15160 27480
rect 14832 27464 14884 27470
rect 14832 27406 14884 27412
rect 14832 26988 14884 26994
rect 14832 26930 14884 26936
rect 14844 26314 14872 26930
rect 14924 26784 14976 26790
rect 14924 26726 14976 26732
rect 14832 26308 14884 26314
rect 14832 26250 14884 26256
rect 14648 26036 14700 26042
rect 14648 25978 14700 25984
rect 14844 25786 14872 26250
rect 14752 25758 14872 25786
rect 14556 25356 14608 25362
rect 14556 25298 14608 25304
rect 14648 25356 14700 25362
rect 14648 25298 14700 25304
rect 14568 24750 14596 25298
rect 14660 24886 14688 25298
rect 14648 24880 14700 24886
rect 14648 24822 14700 24828
rect 14556 24744 14608 24750
rect 14556 24686 14608 24692
rect 14188 23860 14240 23866
rect 14188 23802 14240 23808
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 13912 23656 13964 23662
rect 13912 23598 13964 23604
rect 13912 22636 13964 22642
rect 13912 22578 13964 22584
rect 13360 22568 13412 22574
rect 13360 22510 13412 22516
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12808 22160 12860 22166
rect 12808 22102 12860 22108
rect 12636 21542 12756 21570
rect 12532 21344 12584 21350
rect 12532 21286 12584 21292
rect 12440 20868 12492 20874
rect 12440 20810 12492 20816
rect 12452 19310 12480 20810
rect 12636 20602 12664 21542
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12624 20596 12676 20602
rect 12624 20538 12676 20544
rect 12728 20398 12756 21422
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 13372 21078 13400 22510
rect 13924 22234 13952 22578
rect 13912 22228 13964 22234
rect 13912 22170 13964 22176
rect 13360 21072 13412 21078
rect 13360 21014 13412 21020
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12728 19854 12756 20334
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12728 19666 12756 19790
rect 12728 19638 12848 19666
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12820 19174 12848 19638
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12348 18692 12400 18698
rect 12348 18634 12400 18640
rect 12360 18426 12388 18634
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 12452 17338 12480 18226
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12256 16040 12308 16046
rect 12256 15982 12308 15988
rect 12072 15972 12124 15978
rect 12072 15914 12124 15920
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 12268 15570 12296 15982
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12452 15366 12480 16050
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11796 13456 11848 13462
rect 11796 13398 11848 13404
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11716 9586 11744 13330
rect 11808 12986 11836 13398
rect 11900 12986 11928 14418
rect 11992 13258 12020 14826
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 12256 14476 12308 14482
rect 12256 14418 12308 14424
rect 12268 14074 12296 14418
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12360 14006 12388 14758
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12360 13818 12388 13942
rect 11980 13252 12032 13258
rect 11980 13194 12032 13200
rect 11992 12986 12020 13194
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 12164 13184 12216 13190
rect 12164 13126 12216 13132
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11808 12850 11836 12922
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11808 12753 11836 12786
rect 11794 12744 11850 12753
rect 11900 12714 11928 12922
rect 11794 12679 11850 12688
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11992 12434 12020 12922
rect 11900 12406 12020 12434
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11716 9042 11744 9522
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11518 8392 11574 8401
rect 11440 7886 11468 8366
rect 11518 8327 11574 8336
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11532 7562 11560 8327
rect 11440 7534 11560 7562
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 11256 1834 11284 4626
rect 11348 3194 11376 5782
rect 11440 5234 11468 7534
rect 11520 7472 11572 7478
rect 11520 7414 11572 7420
rect 11532 6730 11560 7414
rect 11716 6866 11744 8978
rect 11808 8090 11836 11494
rect 11900 10470 11928 12406
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11992 10130 12020 12242
rect 12084 10266 12112 13126
rect 12176 11218 12204 13126
rect 12268 12986 12296 13806
rect 12360 13790 12480 13818
rect 12452 13326 12480 13790
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12268 11082 12296 12922
rect 12452 12458 12480 12922
rect 12360 12430 12480 12458
rect 12544 12442 12572 15370
rect 12636 14618 12664 18566
rect 12820 18222 12848 19110
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12808 18216 12860 18222
rect 12808 18158 12860 18164
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12728 16182 12756 17070
rect 12820 16658 12848 18158
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 13372 17746 13400 21014
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13464 19122 13492 20334
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13556 19310 13584 20198
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13464 19094 13584 19122
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 13188 17270 13216 17478
rect 13176 17264 13228 17270
rect 13176 17206 13228 17212
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12716 16176 12768 16182
rect 12716 16118 12768 16124
rect 12728 15638 12756 16118
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12636 12918 12664 13670
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12622 12744 12678 12753
rect 12622 12679 12678 12688
rect 12532 12436 12584 12442
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 12360 10810 12388 12430
rect 12532 12378 12584 12384
rect 12440 12368 12492 12374
rect 12440 12310 12492 12316
rect 12452 12102 12480 12310
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12452 10996 12480 11630
rect 12544 11150 12572 12106
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12452 10968 12572 10996
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12544 10577 12572 10968
rect 12530 10568 12586 10577
rect 12256 10532 12308 10538
rect 12530 10503 12586 10512
rect 12256 10474 12308 10480
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 12162 10024 12218 10033
rect 12162 9959 12218 9968
rect 11888 9920 11940 9926
rect 11886 9888 11888 9897
rect 11940 9888 11942 9897
rect 11886 9823 11942 9832
rect 11900 9178 11928 9823
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11900 6914 11928 8978
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11992 7954 12020 8230
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11992 7546 12020 7890
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 11900 6886 12020 6914
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11532 5302 11560 6666
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11624 5370 11652 5646
rect 11612 5364 11664 5370
rect 11612 5306 11664 5312
rect 11716 5302 11744 6802
rect 11520 5296 11572 5302
rect 11520 5238 11572 5244
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 11900 4826 11928 5102
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11440 3074 11468 4762
rect 11704 4004 11756 4010
rect 11704 3946 11756 3952
rect 11348 3046 11468 3074
rect 11348 2038 11376 3046
rect 11716 2990 11744 3946
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11336 2032 11388 2038
rect 11336 1974 11388 1980
rect 11244 1828 11296 1834
rect 11244 1770 11296 1776
rect 11440 800 11468 2926
rect 11808 800 11836 2994
rect 11992 2378 12020 6886
rect 12084 5166 12112 7414
rect 12176 5778 12204 9959
rect 12268 9654 12296 10474
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12544 9994 12572 10134
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 12360 9518 12388 9930
rect 12440 9648 12492 9654
rect 12492 9608 12572 9636
rect 12440 9590 12492 9596
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12348 9376 12400 9382
rect 12348 9318 12400 9324
rect 12360 7002 12388 9318
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12452 6662 12480 8910
rect 12544 8566 12572 9608
rect 12636 8634 12664 12679
rect 12728 11898 12756 14214
rect 12820 13802 12848 14758
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13096 14074 13124 14350
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13372 13410 13400 15438
rect 13280 13382 13400 13410
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12820 12238 12848 12786
rect 13004 12646 13032 13262
rect 13280 13172 13308 13382
rect 13360 13320 13412 13326
rect 13464 13308 13492 18566
rect 13556 17134 13584 19094
rect 13544 17128 13596 17134
rect 13544 17070 13596 17076
rect 13648 17066 13676 20538
rect 14016 20058 14044 23666
rect 14188 23112 14240 23118
rect 14188 23054 14240 23060
rect 14096 23044 14148 23050
rect 14096 22986 14148 22992
rect 14108 22778 14136 22986
rect 14200 22778 14228 23054
rect 14752 22778 14780 25758
rect 14832 25696 14884 25702
rect 14832 25638 14884 25644
rect 14844 25362 14872 25638
rect 14832 25356 14884 25362
rect 14832 25298 14884 25304
rect 14844 24954 14872 25298
rect 14832 24948 14884 24954
rect 14832 24890 14884 24896
rect 14936 23866 14964 26726
rect 15016 26444 15068 26450
rect 15016 26386 15068 26392
rect 15028 25702 15056 26386
rect 15120 26382 15148 27474
rect 15200 27124 15252 27130
rect 15200 27066 15252 27072
rect 15212 26450 15240 27066
rect 15200 26444 15252 26450
rect 15200 26386 15252 26392
rect 15108 26376 15160 26382
rect 15108 26318 15160 26324
rect 15016 25696 15068 25702
rect 15016 25638 15068 25644
rect 15200 25288 15252 25294
rect 15200 25230 15252 25236
rect 15016 24744 15068 24750
rect 15016 24686 15068 24692
rect 14924 23860 14976 23866
rect 14924 23802 14976 23808
rect 14096 22772 14148 22778
rect 14096 22714 14148 22720
rect 14188 22772 14240 22778
rect 14188 22714 14240 22720
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 14096 22432 14148 22438
rect 14096 22374 14148 22380
rect 14108 22030 14136 22374
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 14108 21486 14136 21966
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14844 21554 14872 21830
rect 14832 21548 14884 21554
rect 14832 21490 14884 21496
rect 14096 21480 14148 21486
rect 14096 21422 14148 21428
rect 14556 21412 14608 21418
rect 14556 21354 14608 21360
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 14384 20398 14412 21286
rect 14372 20392 14424 20398
rect 14372 20334 14424 20340
rect 14004 20052 14056 20058
rect 14004 19994 14056 20000
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 14280 18624 14332 18630
rect 14280 18566 14332 18572
rect 13832 18426 13860 18566
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13832 17814 13860 18362
rect 14188 18216 14240 18222
rect 13910 18184 13966 18193
rect 13910 18119 13966 18128
rect 14186 18184 14188 18193
rect 14240 18184 14242 18193
rect 14186 18119 14242 18128
rect 13820 17808 13872 17814
rect 13820 17750 13872 17756
rect 13728 17604 13780 17610
rect 13728 17546 13780 17552
rect 13740 17338 13768 17546
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13832 16726 13860 16934
rect 13820 16720 13872 16726
rect 13820 16662 13872 16668
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13556 16454 13584 16594
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13556 13530 13584 16390
rect 13648 14890 13676 16526
rect 13636 14884 13688 14890
rect 13636 14826 13688 14832
rect 13924 14362 13952 18119
rect 14292 17678 14320 18566
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14384 16522 14412 19110
rect 14372 16516 14424 16522
rect 14372 16458 14424 16464
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14292 16114 14320 16390
rect 14384 16182 14412 16458
rect 14372 16176 14424 16182
rect 14372 16118 14424 16124
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14292 15978 14320 16050
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14280 15972 14332 15978
rect 14280 15914 14332 15920
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13740 14334 13952 14362
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13412 13280 13492 13308
rect 13360 13262 13412 13268
rect 13280 13144 13400 13172
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 13096 12753 13124 12854
rect 13082 12744 13138 12753
rect 13082 12679 13138 12688
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 13280 11778 13308 12038
rect 13372 11898 13400 13144
rect 13452 12912 13504 12918
rect 13452 12854 13504 12860
rect 13464 12238 13492 12854
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13450 11928 13506 11937
rect 13360 11892 13412 11898
rect 13450 11863 13452 11872
rect 13360 11834 13412 11840
rect 13504 11863 13506 11872
rect 13452 11834 13504 11840
rect 13280 11750 13400 11778
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 13372 11286 13400 11750
rect 13556 11370 13584 12582
rect 13464 11342 13584 11370
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 12900 11280 12952 11286
rect 13084 11280 13136 11286
rect 12952 11228 13084 11234
rect 12900 11222 13136 11228
rect 13360 11280 13412 11286
rect 13360 11222 13412 11228
rect 12714 10840 12770 10849
rect 12714 10775 12716 10784
rect 12768 10775 12770 10784
rect 12716 10746 12768 10752
rect 12820 10674 12848 11222
rect 12912 11206 13124 11222
rect 12900 11144 12952 11150
rect 12952 11104 13400 11132
rect 12900 11086 12952 11092
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 12728 10062 12756 10542
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12808 9920 12860 9926
rect 12714 9888 12770 9897
rect 12808 9862 12860 9868
rect 12714 9823 12770 9832
rect 12728 9722 12756 9823
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12820 9178 12848 9862
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 13372 9110 13400 11104
rect 13464 10742 13492 11342
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13452 10736 13504 10742
rect 13452 10678 13504 10684
rect 13450 10160 13506 10169
rect 13556 10130 13584 11154
rect 13648 10538 13676 14282
rect 13740 12306 13768 14334
rect 13912 14272 13964 14278
rect 13910 14240 13912 14249
rect 13964 14240 13966 14249
rect 13910 14175 13966 14184
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13832 13394 13860 13806
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13740 11694 13768 12242
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 13636 10532 13688 10538
rect 13636 10474 13688 10480
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13450 10095 13506 10104
rect 13544 10124 13596 10130
rect 13360 9104 13412 9110
rect 13360 9046 13412 9052
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 13360 8424 13412 8430
rect 13360 8366 13412 8372
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12636 7546 12664 7686
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12530 7440 12586 7449
rect 12530 7375 12586 7384
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12268 5914 12296 6190
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12164 5772 12216 5778
rect 12164 5714 12216 5720
rect 12544 5710 12572 7375
rect 12820 6458 12848 8298
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 13372 7886 13400 8366
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12268 4049 12296 4082
rect 12624 4072 12676 4078
rect 12254 4040 12310 4049
rect 12624 4014 12676 4020
rect 12254 3975 12310 3984
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12176 2446 12204 3878
rect 12636 3754 12664 4014
rect 12452 3726 12664 3754
rect 12452 2446 12480 3726
rect 12636 3641 12664 3726
rect 12622 3632 12678 3641
rect 12532 3596 12584 3602
rect 12622 3567 12678 3576
rect 12532 3538 12584 3544
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 11980 2372 12032 2378
rect 11980 2314 12032 2320
rect 12176 800 12204 2382
rect 12544 800 12572 3538
rect 12728 1902 12756 6258
rect 13372 6186 13400 7686
rect 13464 7206 13492 10095
rect 13544 10066 13596 10072
rect 13556 9042 13584 10066
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13648 7698 13676 10202
rect 13740 9382 13768 11018
rect 13832 9450 13860 12718
rect 13924 12442 13952 13126
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 14016 11898 14044 15846
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 14108 12782 14136 13670
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14200 12374 14228 15302
rect 14292 15162 14320 15302
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14384 14521 14412 15982
rect 14370 14512 14426 14521
rect 14370 14447 14426 14456
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 14188 12368 14240 12374
rect 14188 12310 14240 12316
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 14004 11892 14056 11898
rect 14004 11834 14056 11840
rect 13924 10266 13952 11834
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 14016 11286 14044 11698
rect 14004 11280 14056 11286
rect 14004 11222 14056 11228
rect 14004 11076 14056 11082
rect 14004 11018 14056 11024
rect 14016 10713 14044 11018
rect 14002 10704 14058 10713
rect 14002 10639 14058 10648
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13728 9376 13780 9382
rect 14016 9330 14044 10542
rect 14108 10266 14136 12310
rect 14292 11914 14320 14214
rect 14384 13326 14412 14447
rect 14568 13462 14596 21354
rect 15028 21350 15056 24686
rect 15212 24682 15240 25230
rect 15304 25106 15332 28902
rect 15384 28620 15436 28626
rect 15384 28562 15436 28568
rect 15396 27946 15424 28562
rect 15580 28218 15608 42026
rect 15764 35494 15792 46446
rect 16488 46028 16540 46034
rect 16488 45970 16540 45976
rect 16212 41744 16264 41750
rect 16212 41686 16264 41692
rect 15752 35488 15804 35494
rect 15752 35430 15804 35436
rect 16120 32972 16172 32978
rect 16120 32914 16172 32920
rect 16132 31890 16160 32914
rect 16120 31884 16172 31890
rect 16120 31826 16172 31832
rect 16132 31278 16160 31826
rect 16120 31272 16172 31278
rect 16120 31214 16172 31220
rect 16028 30184 16080 30190
rect 16028 30126 16080 30132
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 15660 29640 15712 29646
rect 15660 29582 15712 29588
rect 15568 28212 15620 28218
rect 15568 28154 15620 28160
rect 15384 27940 15436 27946
rect 15384 27882 15436 27888
rect 15476 27328 15528 27334
rect 15476 27270 15528 27276
rect 15384 25832 15436 25838
rect 15384 25774 15436 25780
rect 15396 25226 15424 25774
rect 15384 25220 15436 25226
rect 15384 25162 15436 25168
rect 15304 25078 15424 25106
rect 15200 24676 15252 24682
rect 15200 24618 15252 24624
rect 15108 24608 15160 24614
rect 15108 24550 15160 24556
rect 15120 24410 15148 24550
rect 15108 24404 15160 24410
rect 15108 24346 15160 24352
rect 15200 23316 15252 23322
rect 15200 23258 15252 23264
rect 15108 22704 15160 22710
rect 15108 22646 15160 22652
rect 15120 21622 15148 22646
rect 15212 22506 15240 23258
rect 15200 22500 15252 22506
rect 15200 22442 15252 22448
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 15108 21616 15160 21622
rect 15108 21558 15160 21564
rect 15120 21350 15148 21558
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 15108 21344 15160 21350
rect 15108 21286 15160 21292
rect 14648 20868 14700 20874
rect 14648 20810 14700 20816
rect 14660 20466 14688 20810
rect 15120 20806 15148 21286
rect 15108 20800 15160 20806
rect 15108 20742 15160 20748
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14660 19786 14688 20402
rect 15108 20324 15160 20330
rect 15108 20266 15160 20272
rect 14648 19780 14700 19786
rect 14648 19722 14700 19728
rect 14660 19174 14688 19722
rect 14832 19236 14884 19242
rect 14832 19178 14884 19184
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14660 16794 14688 19110
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 14752 15366 14780 16050
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14660 14278 14688 14554
rect 14752 14346 14780 15302
rect 14740 14340 14792 14346
rect 14740 14282 14792 14288
rect 14648 14272 14700 14278
rect 14648 14214 14700 14220
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14556 13456 14608 13462
rect 14556 13398 14608 13404
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14384 12646 14412 12922
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14568 12424 14596 13262
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14660 12889 14688 13126
rect 14646 12880 14702 12889
rect 14646 12815 14702 12824
rect 14752 12434 14780 13466
rect 14476 12396 14596 12424
rect 14660 12406 14780 12434
rect 14370 12064 14426 12073
rect 14370 11999 14426 12008
rect 14200 11886 14320 11914
rect 14200 11830 14228 11886
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14188 11280 14240 11286
rect 14188 11222 14240 11228
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 13728 9318 13780 9324
rect 13832 9302 14044 9330
rect 13728 8560 13780 8566
rect 13832 8537 13860 9302
rect 14108 9194 14136 9454
rect 13924 9166 14136 9194
rect 13728 8502 13780 8508
rect 13818 8528 13874 8537
rect 13740 7886 13768 8502
rect 13818 8463 13874 8472
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13556 7670 13676 7698
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13556 6882 13584 7670
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13464 6854 13584 6882
rect 13360 6180 13412 6186
rect 13360 6122 13412 6128
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 13464 5642 13492 6854
rect 13542 6760 13598 6769
rect 13542 6695 13598 6704
rect 13556 6662 13584 6695
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13648 6254 13676 7482
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13452 5636 13504 5642
rect 13452 5578 13504 5584
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 13464 4570 13492 5578
rect 13648 5370 13676 6190
rect 13740 6186 13768 6734
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13372 4542 13492 4570
rect 13372 4146 13400 4542
rect 13452 4480 13504 4486
rect 13452 4422 13504 4428
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12716 1896 12768 1902
rect 12716 1838 12768 1844
rect 12820 1714 12848 3538
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13464 2582 13492 4422
rect 13832 3738 13860 8463
rect 13924 5794 13952 9166
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 14016 7750 14044 7890
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 14016 5914 14044 6326
rect 14004 5908 14056 5914
rect 14004 5850 14056 5856
rect 13924 5766 14044 5794
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 13924 4146 13952 4966
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14016 4026 14044 5766
rect 13924 3998 14044 4026
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 13924 3194 13952 3998
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13452 2576 13504 2582
rect 13452 2518 13504 2524
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12820 1686 12940 1714
rect 12912 800 12940 1686
rect 13280 800 13308 2314
rect 13648 800 13676 2926
rect 14016 800 14044 3538
rect 14108 3058 14136 8502
rect 14200 6866 14228 11222
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14292 10849 14320 10950
rect 14278 10840 14334 10849
rect 14278 10775 14334 10784
rect 14278 9072 14334 9081
rect 14278 9007 14334 9016
rect 14292 7478 14320 9007
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 14188 6860 14240 6866
rect 14188 6802 14240 6808
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14186 6352 14242 6361
rect 14186 6287 14188 6296
rect 14240 6287 14242 6296
rect 14188 6258 14240 6264
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14200 4214 14228 5306
rect 14292 4622 14320 6598
rect 14384 5914 14412 11999
rect 14476 10606 14504 12396
rect 14660 12238 14688 12406
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14464 10600 14516 10606
rect 14462 10568 14464 10577
rect 14516 10568 14518 10577
rect 14462 10503 14518 10512
rect 14556 10056 14608 10062
rect 14556 9998 14608 10004
rect 14568 9722 14596 9998
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14568 9518 14596 9658
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14568 9042 14596 9454
rect 14660 9450 14688 12174
rect 14844 12050 14872 19178
rect 15120 19174 15148 20266
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 15212 17882 15240 21830
rect 15396 21622 15424 25078
rect 15384 21616 15436 21622
rect 15384 21558 15436 21564
rect 15488 20777 15516 27270
rect 15580 26314 15608 28154
rect 15568 26308 15620 26314
rect 15568 26250 15620 26256
rect 15672 25158 15700 29582
rect 15948 29238 15976 29990
rect 16040 29714 16068 30126
rect 16028 29708 16080 29714
rect 16028 29650 16080 29656
rect 16120 29504 16172 29510
rect 16120 29446 16172 29452
rect 15936 29232 15988 29238
rect 15936 29174 15988 29180
rect 15752 29028 15804 29034
rect 16132 28994 16160 29446
rect 15752 28970 15804 28976
rect 15764 27062 15792 28970
rect 15948 28966 16160 28994
rect 15752 27056 15804 27062
rect 15752 26998 15804 27004
rect 15660 25152 15712 25158
rect 15660 25094 15712 25100
rect 15752 25152 15804 25158
rect 15752 25094 15804 25100
rect 15672 24954 15700 25094
rect 15660 24948 15712 24954
rect 15660 24890 15712 24896
rect 15672 24857 15700 24890
rect 15658 24848 15714 24857
rect 15658 24783 15714 24792
rect 15568 24608 15620 24614
rect 15568 24550 15620 24556
rect 15474 20768 15530 20777
rect 15474 20703 15530 20712
rect 15580 20602 15608 24550
rect 15660 23656 15712 23662
rect 15660 23598 15712 23604
rect 15672 23118 15700 23598
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15764 22166 15792 25094
rect 15948 24886 15976 28966
rect 16028 28416 16080 28422
rect 16028 28358 16080 28364
rect 16040 27402 16068 28358
rect 16224 28098 16252 41686
rect 16304 37324 16356 37330
rect 16304 37266 16356 37272
rect 16316 28490 16344 37266
rect 16500 34950 16528 45970
rect 16960 45554 16988 53926
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 18696 52964 18748 52970
rect 18696 52906 18748 52912
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 18604 50720 18656 50726
rect 18604 50662 18656 50668
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 17592 48068 17644 48074
rect 17592 48010 17644 48016
rect 16776 45526 16988 45554
rect 16580 43988 16632 43994
rect 16580 43930 16632 43936
rect 16488 34944 16540 34950
rect 16488 34886 16540 34892
rect 16592 32978 16620 43930
rect 16776 33114 16804 45526
rect 16856 44192 16908 44198
rect 16856 44134 16908 44140
rect 16764 33108 16816 33114
rect 16764 33050 16816 33056
rect 16580 32972 16632 32978
rect 16580 32914 16632 32920
rect 16776 32910 16804 33050
rect 16764 32904 16816 32910
rect 16764 32846 16816 32852
rect 16672 32496 16724 32502
rect 16672 32438 16724 32444
rect 16580 32224 16632 32230
rect 16580 32166 16632 32172
rect 16592 31822 16620 32166
rect 16580 31816 16632 31822
rect 16580 31758 16632 31764
rect 16592 31142 16620 31758
rect 16684 31686 16712 32438
rect 16764 32360 16816 32366
rect 16764 32302 16816 32308
rect 16776 31822 16804 32302
rect 16764 31816 16816 31822
rect 16764 31758 16816 31764
rect 16672 31680 16724 31686
rect 16672 31622 16724 31628
rect 16580 31136 16632 31142
rect 16580 31078 16632 31084
rect 16580 30388 16632 30394
rect 16580 30330 16632 30336
rect 16488 30116 16540 30122
rect 16488 30058 16540 30064
rect 16500 29782 16528 30058
rect 16488 29776 16540 29782
rect 16488 29718 16540 29724
rect 16500 29510 16528 29718
rect 16488 29504 16540 29510
rect 16488 29446 16540 29452
rect 16488 28688 16540 28694
rect 16488 28630 16540 28636
rect 16304 28484 16356 28490
rect 16304 28426 16356 28432
rect 16500 28422 16528 28630
rect 16488 28416 16540 28422
rect 16488 28358 16540 28364
rect 16224 28082 16344 28098
rect 16224 28076 16356 28082
rect 16224 28070 16304 28076
rect 16304 28018 16356 28024
rect 16316 27878 16344 28018
rect 16304 27872 16356 27878
rect 16304 27814 16356 27820
rect 16120 27600 16172 27606
rect 16120 27542 16172 27548
rect 16028 27396 16080 27402
rect 16028 27338 16080 27344
rect 16028 26580 16080 26586
rect 16028 26522 16080 26528
rect 16040 26314 16068 26522
rect 16028 26308 16080 26314
rect 16028 26250 16080 26256
rect 15936 24880 15988 24886
rect 15936 24822 15988 24828
rect 15844 23792 15896 23798
rect 15844 23734 15896 23740
rect 15752 22160 15804 22166
rect 15752 22102 15804 22108
rect 15752 20868 15804 20874
rect 15752 20810 15804 20816
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15764 20058 15792 20810
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15764 19310 15792 19994
rect 15856 19922 15884 23734
rect 15844 19916 15896 19922
rect 15896 19876 16068 19904
rect 15844 19858 15896 19864
rect 15844 19780 15896 19786
rect 15844 19722 15896 19728
rect 15752 19304 15804 19310
rect 15752 19246 15804 19252
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15488 16590 15516 17478
rect 15568 17128 15620 17134
rect 15568 17070 15620 17076
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 15028 16250 15056 16390
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 15028 15706 15056 15982
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15396 13394 15424 14418
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 14752 12022 14872 12050
rect 14752 11286 14780 12022
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 14740 11280 14792 11286
rect 14740 11222 14792 11228
rect 14844 10198 14872 11834
rect 14832 10192 14884 10198
rect 14832 10134 14884 10140
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14648 9444 14700 9450
rect 14648 9386 14700 9392
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 14568 8634 14596 8978
rect 14660 8838 14688 9114
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14648 8492 14700 8498
rect 14568 8452 14648 8480
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14476 7478 14504 7822
rect 14464 7472 14516 7478
rect 14464 7414 14516 7420
rect 14372 5908 14424 5914
rect 14372 5850 14424 5856
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14188 4208 14240 4214
rect 14188 4150 14240 4156
rect 14384 3670 14412 5850
rect 14476 5302 14504 7414
rect 14464 5296 14516 5302
rect 14464 5238 14516 5244
rect 14476 4842 14504 5238
rect 14568 4978 14596 8452
rect 14648 8434 14700 8440
rect 14646 7984 14702 7993
rect 14646 7919 14702 7928
rect 14660 7886 14688 7919
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14648 6928 14700 6934
rect 14648 6870 14700 6876
rect 14660 6730 14688 6870
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14568 4950 14688 4978
rect 14476 4814 14596 4842
rect 14568 4486 14596 4814
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14372 3664 14424 3670
rect 14372 3606 14424 3612
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14200 2774 14228 3130
rect 14108 2746 14228 2774
rect 14108 2446 14136 2746
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14384 800 14412 2450
rect 14476 2446 14504 4422
rect 14568 4282 14596 4422
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 14660 2961 14688 4950
rect 14752 4622 14780 9862
rect 14844 8838 14872 10134
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14832 7948 14884 7954
rect 14832 7890 14884 7896
rect 14844 7002 14872 7890
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 14936 5250 14964 13262
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 15028 12170 15056 12582
rect 15120 12434 15148 12786
rect 15120 12406 15240 12434
rect 15212 12374 15240 12406
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15016 11824 15068 11830
rect 15016 11766 15068 11772
rect 15028 10130 15056 11766
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 15120 9178 15148 11698
rect 15212 11082 15240 11834
rect 15304 11354 15332 13126
rect 15396 11762 15424 13126
rect 15488 12889 15516 14758
rect 15580 14074 15608 17070
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15672 16250 15700 16458
rect 15660 16244 15712 16250
rect 15660 16186 15712 16192
rect 15764 15450 15792 17614
rect 15856 16454 15884 19722
rect 16040 17218 16068 19876
rect 16132 19378 16160 27542
rect 16316 26314 16344 27814
rect 16500 27334 16528 28358
rect 16488 27328 16540 27334
rect 16488 27270 16540 27276
rect 16304 26308 16356 26314
rect 16304 26250 16356 26256
rect 16304 26036 16356 26042
rect 16304 25978 16356 25984
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 16040 17190 16160 17218
rect 16132 17134 16160 17190
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 15936 17060 15988 17066
rect 15936 17002 15988 17008
rect 16028 17060 16080 17066
rect 16028 17002 16080 17008
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15672 15422 15792 15450
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15474 12880 15530 12889
rect 15474 12815 15476 12824
rect 15528 12815 15530 12824
rect 15476 12786 15528 12792
rect 15580 12782 15608 13738
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15292 11076 15344 11082
rect 15396 11064 15424 11290
rect 15344 11036 15424 11064
rect 15292 11018 15344 11024
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 14844 5222 14964 5250
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14740 2984 14792 2990
rect 14646 2952 14702 2961
rect 14740 2926 14792 2932
rect 14646 2887 14702 2896
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 14752 800 14780 2926
rect 14844 2854 14872 5222
rect 14924 5092 14976 5098
rect 14924 5034 14976 5040
rect 14936 4690 14964 5034
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 14924 4548 14976 4554
rect 14924 4490 14976 4496
rect 14936 3738 14964 4490
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 15028 3466 15056 8774
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 15120 7993 15148 8434
rect 15106 7984 15162 7993
rect 15106 7919 15162 7928
rect 15212 7750 15240 11018
rect 15476 11008 15528 11014
rect 15476 10950 15528 10956
rect 15384 10736 15436 10742
rect 15384 10678 15436 10684
rect 15396 10538 15424 10678
rect 15384 10532 15436 10538
rect 15384 10474 15436 10480
rect 15488 9926 15516 10950
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15580 9738 15608 12038
rect 15672 11937 15700 15422
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15764 15162 15792 15302
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15948 15026 15976 17002
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15658 11928 15714 11937
rect 15658 11863 15714 11872
rect 15672 11762 15700 11863
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15672 9994 15700 10202
rect 15660 9988 15712 9994
rect 15660 9930 15712 9936
rect 15396 9710 15608 9738
rect 15396 9586 15424 9710
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15304 7818 15332 9114
rect 15396 8838 15424 9522
rect 15764 9518 15792 13330
rect 15856 13190 15884 14758
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15934 12744 15990 12753
rect 15856 12306 15884 12718
rect 15934 12679 15990 12688
rect 15844 12300 15896 12306
rect 15844 12242 15896 12248
rect 15856 10130 15884 12242
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15844 9920 15896 9926
rect 15844 9862 15896 9868
rect 15856 9722 15884 9862
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 15568 9512 15620 9518
rect 15568 9454 15620 9460
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15580 9110 15608 9454
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15568 9104 15620 9110
rect 15568 9046 15620 9052
rect 15672 8838 15700 9318
rect 15764 9110 15792 9454
rect 15752 9104 15804 9110
rect 15752 9046 15804 9052
rect 15856 9058 15884 9658
rect 15948 9382 15976 12679
rect 16040 12102 16068 17002
rect 16224 16538 16252 19314
rect 16316 17814 16344 25978
rect 16500 25498 16528 27270
rect 16592 26994 16620 30330
rect 16684 28082 16712 31622
rect 16776 31346 16804 31758
rect 16764 31340 16816 31346
rect 16764 31282 16816 31288
rect 16764 31136 16816 31142
rect 16764 31078 16816 31084
rect 16672 28076 16724 28082
rect 16672 28018 16724 28024
rect 16776 28014 16804 31078
rect 16868 30258 16896 44134
rect 17132 32904 17184 32910
rect 17132 32846 17184 32852
rect 17040 32768 17092 32774
rect 17040 32710 17092 32716
rect 17052 32570 17080 32710
rect 17040 32564 17092 32570
rect 17040 32506 17092 32512
rect 17144 31754 17172 32846
rect 17052 31726 17172 31754
rect 16856 30252 16908 30258
rect 16856 30194 16908 30200
rect 16868 28994 16896 30194
rect 17052 29238 17080 31726
rect 17604 31226 17632 48010
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 18616 37330 18644 50662
rect 18708 41750 18736 52906
rect 20076 49088 20128 49094
rect 20076 49030 20128 49036
rect 19984 44804 20036 44810
rect 19984 44746 20036 44752
rect 19524 43784 19576 43790
rect 19524 43726 19576 43732
rect 18696 41744 18748 41750
rect 18696 41686 18748 41692
rect 18604 37324 18656 37330
rect 18604 37266 18656 37272
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 19536 34082 19564 43726
rect 19996 35018 20024 44746
rect 19984 35012 20036 35018
rect 19984 34954 20036 34960
rect 20088 34218 20116 49030
rect 19904 34190 20116 34218
rect 19536 34066 19748 34082
rect 19536 34060 19760 34066
rect 19536 34054 19708 34060
rect 19432 33992 19484 33998
rect 19432 33934 19484 33940
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 17868 32972 17920 32978
rect 17868 32914 17920 32920
rect 17684 31884 17736 31890
rect 17684 31826 17736 31832
rect 17696 31278 17724 31826
rect 17144 31198 17632 31226
rect 17684 31272 17736 31278
rect 17684 31214 17736 31220
rect 17040 29232 17092 29238
rect 17040 29174 17092 29180
rect 16868 28966 16988 28994
rect 16764 28008 16816 28014
rect 16764 27950 16816 27956
rect 16856 27872 16908 27878
rect 16856 27814 16908 27820
rect 16868 27130 16896 27814
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 16580 26988 16632 26994
rect 16580 26930 16632 26936
rect 16592 26450 16620 26930
rect 16580 26444 16632 26450
rect 16580 26386 16632 26392
rect 16488 25492 16540 25498
rect 16488 25434 16540 25440
rect 16396 25220 16448 25226
rect 16396 25162 16448 25168
rect 16408 24954 16436 25162
rect 16500 25158 16528 25434
rect 16488 25152 16540 25158
rect 16488 25094 16540 25100
rect 16396 24948 16448 24954
rect 16396 24890 16448 24896
rect 16592 24070 16620 26386
rect 16960 26382 16988 28966
rect 17040 26580 17092 26586
rect 17040 26522 17092 26528
rect 16948 26376 17000 26382
rect 16948 26318 17000 26324
rect 16856 25696 16908 25702
rect 16856 25638 16908 25644
rect 16868 25362 16896 25638
rect 16856 25356 16908 25362
rect 16856 25298 16908 25304
rect 17052 24886 17080 26522
rect 17040 24880 17092 24886
rect 17040 24822 17092 24828
rect 17040 24676 17092 24682
rect 17040 24618 17092 24624
rect 16580 24064 16632 24070
rect 16580 24006 16632 24012
rect 16592 23866 16620 24006
rect 16580 23860 16632 23866
rect 16580 23802 16632 23808
rect 16856 23044 16908 23050
rect 16856 22986 16908 22992
rect 16868 22778 16896 22986
rect 16856 22772 16908 22778
rect 16856 22714 16908 22720
rect 16948 22092 17000 22098
rect 16948 22034 17000 22040
rect 16960 21962 16988 22034
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16948 21956 17000 21962
rect 16948 21898 17000 21904
rect 16500 20806 16528 21898
rect 16580 21888 16632 21894
rect 16580 21830 16632 21836
rect 16592 21078 16620 21830
rect 16580 21072 16632 21078
rect 16580 21014 16632 21020
rect 16488 20800 16540 20806
rect 16488 20742 16540 20748
rect 16304 17808 16356 17814
rect 16304 17750 16356 17756
rect 16396 17332 16448 17338
rect 16396 17274 16448 17280
rect 16408 16658 16436 17274
rect 16500 16726 16528 20742
rect 16592 18290 16620 21014
rect 16960 20890 16988 21898
rect 17052 21894 17080 24618
rect 17144 23322 17172 31198
rect 17500 31136 17552 31142
rect 17500 31078 17552 31084
rect 17512 30818 17540 31078
rect 17512 30790 17632 30818
rect 17500 29300 17552 29306
rect 17500 29242 17552 29248
rect 17408 29164 17460 29170
rect 17408 29106 17460 29112
rect 17420 28014 17448 29106
rect 17408 28008 17460 28014
rect 17408 27950 17460 27956
rect 17408 26444 17460 26450
rect 17408 26386 17460 26392
rect 17224 26376 17276 26382
rect 17224 26318 17276 26324
rect 17132 23316 17184 23322
rect 17132 23258 17184 23264
rect 17144 23225 17172 23258
rect 17130 23216 17186 23225
rect 17130 23151 17186 23160
rect 17040 21888 17092 21894
rect 17040 21830 17092 21836
rect 17132 21888 17184 21894
rect 17132 21830 17184 21836
rect 16960 20862 17080 20890
rect 17052 20806 17080 20862
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16684 18902 16712 19790
rect 17052 19718 17080 20742
rect 17144 20534 17172 21830
rect 17132 20528 17184 20534
rect 17132 20470 17184 20476
rect 17144 19990 17172 20470
rect 17132 19984 17184 19990
rect 17132 19926 17184 19932
rect 17040 19712 17092 19718
rect 17040 19654 17092 19660
rect 16672 18896 16724 18902
rect 16672 18838 16724 18844
rect 16670 18728 16726 18737
rect 16670 18663 16726 18672
rect 16684 18426 16712 18663
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16592 17338 16620 18226
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16684 17218 16712 18158
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16856 17604 16908 17610
rect 16856 17546 16908 17552
rect 16592 17190 16712 17218
rect 16488 16720 16540 16726
rect 16488 16662 16540 16668
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16132 16510 16252 16538
rect 16132 15094 16160 16510
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 16224 16250 16252 16390
rect 16212 16244 16264 16250
rect 16212 16186 16264 16192
rect 16120 15088 16172 15094
rect 16120 15030 16172 15036
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 16028 12096 16080 12102
rect 16132 12073 16160 14350
rect 16224 13326 16252 16186
rect 16408 15570 16436 16594
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16396 15428 16448 15434
rect 16396 15370 16448 15376
rect 16408 13852 16436 15370
rect 16592 14958 16620 17190
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16500 14074 16528 14214
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16488 13864 16540 13870
rect 16408 13824 16488 13852
rect 16488 13806 16540 13812
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 16500 12288 16528 13806
rect 16578 13696 16634 13705
rect 16578 13631 16634 13640
rect 16224 12260 16528 12288
rect 16028 12038 16080 12044
rect 16118 12064 16174 12073
rect 16118 11999 16174 12008
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16026 11112 16082 11121
rect 16026 11047 16082 11056
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15292 7812 15344 7818
rect 15292 7754 15344 7760
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15120 5710 15148 7142
rect 15396 6361 15424 8774
rect 15764 7954 15792 9046
rect 15856 9030 15976 9058
rect 15948 8974 15976 9030
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15856 8090 15884 8910
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15844 7812 15896 7818
rect 15844 7754 15896 7760
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15382 6352 15438 6361
rect 15382 6287 15438 6296
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 15212 5817 15240 6054
rect 15198 5808 15254 5817
rect 15198 5743 15200 5752
rect 15252 5743 15254 5752
rect 15384 5772 15436 5778
rect 15200 5714 15252 5720
rect 15384 5714 15436 5720
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 15120 4690 15148 5646
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15016 3460 15068 3466
rect 15016 3402 15068 3408
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 14832 2848 14884 2854
rect 14832 2790 14884 2796
rect 15120 800 15148 2858
rect 15212 2106 15240 5102
rect 15396 4554 15424 5714
rect 15488 5030 15516 6734
rect 15672 6118 15700 7686
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15476 4684 15528 4690
rect 15476 4626 15528 4632
rect 15488 4570 15516 4626
rect 15384 4548 15436 4554
rect 15488 4542 15608 4570
rect 15384 4490 15436 4496
rect 15396 4298 15424 4490
rect 15396 4282 15516 4298
rect 15396 4276 15528 4282
rect 15396 4270 15476 4276
rect 15476 4218 15528 4224
rect 15580 4214 15608 4542
rect 15568 4208 15620 4214
rect 15568 4150 15620 4156
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15200 2100 15252 2106
rect 15200 2042 15252 2048
rect 15488 800 15516 3538
rect 15672 2310 15700 6054
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15764 2650 15792 5102
rect 15856 4690 15884 7754
rect 15948 5846 15976 8910
rect 15936 5840 15988 5846
rect 15936 5782 15988 5788
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 15844 4548 15896 4554
rect 15844 4490 15896 4496
rect 15856 3346 15884 4490
rect 16040 3534 16068 11047
rect 16132 8090 16160 11698
rect 16224 11150 16252 12260
rect 16592 12050 16620 13631
rect 16316 12022 16620 12050
rect 16316 11354 16344 12022
rect 16684 11914 16712 16934
rect 16868 16522 16896 17546
rect 16960 17377 16988 17614
rect 16946 17368 17002 17377
rect 16946 17303 17002 17312
rect 16960 17270 16988 17303
rect 16948 17264 17000 17270
rect 16948 17206 17000 17212
rect 16948 17128 17000 17134
rect 16948 17070 17000 17076
rect 16960 16726 16988 17070
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 16856 16516 16908 16522
rect 16856 16458 16908 16464
rect 16868 16250 16896 16458
rect 16856 16244 16908 16250
rect 16856 16186 16908 16192
rect 16960 15434 16988 16662
rect 16948 15428 17000 15434
rect 16948 15370 17000 15376
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16408 11886 16712 11914
rect 16776 11898 16804 15302
rect 16856 14544 16908 14550
rect 16908 14504 16988 14532
rect 16856 14486 16908 14492
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16868 12434 16896 13806
rect 16960 12986 16988 14504
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 16868 12406 16988 12434
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16764 11892 16816 11898
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16316 7478 16344 11290
rect 16408 8922 16436 11886
rect 16764 11834 16816 11840
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16488 10600 16540 10606
rect 16486 10568 16488 10577
rect 16540 10568 16542 10577
rect 16486 10503 16542 10512
rect 16500 9042 16528 10503
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16408 8894 16528 8922
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16304 7472 16356 7478
rect 16304 7414 16356 7420
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 15856 3318 16068 3346
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 15660 2304 15712 2310
rect 15660 2246 15712 2252
rect 15856 800 15884 2926
rect 16040 2650 16068 3318
rect 16028 2644 16080 2650
rect 16028 2586 16080 2592
rect 16040 2514 16068 2586
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 16132 2446 16160 6190
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16224 800 16252 4014
rect 16408 3398 16436 8026
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16500 3194 16528 8894
rect 16592 7886 16620 11698
rect 16672 11688 16724 11694
rect 16672 11630 16724 11636
rect 16684 11286 16712 11630
rect 16672 11280 16724 11286
rect 16672 11222 16724 11228
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16684 7342 16712 11222
rect 16868 10674 16896 12242
rect 16960 12170 16988 12406
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16960 11218 16988 12106
rect 17052 11898 17080 18566
rect 17144 15706 17172 18566
rect 17236 17814 17264 26318
rect 17316 23520 17368 23526
rect 17316 23462 17368 23468
rect 17328 19514 17356 23462
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17316 18760 17368 18766
rect 17420 18748 17448 26386
rect 17512 20346 17540 29242
rect 17604 27334 17632 30790
rect 17696 29458 17724 31214
rect 17696 29430 17816 29458
rect 17684 27940 17736 27946
rect 17684 27882 17736 27888
rect 17592 27328 17644 27334
rect 17592 27270 17644 27276
rect 17592 26580 17644 26586
rect 17592 26522 17644 26528
rect 17604 25974 17632 26522
rect 17592 25968 17644 25974
rect 17592 25910 17644 25916
rect 17604 25129 17632 25910
rect 17590 25120 17646 25129
rect 17590 25055 17646 25064
rect 17696 24206 17724 27882
rect 17788 27538 17816 29430
rect 17880 29306 17908 32914
rect 19444 32910 19472 33934
rect 19536 33522 19564 34054
rect 19708 34002 19760 34008
rect 19800 33924 19852 33930
rect 19800 33866 19852 33872
rect 19524 33516 19576 33522
rect 19524 33458 19576 33464
rect 19812 33454 19840 33866
rect 19800 33448 19852 33454
rect 19800 33390 19852 33396
rect 19432 32904 19484 32910
rect 19432 32846 19484 32852
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 19444 32230 19472 32846
rect 18972 32224 19024 32230
rect 18972 32166 19024 32172
rect 19432 32224 19484 32230
rect 19432 32166 19484 32172
rect 18984 32026 19012 32166
rect 18512 32020 18564 32026
rect 18512 31962 18564 31968
rect 18972 32020 19024 32026
rect 18972 31962 19024 31968
rect 18524 31754 18552 31962
rect 19444 31822 19472 32166
rect 19708 31884 19760 31890
rect 19708 31826 19760 31832
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 18524 31726 18736 31754
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 18708 31278 18736 31726
rect 18972 31680 19024 31686
rect 18972 31622 19024 31628
rect 18984 31414 19012 31622
rect 18972 31408 19024 31414
rect 18972 31350 19024 31356
rect 18696 31272 18748 31278
rect 18696 31214 18748 31220
rect 18708 30938 18736 31214
rect 18984 30938 19012 31350
rect 18696 30932 18748 30938
rect 18696 30874 18748 30880
rect 18972 30932 19024 30938
rect 18972 30874 19024 30880
rect 18984 30666 19012 30874
rect 19444 30802 19472 31758
rect 19720 31482 19748 31826
rect 19708 31476 19760 31482
rect 19708 31418 19760 31424
rect 19432 30796 19484 30802
rect 19432 30738 19484 30744
rect 18972 30660 19024 30666
rect 18972 30602 19024 30608
rect 18788 30592 18840 30598
rect 18788 30534 18840 30540
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 18328 30320 18380 30326
rect 18328 30262 18380 30268
rect 18340 29578 18368 30262
rect 18420 29776 18472 29782
rect 18420 29718 18472 29724
rect 18328 29572 18380 29578
rect 18328 29514 18380 29520
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 17868 29300 17920 29306
rect 17868 29242 17920 29248
rect 17868 29164 17920 29170
rect 17868 29106 17920 29112
rect 17776 27532 17828 27538
rect 17776 27474 17828 27480
rect 17776 25764 17828 25770
rect 17776 25706 17828 25712
rect 17788 25294 17816 25706
rect 17776 25288 17828 25294
rect 17776 25230 17828 25236
rect 17880 24732 17908 29106
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 17960 28008 18012 28014
rect 17960 27950 18012 27956
rect 17972 27470 18000 27950
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 18328 26240 18380 26246
rect 18328 26182 18380 26188
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 18340 26042 18368 26182
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 18432 25974 18460 29718
rect 18800 29510 18828 30534
rect 18984 30394 19012 30602
rect 18972 30388 19024 30394
rect 18972 30330 19024 30336
rect 19800 30048 19852 30054
rect 19800 29990 19852 29996
rect 19340 29708 19392 29714
rect 19340 29650 19392 29656
rect 18880 29640 18932 29646
rect 18880 29582 18932 29588
rect 18788 29504 18840 29510
rect 18616 29464 18788 29492
rect 18512 27872 18564 27878
rect 18512 27814 18564 27820
rect 18420 25968 18472 25974
rect 18420 25910 18472 25916
rect 18524 25786 18552 27814
rect 18616 25838 18644 29464
rect 18788 29446 18840 29452
rect 18892 28762 18920 29582
rect 19156 29504 19208 29510
rect 19156 29446 19208 29452
rect 19168 29306 19196 29446
rect 19156 29300 19208 29306
rect 19156 29242 19208 29248
rect 18880 28756 18932 28762
rect 18880 28698 18932 28704
rect 18972 28620 19024 28626
rect 18972 28562 19024 28568
rect 18880 28484 18932 28490
rect 18880 28426 18932 28432
rect 18696 28416 18748 28422
rect 18696 28358 18748 28364
rect 18432 25758 18552 25786
rect 18604 25832 18656 25838
rect 18604 25774 18656 25780
rect 18328 25288 18380 25294
rect 18328 25230 18380 25236
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 18340 24954 18368 25230
rect 18328 24948 18380 24954
rect 18328 24890 18380 24896
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 17788 24704 17908 24732
rect 18144 24744 18196 24750
rect 17684 24200 17736 24206
rect 17684 24142 17736 24148
rect 17592 20800 17644 20806
rect 17592 20742 17644 20748
rect 17604 20534 17632 20742
rect 17592 20528 17644 20534
rect 17592 20470 17644 20476
rect 17512 20318 17632 20346
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17368 18720 17448 18748
rect 17316 18702 17368 18708
rect 17224 17808 17276 17814
rect 17224 17750 17276 17756
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17222 16280 17278 16289
rect 17222 16215 17278 16224
rect 17236 16182 17264 16215
rect 17224 16176 17276 16182
rect 17224 16118 17276 16124
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 17236 15162 17264 16118
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17328 15337 17356 15846
rect 17314 15328 17370 15337
rect 17314 15263 17370 15272
rect 17224 15156 17276 15162
rect 17224 15098 17276 15104
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17144 14006 17172 14418
rect 17132 14000 17184 14006
rect 17132 13942 17184 13948
rect 17132 13456 17184 13462
rect 17132 13398 17184 13404
rect 17144 12714 17172 13398
rect 17420 12986 17448 17478
rect 17512 15366 17540 18770
rect 17604 18630 17632 20318
rect 17592 18624 17644 18630
rect 17592 18566 17644 18572
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17604 17338 17632 17682
rect 17696 17610 17724 24142
rect 17788 23866 17816 24704
rect 18144 24686 18196 24692
rect 18156 24614 18184 24686
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 18144 24608 18196 24614
rect 18144 24550 18196 24556
rect 17776 23860 17828 23866
rect 17776 23802 17828 23808
rect 17788 23526 17816 23802
rect 17776 23520 17828 23526
rect 17776 23462 17828 23468
rect 17788 22982 17816 23462
rect 17776 22976 17828 22982
rect 17776 22918 17828 22924
rect 17880 19922 17908 24550
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 18340 23118 18368 24754
rect 18432 24018 18460 25758
rect 18708 25242 18736 28358
rect 18892 28218 18920 28426
rect 18880 28212 18932 28218
rect 18880 28154 18932 28160
rect 18788 28076 18840 28082
rect 18788 28018 18840 28024
rect 18800 27878 18828 28018
rect 18788 27872 18840 27878
rect 18788 27814 18840 27820
rect 18616 25214 18736 25242
rect 18512 25152 18564 25158
rect 18512 25094 18564 25100
rect 18524 24206 18552 25094
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 18432 23990 18552 24018
rect 18420 23180 18472 23186
rect 18420 23122 18472 23128
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 18340 22778 18368 23054
rect 18328 22772 18380 22778
rect 18328 22714 18380 22720
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18432 20466 18460 23122
rect 18420 20460 18472 20466
rect 18420 20402 18472 20408
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17788 17610 17816 18702
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 18340 17814 18368 18022
rect 17868 17808 17920 17814
rect 17868 17750 17920 17756
rect 18328 17808 18380 17814
rect 18328 17750 18380 17756
rect 17684 17604 17736 17610
rect 17684 17546 17736 17552
rect 17776 17604 17828 17610
rect 17776 17546 17828 17552
rect 17880 17542 17908 17750
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 17604 13870 17632 17274
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17776 16720 17828 16726
rect 17776 16662 17828 16668
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17498 13560 17554 13569
rect 17498 13495 17554 13504
rect 17512 13326 17540 13495
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17132 12708 17184 12714
rect 17132 12650 17184 12656
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 17236 11558 17264 12786
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17328 12238 17356 12378
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16960 10062 16988 11154
rect 17236 10810 17264 11290
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 17052 10169 17080 10610
rect 17038 10160 17094 10169
rect 17038 10095 17094 10104
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16684 6730 16712 7142
rect 16672 6724 16724 6730
rect 16672 6666 16724 6672
rect 16684 5642 16712 6666
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 16684 4486 16712 5578
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 16592 800 16620 3062
rect 16776 2446 16804 9862
rect 16960 9518 16988 9998
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16868 8838 16896 9318
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16868 8566 16896 8774
rect 16856 8560 16908 8566
rect 16856 8502 16908 8508
rect 16960 6798 16988 9454
rect 17132 9376 17184 9382
rect 17132 9318 17184 9324
rect 17144 8974 17172 9318
rect 17420 9178 17448 11018
rect 17512 9654 17540 11086
rect 17696 10810 17724 15846
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17696 10656 17724 10746
rect 17788 10742 17816 16662
rect 17880 16658 17908 17070
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 18248 15450 18276 15642
rect 18340 15570 18368 17750
rect 18328 15564 18380 15570
rect 18328 15506 18380 15512
rect 18248 15422 18368 15450
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17880 11778 17908 13806
rect 18340 13734 18368 15422
rect 18328 13728 18380 13734
rect 18432 13705 18460 19654
rect 18328 13670 18380 13676
rect 18418 13696 18474 13705
rect 18418 13631 18474 13640
rect 18328 13252 18380 13258
rect 18328 13194 18380 13200
rect 18420 13252 18472 13258
rect 18420 13194 18472 13200
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17880 11750 18000 11778
rect 17868 11688 17920 11694
rect 17868 11630 17920 11636
rect 17880 11286 17908 11630
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 17972 11064 18000 11750
rect 17880 11036 18000 11064
rect 17880 10792 17908 11036
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17880 10764 18000 10792
rect 17776 10736 17828 10742
rect 17776 10678 17828 10684
rect 17604 10628 17724 10656
rect 17604 10554 17632 10628
rect 17604 10526 17816 10554
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17592 10192 17644 10198
rect 17592 10134 17644 10140
rect 17604 9926 17632 10134
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17500 9648 17552 9654
rect 17500 9590 17552 9596
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16960 5778 16988 6734
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16868 4758 16896 5510
rect 16856 4752 16908 4758
rect 16856 4694 16908 4700
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16960 800 16988 2790
rect 17052 1970 17080 7142
rect 17144 3466 17172 8910
rect 17512 8906 17540 9114
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17222 8528 17278 8537
rect 17222 8463 17224 8472
rect 17276 8463 17278 8472
rect 17224 8434 17276 8440
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17420 6866 17448 8366
rect 17604 7342 17632 9318
rect 17592 7336 17644 7342
rect 17592 7278 17644 7284
rect 17408 6860 17460 6866
rect 17408 6802 17460 6808
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17236 4282 17264 6258
rect 17316 6248 17368 6254
rect 17316 6190 17368 6196
rect 17328 5370 17356 6190
rect 17420 5914 17448 6802
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 17408 3664 17460 3670
rect 17512 3641 17540 3878
rect 17408 3606 17460 3612
rect 17498 3632 17554 3641
rect 17132 3460 17184 3466
rect 17132 3402 17184 3408
rect 17224 2916 17276 2922
rect 17224 2858 17276 2864
rect 17236 2774 17264 2858
rect 17236 2746 17356 2774
rect 17328 2514 17356 2746
rect 17316 2508 17368 2514
rect 17316 2450 17368 2456
rect 17420 2258 17448 3606
rect 17696 3602 17724 10406
rect 17788 8838 17816 10526
rect 17972 9976 18000 10764
rect 18340 10742 18368 13194
rect 18432 12186 18460 13194
rect 18524 12442 18552 23990
rect 18616 19854 18644 25214
rect 18800 24954 18828 27814
rect 18892 27674 18920 28154
rect 18880 27668 18932 27674
rect 18880 27610 18932 27616
rect 18892 27062 18920 27610
rect 18880 27056 18932 27062
rect 18880 26998 18932 27004
rect 18984 26790 19012 28562
rect 19352 28558 19380 29650
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 19156 27872 19208 27878
rect 19156 27814 19208 27820
rect 18972 26784 19024 26790
rect 18972 26726 19024 26732
rect 18880 26036 18932 26042
rect 18880 25978 18932 25984
rect 18892 25498 18920 25978
rect 18880 25492 18932 25498
rect 18880 25434 18932 25440
rect 18788 24948 18840 24954
rect 18788 24890 18840 24896
rect 18892 24886 18920 25434
rect 18880 24880 18932 24886
rect 18880 24822 18932 24828
rect 18696 24608 18748 24614
rect 18696 24550 18748 24556
rect 18708 22982 18736 24550
rect 18984 24274 19012 26726
rect 19064 25220 19116 25226
rect 19064 25162 19116 25168
rect 18972 24268 19024 24274
rect 18972 24210 19024 24216
rect 18880 24132 18932 24138
rect 18880 24074 18932 24080
rect 18788 24064 18840 24070
rect 18788 24006 18840 24012
rect 18800 23866 18828 24006
rect 18892 23866 18920 24074
rect 19076 23866 19104 25162
rect 19168 24426 19196 27814
rect 19352 27146 19380 28494
rect 19708 28416 19760 28422
rect 19708 28358 19760 28364
rect 19720 28218 19748 28358
rect 19708 28212 19760 28218
rect 19708 28154 19760 28160
rect 19260 27130 19472 27146
rect 19248 27124 19472 27130
rect 19300 27118 19472 27124
rect 19248 27066 19300 27072
rect 19444 26450 19472 27118
rect 19432 26444 19484 26450
rect 19432 26386 19484 26392
rect 19340 25220 19392 25226
rect 19340 25162 19392 25168
rect 19352 24954 19380 25162
rect 19340 24948 19392 24954
rect 19340 24890 19392 24896
rect 19444 24818 19472 26386
rect 19432 24812 19484 24818
rect 19432 24754 19484 24760
rect 19168 24398 19288 24426
rect 19156 24336 19208 24342
rect 19156 24278 19208 24284
rect 18788 23860 18840 23866
rect 18788 23802 18840 23808
rect 18880 23860 18932 23866
rect 18880 23802 18932 23808
rect 19064 23860 19116 23866
rect 19064 23802 19116 23808
rect 18696 22976 18748 22982
rect 18696 22918 18748 22924
rect 18708 22642 18736 22918
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18800 22094 18828 23802
rect 18892 23497 18920 23802
rect 19064 23520 19116 23526
rect 18878 23488 18934 23497
rect 19064 23462 19116 23468
rect 18878 23423 18934 23432
rect 18880 23248 18932 23254
rect 18880 23190 18932 23196
rect 18708 22066 18828 22094
rect 18708 20942 18736 22066
rect 18696 20936 18748 20942
rect 18696 20878 18748 20884
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18788 20460 18840 20466
rect 18788 20402 18840 20408
rect 18708 20262 18736 20402
rect 18696 20256 18748 20262
rect 18696 20198 18748 20204
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18708 18222 18736 20198
rect 18696 18216 18748 18222
rect 18696 18158 18748 18164
rect 18696 17536 18748 17542
rect 18696 17478 18748 17484
rect 18708 16998 18736 17478
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18708 16250 18736 16390
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 18800 16046 18828 20402
rect 18892 17746 18920 23190
rect 18972 22976 19024 22982
rect 18972 22918 19024 22924
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 18984 17270 19012 22918
rect 19076 22778 19104 23462
rect 19064 22772 19116 22778
rect 19064 22714 19116 22720
rect 19062 22672 19118 22681
rect 19062 22607 19118 22616
rect 19076 21486 19104 22607
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 19076 21350 19104 21422
rect 19064 21344 19116 21350
rect 19064 21286 19116 21292
rect 19076 21146 19104 21286
rect 19064 21140 19116 21146
rect 19064 21082 19116 21088
rect 19168 20466 19196 24278
rect 19260 24206 19288 24398
rect 19444 24274 19472 24754
rect 19432 24268 19484 24274
rect 19432 24210 19484 24216
rect 19248 24200 19300 24206
rect 19248 24142 19300 24148
rect 19248 23520 19300 23526
rect 19248 23462 19300 23468
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 19260 23118 19288 23462
rect 19248 23112 19300 23118
rect 19248 23054 19300 23060
rect 19248 22772 19300 22778
rect 19248 22714 19300 22720
rect 19260 20942 19288 22714
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 18972 17264 19024 17270
rect 18972 17206 19024 17212
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18696 15972 18748 15978
rect 18696 15914 18748 15920
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18512 12436 18564 12442
rect 18616 12434 18644 15846
rect 18708 13326 18736 15914
rect 18892 13870 18920 17070
rect 18972 16992 19024 16998
rect 18972 16934 19024 16940
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18616 12406 18736 12434
rect 18512 12378 18564 12384
rect 18604 12368 18656 12374
rect 18604 12310 18656 12316
rect 18432 12158 18552 12186
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18432 11898 18460 12038
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18524 11558 18552 12158
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 18616 11218 18644 12310
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18328 10736 18380 10742
rect 18328 10678 18380 10684
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 18064 10033 18092 10406
rect 18432 10282 18460 10746
rect 18604 10736 18656 10742
rect 18604 10678 18656 10684
rect 18432 10254 18552 10282
rect 18328 10192 18380 10198
rect 18328 10134 18380 10140
rect 17880 9948 18000 9976
rect 18050 10024 18106 10033
rect 18050 9959 18106 9968
rect 17880 9674 17908 9948
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17880 9646 18000 9674
rect 17972 9382 18000 9646
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 18064 9194 18092 9590
rect 17880 9166 18092 9194
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17776 8356 17828 8362
rect 17776 8298 17828 8304
rect 17788 8090 17816 8298
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 17788 4146 17816 7210
rect 17880 6866 17908 9166
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17972 8945 18000 8978
rect 17958 8936 18014 8945
rect 17958 8871 18014 8880
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18248 8362 18276 8434
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 17972 7886 18000 8230
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18340 7546 18368 10134
rect 18524 9926 18552 10254
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18420 8492 18472 8498
rect 18420 8434 18472 8440
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17880 6730 17908 6802
rect 17868 6724 17920 6730
rect 17868 6666 17920 6672
rect 17880 6458 17908 6666
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17868 5296 17920 5302
rect 18340 5273 18368 6394
rect 17868 5238 17920 5244
rect 18326 5264 18382 5273
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17498 3567 17554 3576
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 17684 3460 17736 3466
rect 17684 3402 17736 3408
rect 17328 2230 17448 2258
rect 17040 1964 17092 1970
rect 17040 1906 17092 1912
rect 17328 800 17356 2230
rect 17696 800 17724 3402
rect 17880 3194 17908 5238
rect 18326 5199 18382 5208
rect 18432 5098 18460 8434
rect 18524 8362 18552 9862
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18524 6934 18552 7278
rect 18512 6928 18564 6934
rect 18512 6870 18564 6876
rect 18524 5234 18552 6870
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18420 5092 18472 5098
rect 18420 5034 18472 5040
rect 18524 4690 18552 5170
rect 18512 4684 18564 4690
rect 18512 4626 18564 4632
rect 18328 4548 18380 4554
rect 18328 4490 18380 4496
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18340 3670 18368 4490
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 18328 3664 18380 3670
rect 18328 3606 18380 3612
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18432 1170 18460 4014
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18340 1142 18460 1170
rect 18064 870 18184 898
rect 18064 800 18092 870
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18156 762 18184 870
rect 18340 762 18368 1142
rect 18524 1034 18552 3674
rect 18616 3058 18644 10678
rect 18708 10033 18736 12406
rect 18800 12306 18828 12786
rect 18892 12782 18920 13806
rect 18880 12776 18932 12782
rect 18880 12718 18932 12724
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18788 12300 18840 12306
rect 18788 12242 18840 12248
rect 18892 10810 18920 12378
rect 18984 12374 19012 16934
rect 18972 12368 19024 12374
rect 18972 12310 19024 12316
rect 18972 12096 19024 12102
rect 18972 12038 19024 12044
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18800 10169 18828 10610
rect 18786 10160 18842 10169
rect 18786 10095 18842 10104
rect 18694 10024 18750 10033
rect 18694 9959 18750 9968
rect 18786 9888 18842 9897
rect 18786 9823 18842 9832
rect 18694 9480 18750 9489
rect 18694 9415 18750 9424
rect 18708 8906 18736 9415
rect 18696 8900 18748 8906
rect 18696 8842 18748 8848
rect 18800 8022 18828 9823
rect 18878 9752 18934 9761
rect 18878 9687 18934 9696
rect 18892 9518 18920 9687
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 18892 8430 18920 9318
rect 18880 8424 18932 8430
rect 18880 8366 18932 8372
rect 18788 8016 18840 8022
rect 18788 7958 18840 7964
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18800 5710 18828 7686
rect 18880 7472 18932 7478
rect 18880 7414 18932 7420
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18892 3913 18920 7414
rect 18878 3904 18934 3913
rect 18878 3839 18934 3848
rect 18788 3664 18840 3670
rect 18788 3606 18840 3612
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18708 2650 18736 3538
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 18432 1006 18552 1034
rect 18432 800 18460 1006
rect 18800 800 18828 3606
rect 18984 3058 19012 12038
rect 19076 9994 19104 20198
rect 19168 19378 19196 20266
rect 19352 19394 19380 23462
rect 19444 20602 19472 24210
rect 19616 23724 19668 23730
rect 19616 23666 19668 23672
rect 19524 23656 19576 23662
rect 19524 23598 19576 23604
rect 19536 23322 19564 23598
rect 19524 23316 19576 23322
rect 19524 23258 19576 23264
rect 19536 22681 19564 23258
rect 19628 22778 19656 23666
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19522 22672 19578 22681
rect 19522 22607 19578 22616
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19536 19514 19564 21286
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 19616 20800 19668 20806
rect 19616 20742 19668 20748
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 19248 19372 19300 19378
rect 19352 19366 19472 19394
rect 19248 19314 19300 19320
rect 19156 15972 19208 15978
rect 19156 15914 19208 15920
rect 19168 15706 19196 15914
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 19168 14006 19196 15642
rect 19260 15094 19288 19314
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19352 17678 19380 19246
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19444 17490 19472 19366
rect 19352 17462 19472 17490
rect 19352 16182 19380 17462
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19444 16114 19472 16390
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19156 14000 19208 14006
rect 19156 13942 19208 13948
rect 19352 13138 19380 14214
rect 19444 13326 19472 16050
rect 19536 15366 19564 16390
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19628 15162 19656 20742
rect 19720 15434 19748 20946
rect 19812 20466 19840 29990
rect 19904 26586 19932 34190
rect 20180 34082 20208 53994
rect 22100 53984 22152 53990
rect 22100 53926 22152 53932
rect 21088 43716 21140 43722
rect 21088 43658 21140 43664
rect 20260 41472 20312 41478
rect 20260 41414 20312 41420
rect 20088 34054 20208 34082
rect 20088 30682 20116 34054
rect 20088 30654 20208 30682
rect 20076 30592 20128 30598
rect 20076 30534 20128 30540
rect 20088 30394 20116 30534
rect 20076 30388 20128 30394
rect 20076 30330 20128 30336
rect 19984 30184 20036 30190
rect 19984 30126 20036 30132
rect 19996 29510 20024 30126
rect 19984 29504 20036 29510
rect 19984 29446 20036 29452
rect 19996 29238 20024 29446
rect 19984 29232 20036 29238
rect 19984 29174 20036 29180
rect 19984 27668 20036 27674
rect 19984 27610 20036 27616
rect 19996 27384 20024 27610
rect 20076 27396 20128 27402
rect 19996 27356 20076 27384
rect 19996 27130 20024 27356
rect 20076 27338 20128 27344
rect 19984 27124 20036 27130
rect 19984 27066 20036 27072
rect 19892 26580 19944 26586
rect 19892 26522 19944 26528
rect 19996 26568 20024 27066
rect 20076 26580 20128 26586
rect 19996 26540 20076 26568
rect 19996 26314 20024 26540
rect 20076 26522 20128 26528
rect 19984 26308 20036 26314
rect 19984 26250 20036 26256
rect 20180 26042 20208 30654
rect 20168 26036 20220 26042
rect 20168 25978 20220 25984
rect 20076 25220 20128 25226
rect 20076 25162 20128 25168
rect 19892 25152 19944 25158
rect 19892 25094 19944 25100
rect 19904 24993 19932 25094
rect 19890 24984 19946 24993
rect 19890 24919 19946 24928
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19904 23662 19932 24006
rect 19892 23656 19944 23662
rect 19892 23598 19944 23604
rect 20088 21894 20116 25162
rect 20180 25106 20208 25978
rect 20272 25498 20300 41414
rect 20628 35488 20680 35494
rect 20628 35430 20680 35436
rect 20444 35012 20496 35018
rect 20444 34954 20496 34960
rect 20456 31346 20484 34954
rect 20536 33448 20588 33454
rect 20536 33390 20588 33396
rect 20444 31340 20496 31346
rect 20444 31282 20496 31288
rect 20456 31142 20484 31282
rect 20444 31136 20496 31142
rect 20444 31078 20496 31084
rect 20548 30190 20576 33390
rect 20536 30184 20588 30190
rect 20536 30126 20588 30132
rect 20640 29306 20668 35430
rect 20812 34740 20864 34746
rect 20812 34682 20864 34688
rect 20824 29646 20852 34682
rect 21100 34406 21128 43658
rect 21364 41540 21416 41546
rect 21364 41482 21416 41488
rect 21376 35894 21404 41482
rect 21916 39296 21968 39302
rect 21916 39238 21968 39244
rect 21284 35866 21404 35894
rect 21180 35488 21232 35494
rect 21180 35430 21232 35436
rect 21088 34400 21140 34406
rect 21088 34342 21140 34348
rect 21192 33862 21220 35430
rect 21180 33856 21232 33862
rect 21180 33798 21232 33804
rect 21192 32366 21220 33798
rect 21180 32360 21232 32366
rect 21180 32302 21232 32308
rect 20904 32224 20956 32230
rect 20904 32166 20956 32172
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20628 29300 20680 29306
rect 20628 29242 20680 29248
rect 20352 29232 20404 29238
rect 20352 29174 20404 29180
rect 20260 25492 20312 25498
rect 20260 25434 20312 25440
rect 20272 25294 20300 25434
rect 20260 25288 20312 25294
rect 20260 25230 20312 25236
rect 20180 25078 20300 25106
rect 20168 22568 20220 22574
rect 20168 22510 20220 22516
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 20088 21622 20116 21830
rect 20076 21616 20128 21622
rect 20076 21558 20128 21564
rect 20180 21486 20208 22510
rect 20272 21894 20300 25078
rect 20364 23730 20392 29174
rect 20916 29102 20944 32166
rect 20996 31680 21048 31686
rect 20996 31622 21048 31628
rect 21008 30666 21036 31622
rect 21180 31136 21232 31142
rect 21180 31078 21232 31084
rect 20996 30660 21048 30666
rect 20996 30602 21048 30608
rect 20904 29096 20956 29102
rect 20904 29038 20956 29044
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20640 28150 20668 28494
rect 20916 28490 20944 29038
rect 21008 28626 21036 30602
rect 20996 28620 21048 28626
rect 20996 28562 21048 28568
rect 20904 28484 20956 28490
rect 20904 28426 20956 28432
rect 20628 28144 20680 28150
rect 20628 28086 20680 28092
rect 21088 26512 21140 26518
rect 21088 26454 21140 26460
rect 20996 26444 21048 26450
rect 20996 26386 21048 26392
rect 20444 24744 20496 24750
rect 20444 24686 20496 24692
rect 20456 24410 20484 24686
rect 20444 24404 20496 24410
rect 20444 24346 20496 24352
rect 20352 23724 20404 23730
rect 20352 23666 20404 23672
rect 20456 23186 20484 24346
rect 20812 23724 20864 23730
rect 20812 23666 20864 23672
rect 20824 23186 20852 23666
rect 21008 23662 21036 26386
rect 21100 24818 21128 26454
rect 21192 25702 21220 31078
rect 21180 25696 21232 25702
rect 21180 25638 21232 25644
rect 21088 24812 21140 24818
rect 21088 24754 21140 24760
rect 21100 24342 21128 24754
rect 21088 24336 21140 24342
rect 21088 24278 21140 24284
rect 20996 23656 21048 23662
rect 20996 23598 21048 23604
rect 20444 23180 20496 23186
rect 20444 23122 20496 23128
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20812 22704 20864 22710
rect 20812 22646 20864 22652
rect 20720 22432 20772 22438
rect 20720 22374 20772 22380
rect 20352 22092 20404 22098
rect 20352 22034 20404 22040
rect 20260 21888 20312 21894
rect 20260 21830 20312 21836
rect 20272 21690 20300 21830
rect 20260 21684 20312 21690
rect 20260 21626 20312 21632
rect 20168 21480 20220 21486
rect 20168 21422 20220 21428
rect 19800 20460 19852 20466
rect 19800 20402 19852 20408
rect 19800 20256 19852 20262
rect 19800 20198 19852 20204
rect 19812 16726 19840 20198
rect 20180 19786 20208 21422
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 19892 17536 19944 17542
rect 19892 17478 19944 17484
rect 19800 16720 19852 16726
rect 19800 16662 19852 16668
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 19708 15428 19760 15434
rect 19708 15370 19760 15376
rect 19616 15156 19668 15162
rect 19616 15098 19668 15104
rect 19524 14544 19576 14550
rect 19524 14486 19576 14492
rect 19536 14006 19564 14486
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19628 14006 19656 14350
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 19616 14000 19668 14006
rect 19616 13942 19668 13948
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19352 13110 19564 13138
rect 19430 13016 19486 13025
rect 19430 12951 19432 12960
rect 19484 12951 19486 12960
rect 19432 12922 19484 12928
rect 19248 12776 19300 12782
rect 19248 12718 19300 12724
rect 19260 12238 19288 12718
rect 19432 12640 19484 12646
rect 19432 12582 19484 12588
rect 19444 12434 19472 12582
rect 19352 12406 19472 12434
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19064 9988 19116 9994
rect 19064 9930 19116 9936
rect 19064 9648 19116 9654
rect 19064 9590 19116 9596
rect 19076 8401 19104 9590
rect 19062 8392 19118 8401
rect 19062 8327 19118 8336
rect 19064 8084 19116 8090
rect 19064 8026 19116 8032
rect 19076 7546 19104 8026
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 19168 4026 19196 11494
rect 19352 11014 19380 12406
rect 19536 11898 19564 13110
rect 19720 12170 19748 15370
rect 19812 13025 19840 16050
rect 19904 14958 19932 17478
rect 20180 17338 20208 19722
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20272 16658 20300 19858
rect 20364 16998 20392 22034
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20548 18714 20576 20198
rect 20732 19514 20760 22374
rect 20824 20602 20852 22646
rect 20904 22636 20956 22642
rect 20904 22578 20956 22584
rect 21088 22636 21140 22642
rect 21192 22624 21220 25638
rect 21140 22596 21220 22624
rect 21088 22578 21140 22584
rect 20916 21146 20944 22578
rect 21100 22506 21128 22578
rect 21088 22500 21140 22506
rect 21088 22442 21140 22448
rect 21180 21956 21232 21962
rect 21180 21898 21232 21904
rect 20904 21140 20956 21146
rect 20904 21082 20956 21088
rect 20916 20602 20944 21082
rect 20996 20936 21048 20942
rect 20996 20878 21048 20884
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 21008 20398 21036 20878
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20548 18686 20668 18714
rect 20536 18624 20588 18630
rect 20536 18566 20588 18572
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20260 16652 20312 16658
rect 20260 16594 20312 16600
rect 20272 16182 20300 16594
rect 20444 16516 20496 16522
rect 20444 16458 20496 16464
rect 20260 16176 20312 16182
rect 20260 16118 20312 16124
rect 20272 15570 20300 16118
rect 20456 15706 20484 16458
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20260 15564 20312 15570
rect 20260 15506 20312 15512
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19892 14272 19944 14278
rect 19892 14214 19944 14220
rect 19798 13016 19854 13025
rect 19798 12951 19854 12960
rect 19708 12164 19760 12170
rect 19708 12106 19760 12112
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19536 11762 19564 11834
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 19720 11694 19748 12106
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19340 10260 19392 10266
rect 19340 10202 19392 10208
rect 19352 10130 19380 10202
rect 19248 10124 19300 10130
rect 19248 10066 19300 10072
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19260 7342 19288 10066
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 19260 5409 19288 7278
rect 19246 5400 19302 5409
rect 19246 5335 19302 5344
rect 19076 4010 19196 4026
rect 19064 4004 19196 4010
rect 19116 3998 19196 4004
rect 19064 3946 19116 3952
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 19168 800 19196 3878
rect 19352 3534 19380 8842
rect 19340 3528 19392 3534
rect 19340 3470 19392 3476
rect 19444 2446 19472 11494
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19536 10266 19564 10406
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19812 10010 19840 10950
rect 19628 9982 19840 10010
rect 19628 9110 19656 9982
rect 19812 9926 19840 9982
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19800 9920 19852 9926
rect 19800 9862 19852 9868
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 19628 8022 19656 8910
rect 19616 8016 19668 8022
rect 19616 7958 19668 7964
rect 19522 7032 19578 7041
rect 19522 6967 19578 6976
rect 19536 6798 19564 6967
rect 19628 6934 19656 7958
rect 19616 6928 19668 6934
rect 19720 6905 19748 9862
rect 19904 9674 19932 14214
rect 19996 11830 20024 14962
rect 20168 14612 20220 14618
rect 20168 14554 20220 14560
rect 20076 13388 20128 13394
rect 20076 13330 20128 13336
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 20088 11762 20116 13330
rect 20180 12238 20208 14554
rect 20364 12434 20392 15302
rect 20456 14958 20484 15642
rect 20444 14952 20496 14958
rect 20444 14894 20496 14900
rect 20444 13388 20496 13394
rect 20444 13330 20496 13336
rect 20272 12406 20392 12434
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20180 11898 20208 12174
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 20076 11756 20128 11762
rect 20076 11698 20128 11704
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19996 11150 20024 11630
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 20168 11008 20220 11014
rect 20088 10968 20168 10996
rect 19982 10704 20038 10713
rect 19982 10639 19984 10648
rect 20036 10639 20038 10648
rect 19984 10610 20036 10616
rect 20088 10606 20116 10968
rect 20168 10950 20220 10956
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20076 10600 20128 10606
rect 20076 10542 20128 10548
rect 20180 9926 20208 10746
rect 20272 10130 20300 12406
rect 20456 12306 20484 13330
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20352 10192 20404 10198
rect 20352 10134 20404 10140
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 20180 9722 20208 9862
rect 20272 9722 20300 10066
rect 20168 9716 20220 9722
rect 19904 9646 20116 9674
rect 20168 9658 20220 9664
rect 20260 9716 20312 9722
rect 20260 9658 20312 9664
rect 19800 9376 19852 9382
rect 19800 9318 19852 9324
rect 19812 9058 19840 9318
rect 20088 9178 20116 9646
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20076 9172 20128 9178
rect 20076 9114 20128 9120
rect 19812 9030 19932 9058
rect 19800 8900 19852 8906
rect 19800 8842 19852 8848
rect 19812 7342 19840 8842
rect 19904 7750 19932 9030
rect 19892 7744 19944 7750
rect 19892 7686 19944 7692
rect 19904 7410 19932 7686
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19812 6934 19840 7278
rect 19904 7002 19932 7346
rect 19892 6996 19944 7002
rect 19892 6938 19944 6944
rect 19800 6928 19852 6934
rect 19616 6870 19668 6876
rect 19706 6896 19762 6905
rect 19800 6870 19852 6876
rect 19706 6831 19762 6840
rect 19892 6860 19944 6866
rect 19944 6820 20024 6848
rect 19892 6802 19944 6808
rect 19524 6792 19576 6798
rect 19524 6734 19576 6740
rect 19524 6656 19576 6662
rect 19800 6656 19852 6662
rect 19576 6633 19748 6644
rect 19576 6624 19762 6633
rect 19576 6616 19706 6624
rect 19524 6598 19576 6604
rect 19800 6598 19852 6604
rect 19706 6559 19762 6568
rect 19524 6452 19576 6458
rect 19524 6394 19576 6400
rect 19536 3602 19564 6394
rect 19812 6202 19840 6598
rect 19628 6174 19840 6202
rect 19628 6118 19656 6174
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19800 6112 19852 6118
rect 19800 6054 19852 6060
rect 19706 4584 19762 4593
rect 19812 4554 19840 6054
rect 19996 5914 20024 6820
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 19996 5817 20024 5850
rect 19982 5808 20038 5817
rect 19892 5772 19944 5778
rect 19982 5743 20038 5752
rect 19892 5714 19944 5720
rect 19706 4519 19708 4528
rect 19760 4519 19762 4528
rect 19800 4548 19852 4554
rect 19708 4490 19760 4496
rect 19800 4490 19852 4496
rect 19904 3942 19932 5714
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19524 2916 19576 2922
rect 19524 2858 19576 2864
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19536 800 19564 2858
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 19904 2514 19932 2790
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 19996 2258 20024 4422
rect 20088 3602 20116 9114
rect 20168 6996 20220 7002
rect 20168 6938 20220 6944
rect 20180 5234 20208 6938
rect 20272 6882 20300 9522
rect 20364 7478 20392 10134
rect 20444 9988 20496 9994
rect 20548 9976 20576 18566
rect 20640 14482 20668 18686
rect 20812 18148 20864 18154
rect 20812 18090 20864 18096
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20628 13728 20680 13734
rect 20628 13670 20680 13676
rect 20640 12918 20668 13670
rect 20732 13258 20760 17818
rect 20824 17270 20852 18090
rect 21088 18080 21140 18086
rect 21086 18048 21088 18057
rect 21140 18048 21142 18057
rect 21086 17983 21142 17992
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 20812 17264 20864 17270
rect 20812 17206 20864 17212
rect 20824 15978 20852 17206
rect 20904 17060 20956 17066
rect 20904 17002 20956 17008
rect 20812 15972 20864 15978
rect 20812 15914 20864 15920
rect 20824 15502 20852 15914
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20916 13818 20944 17002
rect 21100 15502 21128 17478
rect 21192 16046 21220 21898
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 21100 13938 21128 15098
rect 21284 14346 21312 35866
rect 21824 35692 21876 35698
rect 21824 35634 21876 35640
rect 21836 34950 21864 35634
rect 21824 34944 21876 34950
rect 21744 34904 21824 34932
rect 21364 34400 21416 34406
rect 21364 34342 21416 34348
rect 21376 33930 21404 34342
rect 21364 33924 21416 33930
rect 21364 33866 21416 33872
rect 21376 33590 21404 33866
rect 21364 33584 21416 33590
rect 21364 33526 21416 33532
rect 21376 33318 21404 33526
rect 21364 33312 21416 33318
rect 21364 33254 21416 33260
rect 21376 32230 21404 33254
rect 21456 32292 21508 32298
rect 21456 32234 21508 32240
rect 21364 32224 21416 32230
rect 21364 32166 21416 32172
rect 21376 31754 21404 32166
rect 21468 32026 21496 32234
rect 21456 32020 21508 32026
rect 21456 31962 21508 31968
rect 21364 31748 21416 31754
rect 21364 31690 21416 31696
rect 21376 31482 21404 31690
rect 21640 31680 21692 31686
rect 21640 31622 21692 31628
rect 21364 31476 21416 31482
rect 21364 31418 21416 31424
rect 21376 30802 21404 31418
rect 21364 30796 21416 30802
rect 21364 30738 21416 30744
rect 21364 28620 21416 28626
rect 21364 28562 21416 28568
rect 21376 23730 21404 28562
rect 21652 28422 21680 31622
rect 21744 31482 21772 34904
rect 21824 34886 21876 34892
rect 21824 32768 21876 32774
rect 21824 32710 21876 32716
rect 21836 32434 21864 32710
rect 21824 32428 21876 32434
rect 21824 32370 21876 32376
rect 21836 32230 21864 32370
rect 21824 32224 21876 32230
rect 21824 32166 21876 32172
rect 21732 31476 21784 31482
rect 21732 31418 21784 31424
rect 21836 29034 21864 32166
rect 21928 31890 21956 39238
rect 22008 35488 22060 35494
rect 22008 35430 22060 35436
rect 21916 31884 21968 31890
rect 21916 31826 21968 31832
rect 22020 31754 22048 35430
rect 21928 31726 22048 31754
rect 21928 30326 21956 31726
rect 22008 31680 22060 31686
rect 22008 31622 22060 31628
rect 22020 31482 22048 31622
rect 22008 31476 22060 31482
rect 22008 31418 22060 31424
rect 21916 30320 21968 30326
rect 21916 30262 21968 30268
rect 22112 30122 22140 53926
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 23400 53582 23428 56063
rect 24504 55214 24532 56200
rect 24766 55448 24822 55457
rect 24766 55383 24822 55392
rect 24412 55186 24532 55214
rect 23388 53576 23440 53582
rect 23388 53518 23440 53524
rect 22836 53440 22888 53446
rect 22836 53382 22888 53388
rect 23940 53440 23992 53446
rect 23940 53382 23992 53388
rect 22848 44198 22876 53382
rect 23756 52896 23808 52902
rect 23756 52838 23808 52844
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 23388 51808 23440 51814
rect 23388 51750 23440 51756
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 23400 48142 23428 51750
rect 23388 48136 23440 48142
rect 23388 48078 23440 48084
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 22836 44192 22888 44198
rect 22836 44134 22888 44140
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 23296 40180 23348 40186
rect 23296 40122 23348 40128
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 22192 35624 22244 35630
rect 22192 35566 22244 35572
rect 22560 35624 22612 35630
rect 22560 35566 22612 35572
rect 22204 32026 22232 35566
rect 22468 34944 22520 34950
rect 22468 34886 22520 34892
rect 22284 34060 22336 34066
rect 22284 34002 22336 34008
rect 22296 33590 22324 34002
rect 22284 33584 22336 33590
rect 22284 33526 22336 33532
rect 22296 32978 22324 33526
rect 22376 33448 22428 33454
rect 22376 33390 22428 33396
rect 22388 33114 22416 33390
rect 22376 33108 22428 33114
rect 22376 33050 22428 33056
rect 22284 32972 22336 32978
rect 22284 32914 22336 32920
rect 22296 32502 22324 32914
rect 22284 32496 22336 32502
rect 22284 32438 22336 32444
rect 22192 32020 22244 32026
rect 22192 31962 22244 31968
rect 22100 30116 22152 30122
rect 22100 30058 22152 30064
rect 21916 30048 21968 30054
rect 21916 29990 21968 29996
rect 21824 29028 21876 29034
rect 21824 28970 21876 28976
rect 21640 28416 21692 28422
rect 21640 28358 21692 28364
rect 21732 28416 21784 28422
rect 21732 28358 21784 28364
rect 21640 27328 21692 27334
rect 21640 27270 21692 27276
rect 21652 26450 21680 27270
rect 21744 26772 21772 28358
rect 21836 28082 21864 28970
rect 21824 28076 21876 28082
rect 21824 28018 21876 28024
rect 21824 26784 21876 26790
rect 21744 26744 21824 26772
rect 21824 26726 21876 26732
rect 21836 26518 21864 26726
rect 21824 26512 21876 26518
rect 21824 26454 21876 26460
rect 21640 26444 21692 26450
rect 21640 26386 21692 26392
rect 21640 25696 21692 25702
rect 21640 25638 21692 25644
rect 21456 24336 21508 24342
rect 21456 24278 21508 24284
rect 21468 23730 21496 24278
rect 21364 23724 21416 23730
rect 21364 23666 21416 23672
rect 21456 23724 21508 23730
rect 21456 23666 21508 23672
rect 21468 21690 21496 23666
rect 21652 23118 21680 25638
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21928 22094 21956 29990
rect 22204 28626 22232 31962
rect 22296 31346 22324 32438
rect 22284 31340 22336 31346
rect 22284 31282 22336 31288
rect 22480 30326 22508 34886
rect 22572 33658 22600 35566
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 22744 35148 22796 35154
rect 22744 35090 22796 35096
rect 22560 33652 22612 33658
rect 22560 33594 22612 33600
rect 22756 33114 22784 35090
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 22928 33856 22980 33862
rect 22928 33798 22980 33804
rect 23204 33856 23256 33862
rect 23204 33798 23256 33804
rect 22940 33454 22968 33798
rect 23216 33658 23244 33798
rect 23204 33652 23256 33658
rect 23204 33594 23256 33600
rect 22928 33448 22980 33454
rect 22848 33396 22928 33402
rect 22848 33390 22980 33396
rect 22848 33374 22968 33390
rect 22744 33108 22796 33114
rect 22744 33050 22796 33056
rect 22744 31952 22796 31958
rect 22744 31894 22796 31900
rect 22560 31748 22612 31754
rect 22560 31690 22612 31696
rect 22468 30320 22520 30326
rect 22468 30262 22520 30268
rect 22468 29504 22520 29510
rect 22468 29446 22520 29452
rect 22192 28620 22244 28626
rect 22192 28562 22244 28568
rect 22204 28218 22232 28562
rect 22284 28552 22336 28558
rect 22284 28494 22336 28500
rect 22192 28212 22244 28218
rect 22192 28154 22244 28160
rect 22100 27940 22152 27946
rect 22100 27882 22152 27888
rect 22112 26926 22140 27882
rect 22100 26920 22152 26926
rect 22100 26862 22152 26868
rect 22112 26586 22140 26862
rect 22296 26586 22324 28494
rect 22376 27872 22428 27878
rect 22376 27814 22428 27820
rect 22388 27402 22416 27814
rect 22376 27396 22428 27402
rect 22376 27338 22428 27344
rect 22376 26784 22428 26790
rect 22376 26726 22428 26732
rect 22100 26580 22152 26586
rect 22100 26522 22152 26528
rect 22284 26580 22336 26586
rect 22284 26522 22336 26528
rect 22284 26444 22336 26450
rect 22284 26386 22336 26392
rect 22296 24750 22324 26386
rect 22388 25770 22416 26726
rect 22480 26042 22508 29446
rect 22572 28558 22600 31690
rect 22652 31408 22704 31414
rect 22652 31350 22704 31356
rect 22664 30938 22692 31350
rect 22652 30932 22704 30938
rect 22652 30874 22704 30880
rect 22652 30660 22704 30666
rect 22652 30602 22704 30608
rect 22560 28552 22612 28558
rect 22560 28494 22612 28500
rect 22560 27872 22612 27878
rect 22560 27814 22612 27820
rect 22572 26874 22600 27814
rect 22664 26994 22692 30602
rect 22756 27130 22784 31894
rect 22848 30326 22876 33374
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 23308 31890 23336 40122
rect 23664 33856 23716 33862
rect 23664 33798 23716 33804
rect 23676 33590 23704 33798
rect 23664 33584 23716 33590
rect 23664 33526 23716 33532
rect 23676 33318 23704 33526
rect 23664 33312 23716 33318
rect 23664 33254 23716 33260
rect 23676 32910 23704 33254
rect 23664 32904 23716 32910
rect 23664 32846 23716 32852
rect 23768 32858 23796 52838
rect 23296 31884 23348 31890
rect 23296 31826 23348 31832
rect 23020 31816 23072 31822
rect 23020 31758 23072 31764
rect 23032 31414 23060 31758
rect 23572 31476 23624 31482
rect 23572 31418 23624 31424
rect 23020 31408 23072 31414
rect 23020 31350 23072 31356
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 22836 30320 22888 30326
rect 22836 30262 22888 30268
rect 23584 30190 23612 31418
rect 23676 31362 23704 32846
rect 23768 32830 23888 32858
rect 23860 32774 23888 32830
rect 23848 32768 23900 32774
rect 23848 32710 23900 32716
rect 23952 32570 23980 53382
rect 24412 53038 24440 55186
rect 24490 54632 24546 54641
rect 24490 54567 24546 54576
rect 24504 53786 24532 54567
rect 24780 53786 24808 55383
rect 25884 54194 25912 56200
rect 25872 54188 25924 54194
rect 25872 54130 25924 54136
rect 25044 53984 25096 53990
rect 25044 53926 25096 53932
rect 25320 53984 25372 53990
rect 25320 53926 25372 53932
rect 25056 53825 25084 53926
rect 25042 53816 25098 53825
rect 24492 53780 24544 53786
rect 24492 53722 24544 53728
rect 24768 53780 24820 53786
rect 25042 53751 25098 53760
rect 24768 53722 24820 53728
rect 24504 53582 24532 53722
rect 24492 53576 24544 53582
rect 24492 53518 24544 53524
rect 24780 53106 24808 53722
rect 25056 53582 25084 53751
rect 25044 53576 25096 53582
rect 25044 53518 25096 53524
rect 24768 53100 24820 53106
rect 24768 53042 24820 53048
rect 25044 53100 25096 53106
rect 25044 53042 25096 53048
rect 24400 53032 24452 53038
rect 25056 53009 25084 53042
rect 24400 52974 24452 52980
rect 25042 53000 25098 53009
rect 24412 52698 24440 52974
rect 25042 52935 25098 52944
rect 24492 52896 24544 52902
rect 24492 52838 24544 52844
rect 24400 52692 24452 52698
rect 24400 52634 24452 52640
rect 24032 48000 24084 48006
rect 24032 47942 24084 47948
rect 24044 43858 24072 47942
rect 24032 43852 24084 43858
rect 24032 43794 24084 43800
rect 24216 43104 24268 43110
rect 24216 43046 24268 43052
rect 23940 32564 23992 32570
rect 23940 32506 23992 32512
rect 23676 31346 23888 31362
rect 23676 31340 23900 31346
rect 23676 31334 23848 31340
rect 23848 31282 23900 31288
rect 23860 31142 23888 31282
rect 23848 31136 23900 31142
rect 23848 31078 23900 31084
rect 23860 30938 23888 31078
rect 23848 30932 23900 30938
rect 23848 30874 23900 30880
rect 22836 30184 22888 30190
rect 22836 30126 22888 30132
rect 23572 30184 23624 30190
rect 23572 30126 23624 30132
rect 22848 29102 22876 30126
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 23388 29776 23440 29782
rect 23388 29718 23440 29724
rect 22836 29096 22888 29102
rect 22836 29038 22888 29044
rect 22848 28014 22876 29038
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 22836 28008 22888 28014
rect 22836 27950 22888 27956
rect 22848 27538 22876 27950
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 22836 27532 22888 27538
rect 22888 27492 22968 27520
rect 22836 27474 22888 27480
rect 22744 27124 22796 27130
rect 22744 27066 22796 27072
rect 22940 27062 22968 27492
rect 22928 27056 22980 27062
rect 22928 26998 22980 27004
rect 22652 26988 22704 26994
rect 22652 26930 22704 26936
rect 23296 26988 23348 26994
rect 23296 26930 23348 26936
rect 22572 26846 22692 26874
rect 22560 26512 22612 26518
rect 22560 26454 22612 26460
rect 22468 26036 22520 26042
rect 22468 25978 22520 25984
rect 22376 25764 22428 25770
rect 22376 25706 22428 25712
rect 22468 25696 22520 25702
rect 22468 25638 22520 25644
rect 22376 25356 22428 25362
rect 22376 25298 22428 25304
rect 22284 24744 22336 24750
rect 22284 24686 22336 24692
rect 22100 24608 22152 24614
rect 22100 24550 22152 24556
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 22020 22234 22048 23666
rect 22112 23594 22140 24550
rect 22192 24268 22244 24274
rect 22192 24210 22244 24216
rect 22100 23588 22152 23594
rect 22100 23530 22152 23536
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22112 22642 22140 22918
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 22008 22228 22060 22234
rect 22008 22170 22060 22176
rect 22204 22098 22232 24210
rect 22296 24138 22324 24686
rect 22284 24132 22336 24138
rect 22284 24074 22336 24080
rect 22284 23588 22336 23594
rect 22284 23530 22336 23536
rect 22296 22114 22324 23530
rect 22388 22778 22416 25298
rect 22376 22772 22428 22778
rect 22376 22714 22428 22720
rect 21836 22066 21956 22094
rect 22192 22092 22244 22098
rect 21456 21684 21508 21690
rect 21456 21626 21508 21632
rect 21468 19854 21496 21626
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 21456 19848 21508 19854
rect 21508 19796 21588 19802
rect 21456 19790 21588 19796
rect 21468 19774 21588 19790
rect 21456 19712 21508 19718
rect 21456 19654 21508 19660
rect 21468 17678 21496 19654
rect 21560 19242 21588 19774
rect 21640 19712 21692 19718
rect 21640 19654 21692 19660
rect 21652 19310 21680 19654
rect 21640 19304 21692 19310
rect 21640 19246 21692 19252
rect 21548 19236 21600 19242
rect 21548 19178 21600 19184
rect 21744 17898 21772 21286
rect 21836 20466 21864 22066
rect 22296 22086 22416 22114
rect 22192 22034 22244 22040
rect 22100 21956 22152 21962
rect 22100 21898 22152 21904
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 22020 21010 22048 21490
rect 22112 21146 22140 21898
rect 22204 21622 22232 22034
rect 22284 21956 22336 21962
rect 22284 21898 22336 21904
rect 22296 21690 22324 21898
rect 22284 21684 22336 21690
rect 22284 21626 22336 21632
rect 22192 21616 22244 21622
rect 22192 21558 22244 21564
rect 22100 21140 22152 21146
rect 22100 21082 22152 21088
rect 22008 21004 22060 21010
rect 22008 20946 22060 20952
rect 21824 20460 21876 20466
rect 21824 20402 21876 20408
rect 22112 19310 22140 21082
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22204 20058 22232 20402
rect 22284 20392 22336 20398
rect 22284 20334 22336 20340
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 21824 19236 21876 19242
rect 21824 19178 21876 19184
rect 21916 19236 21968 19242
rect 21916 19178 21968 19184
rect 21652 17870 21772 17898
rect 21548 17808 21600 17814
rect 21548 17750 21600 17756
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21364 16040 21416 16046
rect 21364 15982 21416 15988
rect 21376 15638 21404 15982
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21364 15632 21416 15638
rect 21364 15574 21416 15580
rect 21364 15428 21416 15434
rect 21364 15370 21416 15376
rect 21376 15026 21404 15370
rect 21364 15020 21416 15026
rect 21364 14962 21416 14968
rect 21272 14340 21324 14346
rect 21272 14282 21324 14288
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 20824 13790 20944 13818
rect 20720 13252 20772 13258
rect 20720 13194 20772 13200
rect 20628 12912 20680 12918
rect 20628 12854 20680 12860
rect 20824 12850 20852 13790
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20996 13728 21048 13734
rect 20996 13670 21048 13676
rect 20812 12844 20864 12850
rect 20812 12786 20864 12792
rect 20810 11792 20866 11801
rect 20810 11727 20866 11736
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20640 10606 20668 11222
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20732 9994 20760 11086
rect 20824 11082 20852 11727
rect 20812 11076 20864 11082
rect 20812 11018 20864 11024
rect 20916 10588 20944 13670
rect 21008 11218 21036 13670
rect 21088 13524 21140 13530
rect 21088 13466 21140 13472
rect 21100 12850 21128 13466
rect 21284 12986 21312 13874
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 21180 12708 21232 12714
rect 21180 12650 21232 12656
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 21192 11150 21220 12650
rect 21272 12300 21324 12306
rect 21272 12242 21324 12248
rect 21180 11144 21232 11150
rect 21180 11086 21232 11092
rect 20996 11076 21048 11082
rect 20996 11018 21048 11024
rect 20824 10560 20944 10588
rect 20496 9948 20576 9976
rect 20720 9988 20772 9994
rect 20444 9930 20496 9936
rect 20720 9930 20772 9936
rect 20628 9920 20680 9926
rect 20628 9862 20680 9868
rect 20640 9654 20668 9862
rect 20628 9648 20680 9654
rect 20628 9590 20680 9596
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 20272 6854 20392 6882
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20272 6118 20300 6734
rect 20364 6458 20392 6854
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20456 6390 20484 6802
rect 20444 6384 20496 6390
rect 20350 6352 20406 6361
rect 20444 6326 20496 6332
rect 20350 6287 20406 6296
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 20168 5228 20220 5234
rect 20220 5188 20300 5216
rect 20168 5170 20220 5176
rect 20168 5092 20220 5098
rect 20168 5034 20220 5040
rect 20180 4826 20208 5034
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20272 4554 20300 5188
rect 20260 4548 20312 4554
rect 20260 4490 20312 4496
rect 20272 4282 20300 4490
rect 20260 4276 20312 4282
rect 20260 4218 20312 4224
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 19904 2230 20024 2258
rect 19904 800 19932 2230
rect 20272 800 20300 3674
rect 20364 3233 20392 6287
rect 20442 5400 20498 5409
rect 20442 5335 20444 5344
rect 20496 5335 20498 5344
rect 20444 5306 20496 5312
rect 20548 3398 20576 8366
rect 20824 8362 20852 10560
rect 20904 9988 20956 9994
rect 20904 9930 20956 9936
rect 20916 9178 20944 9930
rect 20904 9172 20956 9178
rect 20904 9114 20956 9120
rect 20812 8356 20864 8362
rect 20812 8298 20864 8304
rect 20720 7812 20772 7818
rect 20720 7754 20772 7760
rect 20732 7410 20760 7754
rect 20720 7404 20772 7410
rect 20720 7346 20772 7352
rect 20718 7032 20774 7041
rect 20718 6967 20774 6976
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20444 3392 20496 3398
rect 20444 3334 20496 3340
rect 20536 3392 20588 3398
rect 20536 3334 20588 3340
rect 20350 3224 20406 3233
rect 20456 3210 20484 3334
rect 20456 3182 20576 3210
rect 20350 3159 20406 3168
rect 20548 3126 20576 3182
rect 20536 3120 20588 3126
rect 20534 3088 20536 3097
rect 20588 3088 20590 3097
rect 20534 3023 20590 3032
rect 20640 800 20668 5646
rect 18156 734 18368 762
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20732 762 20760 6967
rect 20824 5302 20852 8298
rect 21008 6882 21036 11018
rect 21284 10810 21312 12242
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 21100 9722 21128 10610
rect 21284 10606 21312 10746
rect 21272 10600 21324 10606
rect 21272 10542 21324 10548
rect 21088 9716 21140 9722
rect 21088 9658 21140 9664
rect 21088 9512 21140 9518
rect 21088 9454 21140 9460
rect 21180 9512 21232 9518
rect 21180 9454 21232 9460
rect 20916 6854 21036 6882
rect 20916 5574 20944 6854
rect 20994 6624 21050 6633
rect 20994 6559 21050 6568
rect 20904 5568 20956 5574
rect 20904 5510 20956 5516
rect 20812 5296 20864 5302
rect 20812 5238 20864 5244
rect 21008 4146 21036 6559
rect 21100 5234 21128 9454
rect 21088 5228 21140 5234
rect 21088 5170 21140 5176
rect 21100 4321 21128 5170
rect 21086 4312 21142 4321
rect 21086 4247 21142 4256
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 20916 3194 20944 4082
rect 21192 4049 21220 9454
rect 21272 5160 21324 5166
rect 21272 5102 21324 5108
rect 21284 4826 21312 5102
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 21284 4078 21312 4762
rect 21272 4072 21324 4078
rect 21178 4040 21234 4049
rect 21272 4014 21324 4020
rect 21178 3975 21234 3984
rect 21376 3534 21404 11494
rect 21468 9654 21496 15846
rect 21560 14006 21588 17750
rect 21652 14414 21680 17870
rect 21836 17270 21864 19178
rect 21824 17264 21876 17270
rect 21824 17206 21876 17212
rect 21836 16794 21864 17206
rect 21824 16788 21876 16794
rect 21824 16730 21876 16736
rect 21836 16522 21864 16730
rect 21824 16516 21876 16522
rect 21824 16458 21876 16464
rect 21836 16182 21864 16458
rect 21824 16176 21876 16182
rect 21824 16118 21876 16124
rect 21928 15162 21956 19178
rect 22204 18766 22232 19382
rect 22192 18760 22244 18766
rect 22192 18702 22244 18708
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22112 18290 22140 18566
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 22008 17604 22060 17610
rect 22008 17546 22060 17552
rect 22192 17604 22244 17610
rect 22192 17546 22244 17552
rect 22020 17338 22048 17546
rect 22008 17332 22060 17338
rect 22008 17274 22060 17280
rect 22100 16992 22152 16998
rect 22100 16934 22152 16940
rect 22112 16454 22140 16934
rect 22100 16448 22152 16454
rect 22100 16390 22152 16396
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21548 14000 21600 14006
rect 21548 13942 21600 13948
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21456 9648 21508 9654
rect 21456 9590 21508 9596
rect 21456 8832 21508 8838
rect 21456 8774 21508 8780
rect 21468 5710 21496 8774
rect 21560 6798 21588 13262
rect 21640 13184 21692 13190
rect 21640 13126 21692 13132
rect 21652 9194 21680 13126
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21744 12102 21772 12378
rect 21732 12096 21784 12102
rect 21732 12038 21784 12044
rect 21836 11801 21864 14214
rect 22020 12714 22048 14962
rect 22112 12850 22140 16390
rect 22204 15008 22232 17546
rect 22296 16522 22324 20334
rect 22388 16590 22416 22086
rect 22480 21536 22508 25638
rect 22572 21690 22600 26454
rect 22664 24750 22692 26846
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 22744 26376 22796 26382
rect 22744 26318 22796 26324
rect 22652 24744 22704 24750
rect 22652 24686 22704 24692
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 22480 21508 22600 21536
rect 22468 21412 22520 21418
rect 22468 21354 22520 21360
rect 22480 20466 22508 21354
rect 22468 20460 22520 20466
rect 22468 20402 22520 20408
rect 22572 17218 22600 21508
rect 22756 20534 22784 26318
rect 22836 25764 22888 25770
rect 22836 25706 22888 25712
rect 22744 20528 22796 20534
rect 22744 20470 22796 20476
rect 22848 20346 22876 25706
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 23308 24818 23336 26930
rect 23400 26382 23428 29718
rect 23480 28008 23532 28014
rect 23480 27950 23532 27956
rect 23492 27606 23520 27950
rect 23480 27600 23532 27606
rect 23480 27542 23532 27548
rect 23584 27418 23612 30126
rect 24124 29300 24176 29306
rect 24124 29242 24176 29248
rect 23756 29096 23808 29102
rect 23756 29038 23808 29044
rect 23768 28762 23796 29038
rect 23756 28756 23808 28762
rect 23756 28698 23808 28704
rect 23664 28620 23716 28626
rect 23664 28562 23716 28568
rect 23676 27674 23704 28562
rect 23664 27668 23716 27674
rect 23664 27610 23716 27616
rect 23492 27390 23612 27418
rect 23664 27396 23716 27402
rect 23492 26926 23520 27390
rect 23664 27338 23716 27344
rect 23480 26920 23532 26926
rect 23480 26862 23532 26868
rect 23388 26376 23440 26382
rect 23388 26318 23440 26324
rect 23676 26296 23704 27338
rect 23584 26268 23704 26296
rect 23388 25832 23440 25838
rect 23388 25774 23440 25780
rect 23296 24812 23348 24818
rect 23296 24754 23348 24760
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 23308 24342 23336 24754
rect 23296 24336 23348 24342
rect 23296 24278 23348 24284
rect 23308 23746 23336 24278
rect 23400 23798 23428 25774
rect 23584 24682 23612 26268
rect 23768 26234 23796 28698
rect 23940 28416 23992 28422
rect 23940 28358 23992 28364
rect 23952 28014 23980 28358
rect 23940 28008 23992 28014
rect 23940 27950 23992 27956
rect 23952 27470 23980 27950
rect 24030 27704 24086 27713
rect 24030 27639 24086 27648
rect 23940 27464 23992 27470
rect 23940 27406 23992 27412
rect 24044 26382 24072 27639
rect 24136 27538 24164 29242
rect 24124 27532 24176 27538
rect 24124 27474 24176 27480
rect 24032 26376 24084 26382
rect 24032 26318 24084 26324
rect 23676 26206 23796 26234
rect 23572 24676 23624 24682
rect 23572 24618 23624 24624
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23216 23730 23336 23746
rect 23388 23792 23440 23798
rect 23388 23734 23440 23740
rect 23204 23724 23336 23730
rect 23256 23718 23336 23724
rect 23204 23666 23256 23672
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23296 22568 23348 22574
rect 23296 22510 23348 22516
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23204 22160 23256 22166
rect 23204 22102 23256 22108
rect 23216 21894 23244 22102
rect 23308 22001 23336 22510
rect 23400 22234 23428 23734
rect 23584 23662 23612 24006
rect 23572 23656 23624 23662
rect 23572 23598 23624 23604
rect 23388 22228 23440 22234
rect 23388 22170 23440 22176
rect 23294 21992 23350 22001
rect 23294 21927 23350 21936
rect 23204 21888 23256 21894
rect 23204 21830 23256 21836
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 22664 20318 22876 20346
rect 22664 18358 22692 20318
rect 22744 20256 22796 20262
rect 22744 20198 22796 20204
rect 22756 18766 22784 20198
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22652 18352 22704 18358
rect 22652 18294 22704 18300
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 22836 17672 22888 17678
rect 22836 17614 22888 17620
rect 22480 17190 22600 17218
rect 22376 16584 22428 16590
rect 22376 16526 22428 16532
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 22376 16448 22428 16454
rect 22376 16390 22428 16396
rect 22388 16046 22416 16390
rect 22376 16040 22428 16046
rect 22376 15982 22428 15988
rect 22284 15904 22336 15910
rect 22284 15846 22336 15852
rect 22296 15570 22324 15846
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22204 14980 22416 15008
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22008 12708 22060 12714
rect 22008 12650 22060 12656
rect 21916 12640 21968 12646
rect 21916 12582 21968 12588
rect 22100 12640 22152 12646
rect 22100 12582 22152 12588
rect 21822 11792 21878 11801
rect 21822 11727 21878 11736
rect 21732 11620 21784 11626
rect 21732 11562 21784 11568
rect 21744 11150 21772 11562
rect 21824 11348 21876 11354
rect 21824 11290 21876 11296
rect 21836 11150 21864 11290
rect 21732 11144 21784 11150
rect 21732 11086 21784 11092
rect 21824 11144 21876 11150
rect 21824 11086 21876 11092
rect 21824 10464 21876 10470
rect 21824 10406 21876 10412
rect 21836 10044 21864 10406
rect 21928 10112 21956 12582
rect 22112 12458 22140 12582
rect 22020 12430 22140 12458
rect 22020 12170 22048 12430
rect 22008 12164 22060 12170
rect 22008 12106 22060 12112
rect 22020 12050 22048 12106
rect 22020 12022 22140 12050
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 22020 10266 22048 10746
rect 22112 10470 22140 12022
rect 22204 10538 22232 12786
rect 22296 11558 22324 14758
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 22296 11150 22324 11494
rect 22284 11144 22336 11150
rect 22284 11086 22336 11092
rect 22192 10532 22244 10538
rect 22192 10474 22244 10480
rect 22100 10464 22152 10470
rect 22100 10406 22152 10412
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 22008 10124 22060 10130
rect 21928 10084 22008 10112
rect 22008 10066 22060 10072
rect 22112 10062 22140 10406
rect 22100 10056 22152 10062
rect 21836 10016 21956 10044
rect 21652 9166 21772 9194
rect 21640 7812 21692 7818
rect 21640 7754 21692 7760
rect 21548 6792 21600 6798
rect 21548 6734 21600 6740
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21560 5302 21588 5850
rect 21548 5296 21600 5302
rect 21548 5238 21600 5244
rect 21548 5160 21600 5166
rect 21548 5102 21600 5108
rect 21456 3936 21508 3942
rect 21456 3878 21508 3884
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 21364 2984 21416 2990
rect 21364 2926 21416 2932
rect 21178 2408 21234 2417
rect 21178 2343 21234 2352
rect 21192 2310 21220 2343
rect 21180 2304 21232 2310
rect 21180 2246 21232 2252
rect 20916 870 21036 898
rect 20916 762 20944 870
rect 21008 800 21036 870
rect 21376 800 21404 2926
rect 21468 2446 21496 3878
rect 21560 3738 21588 5102
rect 21548 3732 21600 3738
rect 21548 3674 21600 3680
rect 21652 3466 21680 7754
rect 21744 6798 21772 9166
rect 21824 8016 21876 8022
rect 21824 7958 21876 7964
rect 21836 7886 21864 7958
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 21928 7410 21956 10016
rect 22100 9998 22152 10004
rect 22388 9674 22416 14980
rect 22480 14550 22508 17190
rect 22560 17128 22612 17134
rect 22560 17070 22612 17076
rect 22468 14544 22520 14550
rect 22468 14486 22520 14492
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22480 12646 22508 12786
rect 22572 12714 22600 17070
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22664 13870 22692 16526
rect 22848 16454 22876 17614
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23020 15700 23072 15706
rect 23308 15688 23336 21830
rect 23584 21350 23612 23598
rect 23572 21344 23624 21350
rect 23572 21286 23624 21292
rect 23388 20528 23440 20534
rect 23388 20470 23440 20476
rect 23400 19718 23428 20470
rect 23572 20392 23624 20398
rect 23572 20334 23624 20340
rect 23480 20324 23532 20330
rect 23480 20266 23532 20272
rect 23388 19712 23440 19718
rect 23388 19654 23440 19660
rect 23400 18698 23428 19654
rect 23388 18692 23440 18698
rect 23388 18634 23440 18640
rect 23492 18290 23520 20266
rect 23584 19446 23612 20334
rect 23572 19440 23624 19446
rect 23572 19382 23624 19388
rect 23480 18284 23532 18290
rect 23480 18226 23532 18232
rect 23584 17592 23612 19382
rect 23492 17564 23612 17592
rect 23492 17202 23520 17564
rect 23676 17270 23704 26206
rect 23940 25900 23992 25906
rect 23940 25842 23992 25848
rect 23952 25498 23980 25842
rect 24044 25498 24072 26318
rect 23940 25492 23992 25498
rect 23940 25434 23992 25440
rect 24032 25492 24084 25498
rect 24032 25434 24084 25440
rect 23848 25220 23900 25226
rect 23848 25162 23900 25168
rect 23860 24449 23888 25162
rect 24124 24880 24176 24886
rect 24124 24822 24176 24828
rect 23846 24440 23902 24449
rect 23846 24375 23902 24384
rect 24136 24274 24164 24822
rect 24124 24268 24176 24274
rect 24124 24210 24176 24216
rect 23940 23520 23992 23526
rect 23940 23462 23992 23468
rect 23756 23112 23808 23118
rect 23756 23054 23808 23060
rect 23768 22234 23796 23054
rect 23952 22642 23980 23462
rect 23940 22636 23992 22642
rect 23940 22578 23992 22584
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 24228 22094 24256 43046
rect 24308 42560 24360 42566
rect 24308 42502 24360 42508
rect 24044 22066 24256 22094
rect 23940 20936 23992 20942
rect 23940 20878 23992 20884
rect 23952 20058 23980 20878
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 23846 19544 23902 19553
rect 23846 19479 23902 19488
rect 23860 18834 23888 19479
rect 23952 19446 23980 19994
rect 23940 19440 23992 19446
rect 23940 19382 23992 19388
rect 23848 18828 23900 18834
rect 23848 18770 23900 18776
rect 24044 17882 24072 22066
rect 24216 21684 24268 21690
rect 24216 21626 24268 21632
rect 24124 21616 24176 21622
rect 24228 21570 24256 21626
rect 24176 21564 24256 21570
rect 24124 21558 24256 21564
rect 24136 21542 24256 21558
rect 24136 20534 24164 21542
rect 24124 20528 24176 20534
rect 24124 20470 24176 20476
rect 24136 19786 24164 20470
rect 24124 19780 24176 19786
rect 24124 19722 24176 19728
rect 24136 19446 24164 19722
rect 24124 19440 24176 19446
rect 24124 19382 24176 19388
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 23756 17536 23808 17542
rect 23756 17478 23808 17484
rect 23664 17264 23716 17270
rect 23664 17206 23716 17212
rect 23480 17196 23532 17202
rect 23480 17138 23532 17144
rect 23386 17096 23442 17105
rect 23386 17031 23442 17040
rect 23400 16590 23428 17031
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 23492 15994 23520 17138
rect 23572 16108 23624 16114
rect 23572 16050 23624 16056
rect 23400 15966 23520 15994
rect 23400 15910 23428 15966
rect 23388 15904 23440 15910
rect 23388 15846 23440 15852
rect 23020 15642 23072 15648
rect 23216 15660 23336 15688
rect 23032 15434 23060 15642
rect 23020 15428 23072 15434
rect 23020 15370 23072 15376
rect 23216 15094 23244 15660
rect 23294 15464 23350 15473
rect 23294 15399 23350 15408
rect 23308 15094 23336 15399
rect 23204 15088 23256 15094
rect 23204 15030 23256 15036
rect 23296 15088 23348 15094
rect 23296 15030 23348 15036
rect 22744 14952 22796 14958
rect 22744 14894 22796 14900
rect 22652 13864 22704 13870
rect 22652 13806 22704 13812
rect 22560 12708 22612 12714
rect 22560 12650 22612 12656
rect 22468 12640 22520 12646
rect 22468 12582 22520 12588
rect 22650 12472 22706 12481
rect 22650 12407 22706 12416
rect 22468 12368 22520 12374
rect 22468 12310 22520 12316
rect 22480 10690 22508 12310
rect 22560 11280 22612 11286
rect 22560 11222 22612 11228
rect 22572 10849 22600 11222
rect 22558 10840 22614 10849
rect 22558 10775 22614 10784
rect 22480 10662 22600 10690
rect 22664 10674 22692 12407
rect 22468 10600 22520 10606
rect 22468 10542 22520 10548
rect 22020 9646 22416 9674
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 22020 7154 22048 9646
rect 22100 9580 22152 9586
rect 22100 9522 22152 9528
rect 22112 7886 22140 9522
rect 22480 9382 22508 10542
rect 22468 9376 22520 9382
rect 22388 9324 22468 9330
rect 22388 9318 22520 9324
rect 22388 9302 22508 9318
rect 22192 8492 22244 8498
rect 22192 8434 22244 8440
rect 22100 7880 22152 7886
rect 22100 7822 22152 7828
rect 21836 7126 22048 7154
rect 21732 6792 21784 6798
rect 21732 6734 21784 6740
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 21640 3460 21692 3466
rect 21640 3402 21692 3408
rect 21456 2440 21508 2446
rect 21456 2382 21508 2388
rect 21744 800 21772 6190
rect 21836 4622 21864 7126
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 21928 5914 21956 6734
rect 22008 6316 22060 6322
rect 22112 6304 22140 7822
rect 22060 6276 22140 6304
rect 22008 6258 22060 6264
rect 22008 6180 22060 6186
rect 22008 6122 22060 6128
rect 21916 5908 21968 5914
rect 21916 5850 21968 5856
rect 22020 5846 22048 6122
rect 22008 5840 22060 5846
rect 22008 5782 22060 5788
rect 21916 5364 21968 5370
rect 21916 5306 21968 5312
rect 21824 4616 21876 4622
rect 21824 4558 21876 4564
rect 21822 4312 21878 4321
rect 21822 4247 21878 4256
rect 21836 4146 21864 4247
rect 21824 4140 21876 4146
rect 21824 4082 21876 4088
rect 21928 4078 21956 5306
rect 22008 5228 22060 5234
rect 22008 5170 22060 5176
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 22020 4622 22048 5170
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 21916 4072 21968 4078
rect 21916 4014 21968 4020
rect 21916 3936 21968 3942
rect 21916 3878 21968 3884
rect 21928 3126 21956 3878
rect 22020 3210 22048 4082
rect 22112 3942 22140 5170
rect 22100 3936 22152 3942
rect 22100 3878 22152 3884
rect 22098 3224 22154 3233
rect 22020 3182 22098 3210
rect 22204 3194 22232 8434
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22098 3159 22154 3168
rect 22192 3188 22244 3194
rect 22112 3126 22140 3159
rect 22192 3130 22244 3136
rect 21916 3120 21968 3126
rect 21916 3062 21968 3068
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 21836 2774 21864 2994
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 21836 2746 22048 2774
rect 22020 2258 22048 2746
rect 22112 2514 22140 2858
rect 22296 2650 22324 8366
rect 22388 7954 22416 9302
rect 22468 8424 22520 8430
rect 22468 8366 22520 8372
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22388 4826 22416 7686
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 22284 2644 22336 2650
rect 22284 2586 22336 2592
rect 22192 2576 22244 2582
rect 22192 2518 22244 2524
rect 22100 2508 22152 2514
rect 22100 2450 22152 2456
rect 22020 2230 22140 2258
rect 22112 800 22140 2230
rect 22204 1601 22232 2518
rect 22190 1592 22246 1601
rect 22190 1527 22246 1536
rect 22480 800 22508 8366
rect 22572 8294 22600 10662
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 22664 9586 22692 10610
rect 22756 10062 22784 14894
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 23296 14476 23348 14482
rect 23296 14418 23348 14424
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 23204 13864 23256 13870
rect 23308 13818 23336 14418
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 23256 13812 23336 13818
rect 23204 13806 23336 13812
rect 22848 13394 22876 13806
rect 23216 13790 23336 13806
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22836 13388 22888 13394
rect 22836 13330 22888 13336
rect 22848 12850 22876 13330
rect 23308 12918 23336 13790
rect 23400 13258 23428 14010
rect 23388 13252 23440 13258
rect 23388 13194 23440 13200
rect 23296 12912 23348 12918
rect 23296 12854 23348 12860
rect 22836 12844 22888 12850
rect 22836 12786 22888 12792
rect 22848 12753 22876 12786
rect 22834 12744 22890 12753
rect 22834 12679 22890 12688
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 23388 12640 23440 12646
rect 23584 12628 23612 16050
rect 23768 15994 23796 17478
rect 24320 17218 24348 42502
rect 24504 42090 24532 52838
rect 24952 52420 25004 52426
rect 24952 52362 25004 52368
rect 24964 52193 24992 52362
rect 24950 52184 25006 52193
rect 25056 52154 25084 52935
rect 24950 52119 25006 52128
rect 25044 52148 25096 52154
rect 25044 52090 25096 52096
rect 25332 52018 25360 53926
rect 25872 53440 25924 53446
rect 25872 53382 25924 53388
rect 25320 52012 25372 52018
rect 25320 51954 25372 51960
rect 24950 51368 25006 51377
rect 24950 51303 24952 51312
rect 25004 51303 25006 51312
rect 24952 51274 25004 51280
rect 24952 50924 25004 50930
rect 24952 50866 25004 50872
rect 24964 50561 24992 50866
rect 24950 50552 25006 50561
rect 24950 50487 25006 50496
rect 25504 50176 25556 50182
rect 25504 50118 25556 50124
rect 25516 49842 25544 50118
rect 25504 49836 25556 49842
rect 25504 49778 25556 49784
rect 24676 49768 24728 49774
rect 25516 49745 25544 49778
rect 24676 49710 24728 49716
rect 25502 49736 25558 49745
rect 24492 42084 24544 42090
rect 24492 42026 24544 42032
rect 24688 41478 24716 49710
rect 25502 49671 25558 49680
rect 25136 49156 25188 49162
rect 25136 49098 25188 49104
rect 25148 48929 25176 49098
rect 25134 48920 25190 48929
rect 25134 48855 25190 48864
rect 25136 48544 25188 48550
rect 25136 48486 25188 48492
rect 25148 48142 25176 48486
rect 25136 48136 25188 48142
rect 25134 48104 25136 48113
rect 25188 48104 25190 48113
rect 25134 48039 25190 48048
rect 25320 47660 25372 47666
rect 25320 47602 25372 47608
rect 24952 47456 25004 47462
rect 24952 47398 25004 47404
rect 24768 44396 24820 44402
rect 24768 44338 24820 44344
rect 24780 44033 24808 44338
rect 24858 44296 24914 44305
rect 24858 44231 24914 44240
rect 24872 44198 24900 44231
rect 24860 44192 24912 44198
rect 24860 44134 24912 44140
rect 24766 44024 24822 44033
rect 24766 43959 24822 43968
rect 24676 41472 24728 41478
rect 24676 41414 24728 41420
rect 24676 33312 24728 33318
rect 24676 33254 24728 33260
rect 24768 33312 24820 33318
rect 24768 33254 24820 33260
rect 24688 32842 24716 33254
rect 24676 32836 24728 32842
rect 24676 32778 24728 32784
rect 24688 30410 24716 32778
rect 24780 32609 24808 33254
rect 24964 32910 24992 47398
rect 25332 47297 25360 47602
rect 25318 47288 25374 47297
rect 25318 47223 25374 47232
rect 25320 46912 25372 46918
rect 25320 46854 25372 46860
rect 25332 46578 25360 46854
rect 25320 46572 25372 46578
rect 25320 46514 25372 46520
rect 25332 46481 25360 46514
rect 25318 46472 25374 46481
rect 25318 46407 25374 46416
rect 25688 46368 25740 46374
rect 25688 46310 25740 46316
rect 25320 45960 25372 45966
rect 25320 45902 25372 45908
rect 25332 45665 25360 45902
rect 25318 45656 25374 45665
rect 25318 45591 25374 45600
rect 25320 45280 25372 45286
rect 25320 45222 25372 45228
rect 25332 44878 25360 45222
rect 25320 44872 25372 44878
rect 25318 44840 25320 44849
rect 25372 44840 25374 44849
rect 25318 44775 25374 44784
rect 25228 44736 25280 44742
rect 25228 44678 25280 44684
rect 25136 42628 25188 42634
rect 25136 42570 25188 42576
rect 25148 42401 25176 42570
rect 25134 42392 25190 42401
rect 25134 42327 25190 42336
rect 25136 42016 25188 42022
rect 25136 41958 25188 41964
rect 25148 41614 25176 41958
rect 25136 41608 25188 41614
rect 25134 41576 25136 41585
rect 25188 41576 25190 41585
rect 25134 41511 25190 41520
rect 25044 40928 25096 40934
rect 25044 40870 25096 40876
rect 25056 32978 25084 40870
rect 25136 37868 25188 37874
rect 25136 37810 25188 37816
rect 25148 37505 25176 37810
rect 25134 37496 25190 37505
rect 25134 37431 25190 37440
rect 25136 36032 25188 36038
rect 25136 35974 25188 35980
rect 25044 32972 25096 32978
rect 25044 32914 25096 32920
rect 24952 32904 25004 32910
rect 24952 32846 25004 32852
rect 24860 32768 24912 32774
rect 24860 32710 24912 32716
rect 24766 32600 24822 32609
rect 24872 32586 24900 32710
rect 24872 32558 24992 32586
rect 24766 32535 24822 32544
rect 24768 32496 24820 32502
rect 24768 32438 24820 32444
rect 24780 31686 24808 32438
rect 24768 31680 24820 31686
rect 24768 31622 24820 31628
rect 24780 31142 24808 31622
rect 24768 31136 24820 31142
rect 24768 31078 24820 31084
rect 24596 30382 24716 30410
rect 24492 29640 24544 29646
rect 24492 29582 24544 29588
rect 24504 29510 24532 29582
rect 24492 29504 24544 29510
rect 24492 29446 24544 29452
rect 24504 28529 24532 29446
rect 24596 29306 24624 30382
rect 24780 30274 24808 31078
rect 24860 30320 24912 30326
rect 24780 30268 24860 30274
rect 24780 30262 24912 30268
rect 24780 30246 24900 30262
rect 24872 30054 24900 30246
rect 24860 30048 24912 30054
rect 24860 29990 24912 29996
rect 24860 29572 24912 29578
rect 24860 29514 24912 29520
rect 24872 29345 24900 29514
rect 24858 29336 24914 29345
rect 24584 29300 24636 29306
rect 24858 29271 24914 29280
rect 24584 29242 24636 29248
rect 24964 29186 24992 32558
rect 25044 31952 25096 31958
rect 25044 31894 25096 31900
rect 24872 29158 24992 29186
rect 24676 29028 24728 29034
rect 24676 28970 24728 28976
rect 24490 28520 24546 28529
rect 24490 28455 24546 28464
rect 24400 28416 24452 28422
rect 24400 28358 24452 28364
rect 24412 18902 24440 28358
rect 24688 23066 24716 28970
rect 24768 28688 24820 28694
rect 24768 28630 24820 28636
rect 24780 28506 24808 28630
rect 24872 28626 24900 29158
rect 24952 29096 25004 29102
rect 24952 29038 25004 29044
rect 24860 28620 24912 28626
rect 24860 28562 24912 28568
rect 24964 28558 24992 29038
rect 24952 28552 25004 28558
rect 24780 28478 24900 28506
rect 24952 28494 25004 28500
rect 24768 27600 24820 27606
rect 24768 27542 24820 27548
rect 24780 27130 24808 27542
rect 24768 27124 24820 27130
rect 24768 27066 24820 27072
rect 24872 26790 24900 28478
rect 25056 27538 25084 31894
rect 25148 31278 25176 35974
rect 25240 35086 25268 44678
rect 25504 43648 25556 43654
rect 25504 43590 25556 43596
rect 25516 43382 25544 43590
rect 25504 43376 25556 43382
rect 25504 43318 25556 43324
rect 25516 43217 25544 43318
rect 25502 43208 25558 43217
rect 25502 43143 25558 43152
rect 25320 41132 25372 41138
rect 25320 41074 25372 41080
rect 25332 40769 25360 41074
rect 25318 40760 25374 40769
rect 25318 40695 25374 40704
rect 25504 40384 25556 40390
rect 25504 40326 25556 40332
rect 25516 40118 25544 40326
rect 25504 40112 25556 40118
rect 25504 40054 25556 40060
rect 25516 39953 25544 40054
rect 25502 39944 25558 39953
rect 25502 39879 25558 39888
rect 25320 39432 25372 39438
rect 25320 39374 25372 39380
rect 25332 39137 25360 39374
rect 25318 39128 25374 39137
rect 25318 39063 25374 39072
rect 25320 38752 25372 38758
rect 25320 38694 25372 38700
rect 25332 38350 25360 38694
rect 25320 38344 25372 38350
rect 25318 38312 25320 38321
rect 25372 38312 25374 38321
rect 25318 38247 25374 38256
rect 25412 38208 25464 38214
rect 25412 38150 25464 38156
rect 25320 36168 25372 36174
rect 25320 36110 25372 36116
rect 25332 35873 25360 36110
rect 25424 35894 25452 38150
rect 25504 37120 25556 37126
rect 25504 37062 25556 37068
rect 25516 36854 25544 37062
rect 25504 36848 25556 36854
rect 25504 36790 25556 36796
rect 25516 36689 25544 36790
rect 25502 36680 25558 36689
rect 25502 36615 25558 36624
rect 25596 36644 25648 36650
rect 25596 36586 25648 36592
rect 25318 35864 25374 35873
rect 25424 35866 25544 35894
rect 25318 35799 25374 35808
rect 25320 35488 25372 35494
rect 25320 35430 25372 35436
rect 25332 35086 25360 35430
rect 25228 35080 25280 35086
rect 25320 35080 25372 35086
rect 25228 35022 25280 35028
rect 25318 35048 25320 35057
rect 25372 35048 25374 35057
rect 25318 34983 25374 34992
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25332 34241 25360 34546
rect 25318 34232 25374 34241
rect 25318 34167 25374 34176
rect 25320 33992 25372 33998
rect 25320 33934 25372 33940
rect 25332 33425 25360 33934
rect 25318 33416 25374 33425
rect 25318 33351 25374 33360
rect 25320 33040 25372 33046
rect 25320 32982 25372 32988
rect 25228 32972 25280 32978
rect 25228 32914 25280 32920
rect 25240 32366 25268 32914
rect 25332 32570 25360 32982
rect 25412 32904 25464 32910
rect 25412 32846 25464 32852
rect 25320 32564 25372 32570
rect 25320 32506 25372 32512
rect 25228 32360 25280 32366
rect 25228 32302 25280 32308
rect 25136 31272 25188 31278
rect 25136 31214 25188 31220
rect 25136 31136 25188 31142
rect 25136 31078 25188 31084
rect 25044 27532 25096 27538
rect 25044 27474 25096 27480
rect 24860 26784 24912 26790
rect 24860 26726 24912 26732
rect 24872 26382 24900 26726
rect 24952 26580 25004 26586
rect 24952 26522 25004 26528
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 24858 26072 24914 26081
rect 24858 26007 24914 26016
rect 24872 25974 24900 26007
rect 24860 25968 24912 25974
rect 24860 25910 24912 25916
rect 24872 25430 24900 25910
rect 24860 25424 24912 25430
rect 24860 25366 24912 25372
rect 24964 24970 24992 26522
rect 25044 26512 25096 26518
rect 25044 26454 25096 26460
rect 24872 24942 24992 24970
rect 24766 23624 24822 23633
rect 24766 23559 24822 23568
rect 24504 23038 24716 23066
rect 24400 18896 24452 18902
rect 24400 18838 24452 18844
rect 24504 17338 24532 23038
rect 24584 22976 24636 22982
rect 24584 22918 24636 22924
rect 24596 19514 24624 22918
rect 24780 22574 24808 23559
rect 24768 22568 24820 22574
rect 24768 22510 24820 22516
rect 24872 21298 24900 24942
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 24964 23730 24992 24006
rect 24952 23724 25004 23730
rect 24952 23666 25004 23672
rect 24964 21690 24992 23666
rect 25056 22098 25084 26454
rect 25148 26450 25176 31078
rect 25240 30190 25268 32302
rect 25320 31816 25372 31822
rect 25318 31784 25320 31793
rect 25372 31784 25374 31793
rect 25318 31719 25374 31728
rect 25228 30184 25280 30190
rect 25228 30126 25280 30132
rect 25318 30152 25374 30161
rect 25318 30087 25374 30096
rect 25228 30048 25280 30054
rect 25228 29990 25280 29996
rect 25240 29510 25268 29990
rect 25332 29646 25360 30087
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 25228 29504 25280 29510
rect 25228 29446 25280 29452
rect 25240 27878 25268 29446
rect 25332 29306 25360 29582
rect 25320 29300 25372 29306
rect 25320 29242 25372 29248
rect 25424 29170 25452 32846
rect 25516 31482 25544 35866
rect 25504 31476 25556 31482
rect 25504 31418 25556 31424
rect 25504 31340 25556 31346
rect 25504 31282 25556 31288
rect 25516 30977 25544 31282
rect 25502 30968 25558 30977
rect 25502 30903 25504 30912
rect 25556 30903 25558 30912
rect 25504 30874 25556 30880
rect 25608 30818 25636 36586
rect 25700 35766 25728 46310
rect 25780 37732 25832 37738
rect 25780 37674 25832 37680
rect 25688 35760 25740 35766
rect 25688 35702 25740 35708
rect 25688 34944 25740 34950
rect 25688 34886 25740 34892
rect 25516 30790 25636 30818
rect 25412 29164 25464 29170
rect 25412 29106 25464 29112
rect 25228 27872 25280 27878
rect 25228 27814 25280 27820
rect 25412 27872 25464 27878
rect 25412 27814 25464 27820
rect 25240 27062 25268 27814
rect 25424 27470 25452 27814
rect 25412 27464 25464 27470
rect 25412 27406 25464 27412
rect 25228 27056 25280 27062
rect 25228 26998 25280 27004
rect 25318 26888 25374 26897
rect 25318 26823 25374 26832
rect 25136 26444 25188 26450
rect 25136 26386 25188 26392
rect 25228 26444 25280 26450
rect 25228 26386 25280 26392
rect 25136 26308 25188 26314
rect 25136 26250 25188 26256
rect 25148 26042 25176 26250
rect 25136 26036 25188 26042
rect 25136 25978 25188 25984
rect 25136 25832 25188 25838
rect 25136 25774 25188 25780
rect 25148 25265 25176 25774
rect 25134 25256 25190 25265
rect 25134 25191 25190 25200
rect 25136 25152 25188 25158
rect 25136 25094 25188 25100
rect 25148 24886 25176 25094
rect 25136 24880 25188 24886
rect 25136 24822 25188 24828
rect 25136 24744 25188 24750
rect 25240 24698 25268 26386
rect 25332 25294 25360 26823
rect 25424 26450 25452 27406
rect 25412 26444 25464 26450
rect 25412 26386 25464 26392
rect 25410 26344 25466 26353
rect 25410 26279 25466 26288
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25188 24692 25268 24698
rect 25136 24686 25268 24692
rect 25148 24670 25268 24686
rect 25148 23866 25176 24670
rect 25228 24608 25280 24614
rect 25228 24550 25280 24556
rect 25136 23860 25188 23866
rect 25136 23802 25188 23808
rect 25240 22234 25268 24550
rect 25332 24410 25360 25230
rect 25424 24614 25452 26279
rect 25412 24608 25464 24614
rect 25412 24550 25464 24556
rect 25320 24404 25372 24410
rect 25320 24346 25372 24352
rect 25412 24336 25464 24342
rect 25412 24278 25464 24284
rect 25424 23866 25452 24278
rect 25412 23860 25464 23866
rect 25412 23802 25464 23808
rect 25320 23180 25372 23186
rect 25320 23122 25372 23128
rect 25228 22228 25280 22234
rect 25228 22170 25280 22176
rect 25044 22092 25096 22098
rect 25044 22034 25096 22040
rect 24952 21684 25004 21690
rect 24952 21626 25004 21632
rect 25332 21486 25360 23122
rect 25424 23118 25452 23802
rect 25412 23112 25464 23118
rect 25412 23054 25464 23060
rect 25320 21480 25372 21486
rect 25320 21422 25372 21428
rect 25044 21344 25096 21350
rect 24872 21270 24992 21298
rect 25044 21286 25096 21292
rect 24858 21176 24914 21185
rect 24858 21111 24914 21120
rect 24872 21010 24900 21111
rect 24964 21010 24992 21270
rect 25056 21146 25084 21286
rect 25044 21140 25096 21146
rect 25044 21082 25096 21088
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 24674 20360 24730 20369
rect 24674 20295 24730 20304
rect 24584 19508 24636 19514
rect 24584 19450 24636 19456
rect 24688 18222 24716 20295
rect 24872 18850 24900 20742
rect 24964 19718 24992 20742
rect 25332 20602 25360 21422
rect 25320 20596 25372 20602
rect 25320 20538 25372 20544
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 24952 19712 25004 19718
rect 24952 19654 25004 19660
rect 25148 19514 25176 20334
rect 25412 19780 25464 19786
rect 25412 19722 25464 19728
rect 25424 19514 25452 19722
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 25412 19508 25464 19514
rect 25412 19450 25464 19456
rect 24872 18822 24992 18850
rect 24858 18728 24914 18737
rect 24858 18663 24914 18672
rect 24872 18358 24900 18663
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 24676 18216 24728 18222
rect 24676 18158 24728 18164
rect 24858 17912 24914 17921
rect 24858 17847 24914 17856
rect 24872 17746 24900 17847
rect 24964 17746 24992 18822
rect 25148 17746 25176 19450
rect 25228 18692 25280 18698
rect 25228 18634 25280 18640
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24952 17740 25004 17746
rect 24952 17682 25004 17688
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 25044 17604 25096 17610
rect 25044 17546 25096 17552
rect 24676 17536 24728 17542
rect 24676 17478 24728 17484
rect 24492 17332 24544 17338
rect 24492 17274 24544 17280
rect 24320 17190 24440 17218
rect 23848 16516 23900 16522
rect 23848 16458 23900 16464
rect 24216 16516 24268 16522
rect 24216 16458 24268 16464
rect 23388 12582 23440 12588
rect 23492 12600 23612 12628
rect 23676 15966 23796 15994
rect 22848 12374 22876 12582
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22836 12368 22888 12374
rect 22836 12310 22888 12316
rect 23296 11552 23348 11558
rect 23296 11494 23348 11500
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23308 11336 23336 11494
rect 23216 11308 23336 11336
rect 23216 10452 23244 11308
rect 23296 11212 23348 11218
rect 23296 11154 23348 11160
rect 23308 10577 23336 11154
rect 23400 10742 23428 12582
rect 23388 10736 23440 10742
rect 23388 10678 23440 10684
rect 23294 10568 23350 10577
rect 23294 10503 23350 10512
rect 23388 10464 23440 10470
rect 23216 10424 23336 10452
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 22652 9580 22704 9586
rect 22652 9522 22704 9528
rect 22652 9444 22704 9450
rect 22704 9404 22784 9432
rect 22652 9386 22704 9392
rect 22650 9072 22706 9081
rect 22650 9007 22706 9016
rect 22664 8974 22692 9007
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22560 8288 22612 8294
rect 22560 8230 22612 8236
rect 22652 6452 22704 6458
rect 22652 6394 22704 6400
rect 22560 6384 22612 6390
rect 22560 6326 22612 6332
rect 22572 5137 22600 6326
rect 22558 5128 22614 5137
rect 22558 5063 22614 5072
rect 22560 4004 22612 4010
rect 22560 3946 22612 3952
rect 22572 3194 22600 3946
rect 22664 3738 22692 6394
rect 22756 5710 22784 9404
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22836 7200 22888 7206
rect 22836 7142 22888 7148
rect 22848 6882 22876 7142
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22848 6854 22968 6882
rect 23308 6866 23336 10424
rect 23388 10406 23440 10412
rect 23400 10130 23428 10406
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23400 9518 23428 10066
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 22940 6338 22968 6854
rect 23296 6860 23348 6866
rect 23296 6802 23348 6808
rect 23400 6769 23428 7686
rect 23492 7546 23520 12600
rect 23572 12164 23624 12170
rect 23572 12106 23624 12112
rect 23584 11354 23612 12106
rect 23572 11348 23624 11354
rect 23572 11290 23624 11296
rect 23676 10810 23704 15966
rect 23756 15904 23808 15910
rect 23756 15846 23808 15852
rect 23768 15570 23796 15846
rect 23756 15564 23808 15570
rect 23756 15506 23808 15512
rect 23860 15552 23888 16458
rect 24228 15910 24256 16458
rect 24216 15904 24268 15910
rect 24216 15846 24268 15852
rect 23940 15564 23992 15570
rect 23860 15524 23940 15552
rect 23754 13832 23810 13841
rect 23754 13767 23810 13776
rect 23768 13394 23796 13767
rect 23860 13734 23888 15524
rect 23940 15506 23992 15512
rect 24228 15366 24256 15846
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 24216 15360 24268 15366
rect 24216 15302 24268 15308
rect 23848 13728 23900 13734
rect 23848 13670 23900 13676
rect 23756 13388 23808 13394
rect 23756 13330 23808 13336
rect 23756 11756 23808 11762
rect 23756 11698 23808 11704
rect 23664 10804 23716 10810
rect 23664 10746 23716 10752
rect 23664 8560 23716 8566
rect 23664 8502 23716 8508
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 23478 7440 23534 7449
rect 23478 7375 23480 7384
rect 23532 7375 23534 7384
rect 23480 7346 23532 7352
rect 23572 7268 23624 7274
rect 23572 7210 23624 7216
rect 23386 6760 23442 6769
rect 23386 6695 23442 6704
rect 23296 6656 23348 6662
rect 23296 6598 23348 6604
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 22848 6310 22968 6338
rect 22744 5704 22796 5710
rect 22744 5646 22796 5652
rect 22742 3904 22798 3913
rect 22742 3839 22798 3848
rect 22652 3732 22704 3738
rect 22652 3674 22704 3680
rect 22756 3602 22784 3839
rect 22848 3618 22876 6310
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 23308 5681 23336 6598
rect 23400 6474 23428 6598
rect 23400 6446 23520 6474
rect 23492 6202 23520 6446
rect 23400 6174 23520 6202
rect 23294 5672 23350 5681
rect 23294 5607 23350 5616
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 23400 4706 23428 6174
rect 23480 5160 23532 5166
rect 23480 5102 23532 5108
rect 23308 4678 23428 4706
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22744 3596 22796 3602
rect 22848 3590 22968 3618
rect 22744 3538 22796 3544
rect 22836 3460 22888 3466
rect 22836 3402 22888 3408
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 22848 800 22876 3402
rect 22940 3058 22968 3590
rect 23020 3460 23072 3466
rect 23020 3402 23072 3408
rect 23032 3126 23060 3402
rect 23112 3392 23164 3398
rect 23112 3334 23164 3340
rect 23124 3233 23152 3334
rect 23110 3224 23166 3233
rect 23110 3159 23166 3168
rect 23020 3120 23072 3126
rect 23020 3062 23072 3068
rect 22928 3052 22980 3058
rect 22928 2994 22980 3000
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 23204 2644 23256 2650
rect 23204 2586 23256 2592
rect 23216 800 23244 2586
rect 23308 2310 23336 4678
rect 23386 3632 23442 3641
rect 23386 3567 23442 3576
rect 23400 2774 23428 3567
rect 23492 2990 23520 5102
rect 23584 3126 23612 7210
rect 23676 3194 23704 8502
rect 23768 6458 23796 11698
rect 23952 11150 23980 15302
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 23940 11144 23992 11150
rect 23940 11086 23992 11092
rect 24044 9674 24072 14554
rect 24136 12442 24164 14962
rect 24228 13938 24256 15302
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24228 13818 24256 13874
rect 24228 13790 24348 13818
rect 24216 13456 24268 13462
rect 24216 13398 24268 13404
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 24122 10840 24178 10849
rect 24122 10775 24178 10784
rect 23952 9646 24072 9674
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23860 6934 23888 7686
rect 23848 6928 23900 6934
rect 23848 6870 23900 6876
rect 23756 6452 23808 6458
rect 23756 6394 23808 6400
rect 23860 6254 23888 6870
rect 23848 6248 23900 6254
rect 23848 6190 23900 6196
rect 23848 6112 23900 6118
rect 23848 6054 23900 6060
rect 23860 5710 23888 6054
rect 23952 5710 23980 9646
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 24044 8838 24072 9522
rect 24032 8832 24084 8838
rect 24032 8774 24084 8780
rect 24044 7886 24072 8774
rect 24032 7880 24084 7886
rect 24032 7822 24084 7828
rect 24032 6860 24084 6866
rect 24032 6802 24084 6808
rect 23848 5704 23900 5710
rect 23848 5646 23900 5652
rect 23940 5704 23992 5710
rect 23940 5646 23992 5652
rect 23756 5636 23808 5642
rect 23756 5578 23808 5584
rect 23768 5234 23796 5578
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 24044 4758 24072 6802
rect 24136 6322 24164 10775
rect 24228 8974 24256 13398
rect 24320 13190 24348 13790
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 24320 12986 24348 13126
rect 24308 12980 24360 12986
rect 24308 12922 24360 12928
rect 24320 10554 24348 12922
rect 24412 11898 24440 17190
rect 24584 16040 24636 16046
rect 24584 15982 24636 15988
rect 24492 14408 24544 14414
rect 24492 14350 24544 14356
rect 24504 13530 24532 14350
rect 24492 13524 24544 13530
rect 24492 13466 24544 13472
rect 24492 12232 24544 12238
rect 24492 12174 24544 12180
rect 24400 11892 24452 11898
rect 24400 11834 24452 11840
rect 24504 11014 24532 12174
rect 24492 11008 24544 11014
rect 24492 10950 24544 10956
rect 24320 10538 24440 10554
rect 24320 10532 24452 10538
rect 24320 10526 24400 10532
rect 24400 10474 24452 10480
rect 24412 9518 24440 10474
rect 24596 10266 24624 15982
rect 24688 15570 24716 17478
rect 24860 17196 24912 17202
rect 24860 17138 24912 17144
rect 24768 16584 24820 16590
rect 24768 16526 24820 16532
rect 24780 16250 24808 16526
rect 24872 16522 24900 17138
rect 24860 16516 24912 16522
rect 24860 16458 24912 16464
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24858 14648 24914 14657
rect 24858 14583 24914 14592
rect 24872 14482 24900 14583
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 25056 14414 25084 17546
rect 25134 16280 25190 16289
rect 25134 16215 25190 16224
rect 25148 15094 25176 16215
rect 25136 15088 25188 15094
rect 25136 15030 25188 15036
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 24860 14272 24912 14278
rect 24860 14214 24912 14220
rect 24766 13016 24822 13025
rect 24766 12951 24822 12960
rect 24780 11694 24808 12951
rect 24872 11914 24900 14214
rect 25044 13728 25096 13734
rect 25044 13670 25096 13676
rect 25056 13394 25084 13670
rect 25044 13388 25096 13394
rect 25044 13330 25096 13336
rect 24950 12200 25006 12209
rect 24950 12135 24952 12144
rect 25004 12135 25006 12144
rect 24952 12106 25004 12112
rect 24872 11886 24992 11914
rect 24860 11824 24912 11830
rect 24860 11766 24912 11772
rect 24768 11688 24820 11694
rect 24768 11630 24820 11636
rect 24872 11393 24900 11766
rect 24964 11762 24992 11886
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24858 11384 24914 11393
rect 24858 11319 24914 11328
rect 25044 11076 25096 11082
rect 25044 11018 25096 11024
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24492 10192 24544 10198
rect 24492 10134 24544 10140
rect 24400 9512 24452 9518
rect 24400 9454 24452 9460
rect 24216 8968 24268 8974
rect 24216 8910 24268 8916
rect 24216 7880 24268 7886
rect 24216 7822 24268 7828
rect 24228 7750 24256 7822
rect 24216 7744 24268 7750
rect 24216 7686 24268 7692
rect 24124 6316 24176 6322
rect 24124 6258 24176 6264
rect 24228 6202 24256 7686
rect 24504 6866 24532 10134
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24584 8832 24636 8838
rect 24584 8774 24636 8780
rect 24492 6860 24544 6866
rect 24492 6802 24544 6808
rect 24136 6174 24256 6202
rect 24136 6118 24164 6174
rect 24124 6112 24176 6118
rect 24124 6054 24176 6060
rect 24032 4752 24084 4758
rect 24032 4694 24084 4700
rect 23756 4480 23808 4486
rect 23756 4422 23808 4428
rect 23768 4185 23796 4422
rect 23754 4176 23810 4185
rect 23754 4111 23810 4120
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 23768 3466 23796 3878
rect 24044 3534 24072 4694
rect 24136 4078 24164 6054
rect 24596 5710 24624 8774
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 24584 5568 24636 5574
rect 24584 5510 24636 5516
rect 24216 5092 24268 5098
rect 24216 5034 24268 5040
rect 24124 4072 24176 4078
rect 24124 4014 24176 4020
rect 24032 3528 24084 3534
rect 23938 3496 23994 3505
rect 23756 3460 23808 3466
rect 24032 3470 24084 3476
rect 23938 3431 23994 3440
rect 23756 3402 23808 3408
rect 23664 3188 23716 3194
rect 23664 3130 23716 3136
rect 23572 3120 23624 3126
rect 23756 3120 23808 3126
rect 23572 3062 23624 3068
rect 23754 3088 23756 3097
rect 23808 3088 23810 3097
rect 23754 3023 23810 3032
rect 23480 2984 23532 2990
rect 23480 2926 23532 2932
rect 23400 2746 23612 2774
rect 23296 2304 23348 2310
rect 23296 2246 23348 2252
rect 23584 800 23612 2746
rect 23952 800 23980 3431
rect 24228 3194 24256 5034
rect 24596 3534 24624 5510
rect 24688 4282 24716 9862
rect 24766 9752 24822 9761
rect 24766 9687 24822 9696
rect 24780 8430 24808 9687
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24872 9110 24900 9318
rect 24860 9104 24912 9110
rect 24860 9046 24912 9052
rect 24950 8936 25006 8945
rect 24950 8871 24952 8880
rect 25004 8871 25006 8880
rect 24952 8842 25004 8848
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 25056 8022 25084 11018
rect 25134 8120 25190 8129
rect 25134 8055 25190 8064
rect 25044 8016 25096 8022
rect 25044 7958 25096 7964
rect 25148 7478 25176 8055
rect 25136 7472 25188 7478
rect 25136 7414 25188 7420
rect 24860 7336 24912 7342
rect 24858 7304 24860 7313
rect 24912 7304 24914 7313
rect 24858 7239 24914 7248
rect 25136 6724 25188 6730
rect 25136 6666 25188 6672
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24676 4276 24728 4282
rect 24676 4218 24728 4224
rect 24308 3528 24360 3534
rect 24308 3470 24360 3476
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24216 3188 24268 3194
rect 24216 3130 24268 3136
rect 24320 800 24348 3470
rect 24584 3392 24636 3398
rect 24584 3334 24636 3340
rect 24596 2446 24624 3334
rect 24872 2514 24900 6598
rect 25148 6497 25176 6666
rect 25134 6488 25190 6497
rect 25134 6423 25190 6432
rect 25240 5914 25268 18634
rect 25516 11286 25544 30790
rect 25596 26920 25648 26926
rect 25596 26862 25648 26868
rect 25608 26489 25636 26862
rect 25594 26480 25650 26489
rect 25594 26415 25650 26424
rect 25596 26308 25648 26314
rect 25596 26250 25648 26256
rect 25608 18970 25636 26250
rect 25596 18964 25648 18970
rect 25596 18906 25648 18912
rect 25700 17814 25728 34886
rect 25688 17808 25740 17814
rect 25688 17750 25740 17756
rect 25792 11626 25820 37674
rect 25884 33402 25912 53382
rect 26516 52488 26568 52494
rect 26516 52430 26568 52436
rect 26056 45824 26108 45830
rect 26056 45766 26108 45772
rect 26068 35834 26096 45766
rect 26056 35828 26108 35834
rect 26056 35770 26108 35776
rect 26240 33856 26292 33862
rect 26240 33798 26292 33804
rect 25884 33374 26188 33402
rect 25964 33312 26016 33318
rect 25964 33254 26016 33260
rect 25872 31272 25924 31278
rect 25872 31214 25924 31220
rect 25884 26382 25912 31214
rect 25976 28490 26004 33254
rect 26056 32564 26108 32570
rect 26056 32506 26108 32512
rect 26068 28626 26096 32506
rect 26160 30122 26188 33374
rect 26148 30116 26200 30122
rect 26148 30058 26200 30064
rect 26148 29844 26200 29850
rect 26148 29786 26200 29792
rect 26056 28620 26108 28626
rect 26056 28562 26108 28568
rect 25964 28484 26016 28490
rect 25964 28426 26016 28432
rect 25964 26784 26016 26790
rect 25964 26726 26016 26732
rect 25872 26376 25924 26382
rect 25872 26318 25924 26324
rect 25870 26248 25926 26257
rect 25870 26183 25926 26192
rect 25884 23254 25912 26183
rect 25976 24342 26004 26726
rect 26160 26353 26188 29786
rect 26252 28218 26280 33798
rect 26528 32230 26556 52430
rect 26608 51332 26660 51338
rect 26608 51274 26660 51280
rect 26516 32224 26568 32230
rect 26516 32166 26568 32172
rect 26620 29714 26648 51274
rect 26608 29708 26660 29714
rect 26608 29650 26660 29656
rect 26240 28212 26292 28218
rect 26240 28154 26292 28160
rect 26240 27056 26292 27062
rect 26240 26998 26292 27004
rect 26146 26344 26202 26353
rect 26146 26279 26202 26288
rect 26252 26234 26280 26998
rect 26068 26206 26280 26234
rect 26068 25226 26096 26206
rect 26056 25220 26108 25226
rect 26056 25162 26108 25168
rect 26068 24410 26096 25162
rect 26056 24404 26108 24410
rect 26056 24346 26108 24352
rect 25964 24336 26016 24342
rect 25964 24278 26016 24284
rect 26068 23798 26096 24346
rect 26056 23792 26108 23798
rect 26056 23734 26108 23740
rect 25872 23248 25924 23254
rect 25872 23190 25924 23196
rect 25872 23044 25924 23050
rect 25872 22986 25924 22992
rect 25884 22817 25912 22986
rect 25870 22808 25926 22817
rect 25870 22743 25926 22752
rect 25780 11620 25832 11626
rect 25780 11562 25832 11568
rect 25504 11280 25556 11286
rect 25504 11222 25556 11228
rect 25320 8084 25372 8090
rect 25320 8026 25372 8032
rect 25228 5908 25280 5914
rect 25228 5850 25280 5856
rect 25136 5636 25188 5642
rect 25136 5578 25188 5584
rect 25148 3058 25176 5578
rect 25136 3052 25188 3058
rect 25136 2994 25188 3000
rect 24950 2952 25006 2961
rect 24950 2887 24952 2896
rect 25004 2887 25006 2896
rect 24952 2858 25004 2864
rect 25240 2774 25268 5850
rect 25148 2746 25268 2774
rect 24860 2508 24912 2514
rect 24860 2450 24912 2456
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 25148 2378 25176 2746
rect 25136 2372 25188 2378
rect 25136 2314 25188 2320
rect 25228 2304 25280 2310
rect 25228 2246 25280 2252
rect 25240 1834 25268 2246
rect 25228 1828 25280 1834
rect 25228 1770 25280 1776
rect 20732 734 20944 762
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25332 785 25360 8026
rect 25318 776 25374 785
rect 25318 711 25374 720
<< via2 >>
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 2778 8744 2834 8800
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 3422 6432 3478 6488
rect 3422 4120 3478 4176
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 3514 1808 3570 1864
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 23386 56072 23442 56128
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 9954 18128 10010 18184
rect 8758 12824 8814 12880
rect 5446 2508 5502 2544
rect 5446 2488 5448 2508
rect 5448 2488 5500 2508
rect 5500 2488 5502 2508
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 10230 14476 10286 14512
rect 10230 14456 10232 14476
rect 10232 14456 10284 14476
rect 10284 14456 10286 14476
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 10138 8880 10194 8936
rect 10598 5208 10654 5264
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 11794 12688 11850 12744
rect 11518 8336 11574 8392
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12622 12688 12678 12744
rect 12530 10512 12586 10568
rect 12162 9968 12218 10024
rect 11886 9868 11888 9888
rect 11888 9868 11940 9888
rect 11940 9868 11942 9888
rect 11886 9832 11942 9868
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 13910 18128 13966 18184
rect 14186 18164 14188 18184
rect 14188 18164 14240 18184
rect 14240 18164 14242 18184
rect 14186 18128 14242 18164
rect 13082 12688 13138 12744
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 13450 11892 13506 11928
rect 13450 11872 13452 11892
rect 13452 11872 13504 11892
rect 13504 11872 13506 11892
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12714 10804 12770 10840
rect 12714 10784 12716 10804
rect 12716 10784 12768 10804
rect 12768 10784 12770 10804
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12714 9832 12770 9888
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 13450 10104 13506 10160
rect 13910 14220 13912 14240
rect 13912 14220 13964 14240
rect 13964 14220 13966 14240
rect 13910 14184 13966 14220
rect 12530 7384 12586 7440
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12254 3984 12310 4040
rect 12622 3576 12678 3632
rect 14370 14456 14426 14512
rect 14002 10648 14058 10704
rect 14646 12824 14702 12880
rect 14370 12008 14426 12064
rect 13818 8472 13874 8528
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 13542 6704 13598 6760
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 14278 10784 14334 10840
rect 14278 9016 14334 9072
rect 14186 6316 14242 6352
rect 14186 6296 14188 6316
rect 14188 6296 14240 6316
rect 14240 6296 14242 6316
rect 14462 10548 14464 10568
rect 14464 10548 14516 10568
rect 14516 10548 14518 10568
rect 14462 10512 14518 10548
rect 15658 24792 15714 24848
rect 15474 20712 15530 20768
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 14646 7928 14702 7984
rect 15474 12844 15530 12880
rect 15474 12824 15476 12844
rect 15476 12824 15528 12844
rect 15528 12824 15530 12844
rect 14646 2896 14702 2952
rect 15106 7928 15162 7984
rect 15658 11872 15714 11928
rect 15934 12688 15990 12744
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 17130 23160 17186 23216
rect 16670 18672 16726 18728
rect 16578 13640 16634 13696
rect 16118 12008 16174 12064
rect 16026 11056 16082 11112
rect 15382 6296 15438 6352
rect 15198 5772 15254 5808
rect 15198 5752 15200 5772
rect 15200 5752 15252 5772
rect 15252 5752 15254 5772
rect 16946 17312 17002 17368
rect 16486 10548 16488 10568
rect 16488 10548 16540 10568
rect 16540 10548 16542 10568
rect 16486 10512 16542 10548
rect 17590 25064 17646 25120
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 17222 16224 17278 16280
rect 17314 15272 17370 15328
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17498 13504 17554 13560
rect 17038 10104 17094 10160
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18418 13640 18474 13696
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17222 8492 17278 8528
rect 17222 8472 17224 8492
rect 17224 8472 17276 8492
rect 17276 8472 17278 8492
rect 17498 3576 17554 3632
rect 18878 23432 18934 23488
rect 19062 22616 19118 22672
rect 18050 9968 18106 10024
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17958 8880 18014 8936
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18326 5208 18382 5264
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18786 10104 18842 10160
rect 18694 9968 18750 10024
rect 18786 9832 18842 9888
rect 18694 9424 18750 9480
rect 18878 9696 18934 9752
rect 18878 3848 18934 3904
rect 19522 22616 19578 22672
rect 19890 24928 19946 24984
rect 19430 12980 19486 13016
rect 19430 12960 19432 12980
rect 19432 12960 19484 12980
rect 19484 12960 19486 12980
rect 19062 8336 19118 8392
rect 19798 12960 19854 13016
rect 19246 5344 19302 5400
rect 19522 6976 19578 7032
rect 19982 10668 20038 10704
rect 19982 10648 19984 10668
rect 19984 10648 20036 10668
rect 20036 10648 20038 10668
rect 19706 6840 19762 6896
rect 19706 6568 19762 6624
rect 19706 4548 19762 4584
rect 19982 5752 20038 5808
rect 19706 4528 19708 4548
rect 19708 4528 19760 4548
rect 19760 4528 19762 4548
rect 21086 18028 21088 18048
rect 21088 18028 21140 18048
rect 21140 18028 21142 18048
rect 21086 17992 21142 18028
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 24766 55392 24822 55448
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 24490 54576 24546 54632
rect 25042 53760 25098 53816
rect 25042 52944 25098 53000
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 20810 11736 20866 11792
rect 20350 6296 20406 6352
rect 20442 5364 20498 5400
rect 20442 5344 20444 5364
rect 20444 5344 20496 5364
rect 20496 5344 20498 5364
rect 20718 6976 20774 7032
rect 20350 3168 20406 3224
rect 20534 3068 20536 3088
rect 20536 3068 20588 3088
rect 20588 3068 20590 3088
rect 20534 3032 20590 3068
rect 20994 6568 21050 6624
rect 21086 4256 21142 4312
rect 21178 3984 21234 4040
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 24030 27648 24086 27704
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 23294 21936 23350 21992
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 21822 11736 21878 11792
rect 21178 2352 21234 2408
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 23846 24384 23902 24440
rect 23846 19488 23902 19544
rect 23386 17040 23442 17096
rect 23294 15408 23350 15464
rect 22650 12416 22706 12472
rect 22558 10784 22614 10840
rect 21822 4256 21878 4312
rect 22098 3168 22154 3224
rect 22190 1536 22246 1592
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22834 12688 22890 12744
rect 24950 52128 25006 52184
rect 24950 51332 25006 51368
rect 24950 51312 24952 51332
rect 24952 51312 25004 51332
rect 25004 51312 25006 51332
rect 24950 50496 25006 50552
rect 25502 49680 25558 49736
rect 25134 48864 25190 48920
rect 25134 48084 25136 48104
rect 25136 48084 25188 48104
rect 25188 48084 25190 48104
rect 25134 48048 25190 48084
rect 24858 44240 24914 44296
rect 24766 43968 24822 44024
rect 25318 47232 25374 47288
rect 25318 46416 25374 46472
rect 25318 45600 25374 45656
rect 25318 44820 25320 44840
rect 25320 44820 25372 44840
rect 25372 44820 25374 44840
rect 25318 44784 25374 44820
rect 25134 42336 25190 42392
rect 25134 41556 25136 41576
rect 25136 41556 25188 41576
rect 25188 41556 25190 41576
rect 25134 41520 25190 41556
rect 25134 37440 25190 37496
rect 24766 32544 24822 32600
rect 24858 29280 24914 29336
rect 24490 28464 24546 28520
rect 25502 43152 25558 43208
rect 25318 40704 25374 40760
rect 25502 39888 25558 39944
rect 25318 39072 25374 39128
rect 25318 38292 25320 38312
rect 25320 38292 25372 38312
rect 25372 38292 25374 38312
rect 25318 38256 25374 38292
rect 25502 36624 25558 36680
rect 25318 35808 25374 35864
rect 25318 35028 25320 35048
rect 25320 35028 25372 35048
rect 25372 35028 25374 35048
rect 25318 34992 25374 35028
rect 25318 34176 25374 34232
rect 25318 33360 25374 33416
rect 24858 26016 24914 26072
rect 24766 23568 24822 23624
rect 25318 31764 25320 31784
rect 25320 31764 25372 31784
rect 25372 31764 25374 31784
rect 25318 31728 25374 31764
rect 25318 30096 25374 30152
rect 25502 30932 25558 30968
rect 25502 30912 25504 30932
rect 25504 30912 25556 30932
rect 25556 30912 25558 30932
rect 25318 26832 25374 26888
rect 25134 25200 25190 25256
rect 25410 26288 25466 26344
rect 24858 21120 24914 21176
rect 24674 20304 24730 20360
rect 24858 18672 24914 18728
rect 24858 17856 24914 17912
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 23294 10512 23350 10568
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22650 9016 22706 9072
rect 22558 5072 22614 5128
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 23754 13776 23810 13832
rect 23478 7404 23534 7440
rect 23478 7384 23480 7404
rect 23480 7384 23532 7404
rect 23532 7384 23534 7404
rect 23386 6704 23442 6760
rect 22742 3848 22798 3904
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 23294 5616 23350 5672
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 23110 3168 23166 3224
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 23386 3576 23442 3632
rect 24122 10784 24178 10840
rect 24858 14592 24914 14648
rect 25134 16224 25190 16280
rect 24766 12960 24822 13016
rect 24950 12164 25006 12200
rect 24950 12144 24952 12164
rect 24952 12144 25004 12164
rect 25004 12144 25006 12164
rect 24858 11328 24914 11384
rect 23754 4120 23810 4176
rect 23938 3440 23994 3496
rect 23754 3068 23756 3088
rect 23756 3068 23808 3088
rect 23808 3068 23810 3088
rect 23754 3032 23810 3068
rect 24766 9696 24822 9752
rect 24950 8900 25006 8936
rect 24950 8880 24952 8900
rect 24952 8880 25004 8900
rect 25004 8880 25006 8900
rect 25134 8064 25190 8120
rect 24858 7284 24860 7304
rect 24860 7284 24912 7304
rect 24912 7284 24914 7304
rect 24858 7248 24914 7284
rect 25134 6432 25190 6488
rect 25594 26424 25650 26480
rect 25870 26192 25926 26248
rect 26146 26288 26202 26344
rect 25870 22752 25926 22808
rect 24950 2916 25006 2952
rect 24950 2896 24952 2916
rect 24952 2896 25004 2916
rect 25004 2896 25006 2916
rect 25318 720 25374 776
<< metal3 >>
rect 26200 56266 27000 56296
rect 23430 56206 27000 56266
rect 23430 56133 23490 56206
rect 26200 56176 27000 56206
rect 23381 56128 23490 56133
rect 23381 56072 23386 56128
rect 23442 56072 23490 56128
rect 23381 56070 23490 56072
rect 23381 56067 23447 56070
rect 24761 55450 24827 55453
rect 26200 55450 27000 55480
rect 24761 55448 27000 55450
rect 24761 55392 24766 55448
rect 24822 55392 27000 55448
rect 24761 55390 27000 55392
rect 24761 55387 24827 55390
rect 26200 55360 27000 55390
rect 24485 54634 24551 54637
rect 26200 54634 27000 54664
rect 24485 54632 27000 54634
rect 24485 54576 24490 54632
rect 24546 54576 27000 54632
rect 24485 54574 27000 54576
rect 24485 54571 24551 54574
rect 26200 54544 27000 54574
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 25037 53818 25103 53821
rect 26200 53818 27000 53848
rect 25037 53816 27000 53818
rect 25037 53760 25042 53816
rect 25098 53760 27000 53816
rect 25037 53758 27000 53760
rect 25037 53755 25103 53758
rect 26200 53728 27000 53758
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 25037 53002 25103 53005
rect 26200 53002 27000 53032
rect 25037 53000 27000 53002
rect 25037 52944 25042 53000
rect 25098 52944 27000 53000
rect 25037 52942 27000 52944
rect 25037 52939 25103 52942
rect 26200 52912 27000 52942
rect 2946 52800 3262 52801
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 24945 52186 25011 52189
rect 26200 52186 27000 52216
rect 24945 52184 27000 52186
rect 24945 52128 24950 52184
rect 25006 52128 27000 52184
rect 24945 52126 27000 52128
rect 24945 52123 25011 52126
rect 26200 52096 27000 52126
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 24945 51370 25011 51373
rect 26200 51370 27000 51400
rect 24945 51368 27000 51370
rect 24945 51312 24950 51368
rect 25006 51312 27000 51368
rect 24945 51310 27000 51312
rect 24945 51307 25011 51310
rect 26200 51280 27000 51310
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 2946 50624 3262 50625
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 24945 50554 25011 50557
rect 26200 50554 27000 50584
rect 24945 50552 27000 50554
rect 24945 50496 24950 50552
rect 25006 50496 27000 50552
rect 24945 50494 27000 50496
rect 24945 50491 25011 50494
rect 26200 50464 27000 50494
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 25497 49738 25563 49741
rect 26200 49738 27000 49768
rect 25497 49736 27000 49738
rect 25497 49680 25502 49736
rect 25558 49680 27000 49736
rect 25497 49678 27000 49680
rect 25497 49675 25563 49678
rect 26200 49648 27000 49678
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 25129 48922 25195 48925
rect 26200 48922 27000 48952
rect 25129 48920 27000 48922
rect 25129 48864 25134 48920
rect 25190 48864 27000 48920
rect 25129 48862 27000 48864
rect 25129 48859 25195 48862
rect 26200 48832 27000 48862
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 25129 48106 25195 48109
rect 26200 48106 27000 48136
rect 25129 48104 27000 48106
rect 25129 48048 25134 48104
rect 25190 48048 27000 48104
rect 25129 48046 27000 48048
rect 25129 48043 25195 48046
rect 26200 48016 27000 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 25313 47290 25379 47293
rect 26200 47290 27000 47320
rect 25313 47288 27000 47290
rect 25313 47232 25318 47288
rect 25374 47232 27000 47288
rect 25313 47230 27000 47232
rect 25313 47227 25379 47230
rect 26200 47200 27000 47230
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 25313 46474 25379 46477
rect 26200 46474 27000 46504
rect 25313 46472 27000 46474
rect 25313 46416 25318 46472
rect 25374 46416 27000 46472
rect 25313 46414 27000 46416
rect 25313 46411 25379 46414
rect 26200 46384 27000 46414
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 7946 45728 8262 45729
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 25313 45658 25379 45661
rect 26200 45658 27000 45688
rect 25313 45656 27000 45658
rect 25313 45600 25318 45656
rect 25374 45600 27000 45656
rect 25313 45598 27000 45600
rect 25313 45595 25379 45598
rect 26200 45568 27000 45598
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 25313 44842 25379 44845
rect 26200 44842 27000 44872
rect 25313 44840 27000 44842
rect 25313 44784 25318 44840
rect 25374 44784 27000 44840
rect 25313 44782 27000 44784
rect 25313 44779 25379 44782
rect 26200 44752 27000 44782
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 21398 44236 21404 44300
rect 21468 44298 21474 44300
rect 24853 44298 24919 44301
rect 21468 44296 24919 44298
rect 21468 44240 24858 44296
rect 24914 44240 24919 44296
rect 21468 44238 24919 44240
rect 21468 44236 21474 44238
rect 24853 44235 24919 44238
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 24761 44026 24827 44029
rect 26200 44026 27000 44056
rect 24761 44024 27000 44026
rect 24761 43968 24766 44024
rect 24822 43968 27000 44024
rect 24761 43966 27000 43968
rect 24761 43963 24827 43966
rect 26200 43936 27000 43966
rect 7946 43552 8262 43553
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 25497 43210 25563 43213
rect 26200 43210 27000 43240
rect 25497 43208 27000 43210
rect 25497 43152 25502 43208
rect 25558 43152 27000 43208
rect 25497 43150 27000 43152
rect 25497 43147 25563 43150
rect 26200 43120 27000 43150
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 25129 42394 25195 42397
rect 26200 42394 27000 42424
rect 25129 42392 27000 42394
rect 25129 42336 25134 42392
rect 25190 42336 27000 42392
rect 25129 42334 27000 42336
rect 25129 42331 25195 42334
rect 26200 42304 27000 42334
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 25129 41578 25195 41581
rect 26200 41578 27000 41608
rect 25129 41576 27000 41578
rect 25129 41520 25134 41576
rect 25190 41520 27000 41576
rect 25129 41518 27000 41520
rect 25129 41515 25195 41518
rect 26200 41488 27000 41518
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 2946 40832 3262 40833
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 25313 40762 25379 40765
rect 26200 40762 27000 40792
rect 25313 40760 27000 40762
rect 25313 40704 25318 40760
rect 25374 40704 27000 40760
rect 25313 40702 27000 40704
rect 25313 40699 25379 40702
rect 26200 40672 27000 40702
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 25497 39946 25563 39949
rect 26200 39946 27000 39976
rect 25497 39944 27000 39946
rect 25497 39888 25502 39944
rect 25558 39888 27000 39944
rect 25497 39886 27000 39888
rect 25497 39883 25563 39886
rect 26200 39856 27000 39886
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 25313 39130 25379 39133
rect 26200 39130 27000 39160
rect 25313 39128 27000 39130
rect 25313 39072 25318 39128
rect 25374 39072 27000 39128
rect 25313 39070 27000 39072
rect 25313 39067 25379 39070
rect 26200 39040 27000 39070
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 25313 38314 25379 38317
rect 26200 38314 27000 38344
rect 25313 38312 27000 38314
rect 25313 38256 25318 38312
rect 25374 38256 27000 38312
rect 25313 38254 27000 38256
rect 25313 38251 25379 38254
rect 26200 38224 27000 38254
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 25129 37498 25195 37501
rect 26200 37498 27000 37528
rect 25129 37496 27000 37498
rect 25129 37440 25134 37496
rect 25190 37440 27000 37496
rect 25129 37438 27000 37440
rect 25129 37435 25195 37438
rect 26200 37408 27000 37438
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 25497 36682 25563 36685
rect 26200 36682 27000 36712
rect 25497 36680 27000 36682
rect 25497 36624 25502 36680
rect 25558 36624 27000 36680
rect 25497 36622 27000 36624
rect 25497 36619 25563 36622
rect 26200 36592 27000 36622
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 7946 35936 8262 35937
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 25313 35866 25379 35869
rect 26200 35866 27000 35896
rect 25313 35864 27000 35866
rect 25313 35808 25318 35864
rect 25374 35808 27000 35864
rect 25313 35806 27000 35808
rect 25313 35803 25379 35806
rect 26200 35776 27000 35806
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 25313 35050 25379 35053
rect 26200 35050 27000 35080
rect 25313 35048 27000 35050
rect 25313 34992 25318 35048
rect 25374 34992 27000 35048
rect 25313 34990 27000 34992
rect 25313 34987 25379 34990
rect 26200 34960 27000 34990
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 2946 34304 3262 34305
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 25313 34234 25379 34237
rect 26200 34234 27000 34264
rect 25313 34232 27000 34234
rect 25313 34176 25318 34232
rect 25374 34176 27000 34232
rect 25313 34174 27000 34176
rect 25313 34171 25379 34174
rect 26200 34144 27000 34174
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 25313 33418 25379 33421
rect 26200 33418 27000 33448
rect 25313 33416 27000 33418
rect 25313 33360 25318 33416
rect 25374 33360 27000 33416
rect 25313 33358 27000 33360
rect 25313 33355 25379 33358
rect 26200 33328 27000 33358
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 24761 32602 24827 32605
rect 26200 32602 27000 32632
rect 24761 32600 27000 32602
rect 24761 32544 24766 32600
rect 24822 32544 27000 32600
rect 24761 32542 27000 32544
rect 24761 32539 24827 32542
rect 26200 32512 27000 32542
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 25313 31786 25379 31789
rect 26200 31786 27000 31816
rect 25313 31784 27000 31786
rect 25313 31728 25318 31784
rect 25374 31728 27000 31784
rect 25313 31726 27000 31728
rect 25313 31723 25379 31726
rect 26200 31696 27000 31726
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 2946 31040 3262 31041
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 25497 30970 25563 30973
rect 26200 30970 27000 31000
rect 25497 30968 27000 30970
rect 25497 30912 25502 30968
rect 25558 30912 27000 30968
rect 25497 30910 27000 30912
rect 25497 30907 25563 30910
rect 26200 30880 27000 30910
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 25313 30154 25379 30157
rect 26200 30154 27000 30184
rect 25313 30152 27000 30154
rect 25313 30096 25318 30152
rect 25374 30096 27000 30152
rect 25313 30094 27000 30096
rect 25313 30091 25379 30094
rect 26200 30064 27000 30094
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 24853 29338 24919 29341
rect 26200 29338 27000 29368
rect 24853 29336 27000 29338
rect 24853 29280 24858 29336
rect 24914 29280 27000 29336
rect 24853 29278 27000 29280
rect 24853 29275 24919 29278
rect 26200 29248 27000 29278
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 24485 28522 24551 28525
rect 26200 28522 27000 28552
rect 24485 28520 27000 28522
rect 24485 28464 24490 28520
rect 24546 28464 27000 28520
rect 24485 28462 27000 28464
rect 24485 28459 24551 28462
rect 26200 28432 27000 28462
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 24025 27706 24091 27709
rect 26200 27706 27000 27736
rect 24025 27704 27000 27706
rect 24025 27648 24030 27704
rect 24086 27648 27000 27704
rect 24025 27646 27000 27648
rect 24025 27643 24091 27646
rect 26200 27616 27000 27646
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 25313 26890 25379 26893
rect 26200 26890 27000 26920
rect 25313 26888 27000 26890
rect 25313 26832 25318 26888
rect 25374 26832 27000 26888
rect 25313 26830 27000 26832
rect 25313 26827 25379 26830
rect 26200 26800 27000 26830
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 25589 26482 25655 26485
rect 25454 26480 25655 26482
rect 25454 26424 25594 26480
rect 25650 26424 25655 26480
rect 25454 26422 25655 26424
rect 25454 26349 25514 26422
rect 25589 26419 25655 26422
rect 25405 26344 25514 26349
rect 26141 26346 26207 26349
rect 25405 26288 25410 26344
rect 25466 26288 25514 26344
rect 25405 26286 25514 26288
rect 26006 26344 26207 26346
rect 26006 26288 26146 26344
rect 26202 26288 26207 26344
rect 26006 26286 26207 26288
rect 25405 26283 25471 26286
rect 25865 26250 25931 26253
rect 26006 26250 26066 26286
rect 26141 26283 26207 26286
rect 25865 26248 26066 26250
rect 25865 26192 25870 26248
rect 25926 26192 26066 26248
rect 25865 26190 26066 26192
rect 25865 26187 25931 26190
rect 7946 26144 8262 26145
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 24853 26074 24919 26077
rect 26200 26074 27000 26104
rect 24853 26072 27000 26074
rect 24853 26016 24858 26072
rect 24914 26016 27000 26072
rect 24853 26014 27000 26016
rect 24853 26011 24919 26014
rect 26200 25984 27000 26014
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 25129 25258 25195 25261
rect 26200 25258 27000 25288
rect 25129 25256 27000 25258
rect 25129 25200 25134 25256
rect 25190 25200 27000 25256
rect 25129 25198 27000 25200
rect 25129 25195 25195 25198
rect 26200 25168 27000 25198
rect 17166 25060 17172 25124
rect 17236 25122 17242 25124
rect 17585 25122 17651 25125
rect 17236 25120 17651 25122
rect 17236 25064 17590 25120
rect 17646 25064 17651 25120
rect 17236 25062 17651 25064
rect 17236 25060 17242 25062
rect 17585 25059 17651 25062
rect 7946 25056 8262 25057
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 19885 24988 19951 24989
rect 19885 24984 19932 24988
rect 19996 24986 20002 24988
rect 19885 24928 19890 24984
rect 19885 24924 19932 24928
rect 19996 24926 20042 24986
rect 19996 24924 20002 24926
rect 19885 24923 19951 24924
rect 15653 24850 15719 24853
rect 16430 24850 16436 24852
rect 15653 24848 16436 24850
rect 15653 24792 15658 24848
rect 15714 24792 16436 24848
rect 15653 24790 16436 24792
rect 15653 24787 15719 24790
rect 16430 24788 16436 24790
rect 16500 24788 16506 24852
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 23841 24442 23907 24445
rect 26200 24442 27000 24472
rect 23841 24440 27000 24442
rect 23841 24384 23846 24440
rect 23902 24384 27000 24440
rect 23841 24382 27000 24384
rect 23841 24379 23907 24382
rect 26200 24352 27000 24382
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 24761 23626 24827 23629
rect 26200 23626 27000 23656
rect 24761 23624 27000 23626
rect 24761 23568 24766 23624
rect 24822 23568 27000 23624
rect 24761 23566 27000 23568
rect 24761 23563 24827 23566
rect 26200 23536 27000 23566
rect 18873 23490 18939 23493
rect 19006 23490 19012 23492
rect 18873 23488 19012 23490
rect 18873 23432 18878 23488
rect 18934 23432 19012 23488
rect 18873 23430 19012 23432
rect 18873 23427 18939 23430
rect 19006 23428 19012 23430
rect 19076 23428 19082 23492
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 17125 23218 17191 23221
rect 17350 23218 17356 23220
rect 17125 23216 17356 23218
rect 17125 23160 17130 23216
rect 17186 23160 17356 23216
rect 17125 23158 17356 23160
rect 17125 23155 17191 23158
rect 17350 23156 17356 23158
rect 17420 23156 17426 23220
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 25865 22810 25931 22813
rect 26200 22810 27000 22840
rect 25865 22808 27000 22810
rect 25865 22752 25870 22808
rect 25926 22752 27000 22808
rect 25865 22750 27000 22752
rect 25865 22747 25931 22750
rect 26200 22720 27000 22750
rect 19057 22674 19123 22677
rect 19517 22674 19583 22677
rect 19057 22672 19583 22674
rect 19057 22616 19062 22672
rect 19118 22616 19522 22672
rect 19578 22616 19583 22672
rect 19057 22614 19583 22616
rect 19057 22611 19123 22614
rect 19517 22611 19583 22614
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 23289 21994 23355 21997
rect 26200 21994 27000 22024
rect 23289 21992 27000 21994
rect 23289 21936 23294 21992
rect 23350 21936 27000 21992
rect 23289 21934 27000 21936
rect 23289 21931 23355 21934
rect 26200 21904 27000 21934
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 24853 21178 24919 21181
rect 26200 21178 27000 21208
rect 24853 21176 27000 21178
rect 24853 21120 24858 21176
rect 24914 21120 27000 21176
rect 24853 21118 27000 21120
rect 24853 21115 24919 21118
rect 26200 21088 27000 21118
rect 14038 20708 14044 20772
rect 14108 20770 14114 20772
rect 15469 20770 15535 20773
rect 14108 20768 15535 20770
rect 14108 20712 15474 20768
rect 15530 20712 15535 20768
rect 14108 20710 15535 20712
rect 14108 20708 14114 20710
rect 15469 20707 15535 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 24669 20362 24735 20365
rect 26200 20362 27000 20392
rect 24669 20360 27000 20362
rect 24669 20304 24674 20360
rect 24730 20304 27000 20360
rect 24669 20302 27000 20304
rect 24669 20299 24735 20302
rect 26200 20272 27000 20302
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 23841 19546 23907 19549
rect 26200 19546 27000 19576
rect 23841 19544 27000 19546
rect 23841 19488 23846 19544
rect 23902 19488 27000 19544
rect 23841 19486 27000 19488
rect 23841 19483 23907 19486
rect 26200 19456 27000 19486
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 16665 18730 16731 18733
rect 17534 18730 17540 18732
rect 16665 18728 17540 18730
rect 16665 18672 16670 18728
rect 16726 18672 17540 18728
rect 16665 18670 17540 18672
rect 16665 18667 16731 18670
rect 17534 18668 17540 18670
rect 17604 18730 17610 18732
rect 21398 18730 21404 18732
rect 17604 18670 21404 18730
rect 17604 18668 17610 18670
rect 21398 18668 21404 18670
rect 21468 18668 21474 18732
rect 24853 18730 24919 18733
rect 26200 18730 27000 18760
rect 24853 18728 27000 18730
rect 24853 18672 24858 18728
rect 24914 18672 27000 18728
rect 24853 18670 27000 18672
rect 24853 18667 24919 18670
rect 26200 18640 27000 18670
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 9949 18186 10015 18189
rect 13905 18186 13971 18189
rect 14181 18186 14247 18189
rect 9949 18184 14247 18186
rect 9949 18128 9954 18184
rect 10010 18128 13910 18184
rect 13966 18128 14186 18184
rect 14242 18128 14247 18184
rect 9949 18126 14247 18128
rect 9949 18123 10015 18126
rect 13905 18123 13971 18126
rect 14181 18123 14247 18126
rect 21081 18050 21147 18053
rect 21214 18050 21220 18052
rect 21081 18048 21220 18050
rect 21081 17992 21086 18048
rect 21142 17992 21220 18048
rect 21081 17990 21220 17992
rect 21081 17987 21147 17990
rect 21214 17988 21220 17990
rect 21284 17988 21290 18052
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 24853 17914 24919 17917
rect 26200 17914 27000 17944
rect 24853 17912 27000 17914
rect 24853 17856 24858 17912
rect 24914 17856 27000 17912
rect 24853 17854 27000 17856
rect 24853 17851 24919 17854
rect 26200 17824 27000 17854
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 16941 17370 17007 17373
rect 17166 17370 17172 17372
rect 16941 17368 17172 17370
rect 16941 17312 16946 17368
rect 17002 17312 17172 17368
rect 16941 17310 17172 17312
rect 16941 17307 17007 17310
rect 17166 17308 17172 17310
rect 17236 17308 17242 17372
rect 23381 17098 23447 17101
rect 26200 17098 27000 17128
rect 23381 17096 27000 17098
rect 23381 17040 23386 17096
rect 23442 17040 27000 17096
rect 23381 17038 27000 17040
rect 23381 17035 23447 17038
rect 26200 17008 27000 17038
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 17217 16282 17283 16285
rect 17350 16282 17356 16284
rect 17217 16280 17356 16282
rect 17217 16224 17222 16280
rect 17278 16224 17356 16280
rect 17217 16222 17356 16224
rect 17217 16219 17283 16222
rect 17350 16220 17356 16222
rect 17420 16220 17426 16284
rect 25129 16282 25195 16285
rect 26200 16282 27000 16312
rect 25129 16280 27000 16282
rect 25129 16224 25134 16280
rect 25190 16224 27000 16280
rect 25129 16222 27000 16224
rect 25129 16219 25195 16222
rect 26200 16192 27000 16222
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 23289 15466 23355 15469
rect 26200 15466 27000 15496
rect 23289 15464 27000 15466
rect 23289 15408 23294 15464
rect 23350 15408 27000 15464
rect 23289 15406 27000 15408
rect 23289 15403 23355 15406
rect 26200 15376 27000 15406
rect 16982 15268 16988 15332
rect 17052 15330 17058 15332
rect 17309 15330 17375 15333
rect 17052 15328 17375 15330
rect 17052 15272 17314 15328
rect 17370 15272 17375 15328
rect 17052 15270 17375 15272
rect 17052 15268 17058 15270
rect 17309 15267 17375 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 24853 14650 24919 14653
rect 26200 14650 27000 14680
rect 24853 14648 27000 14650
rect 24853 14592 24858 14648
rect 24914 14592 27000 14648
rect 24853 14590 27000 14592
rect 24853 14587 24919 14590
rect 26200 14560 27000 14590
rect 10225 14514 10291 14517
rect 14365 14514 14431 14517
rect 10225 14512 14431 14514
rect 10225 14456 10230 14512
rect 10286 14456 14370 14512
rect 14426 14456 14431 14512
rect 10225 14454 14431 14456
rect 10225 14451 10291 14454
rect 14365 14451 14431 14454
rect 13905 14244 13971 14245
rect 13854 14180 13860 14244
rect 13924 14242 13971 14244
rect 13924 14240 14016 14242
rect 13966 14184 14016 14240
rect 13924 14182 14016 14184
rect 13924 14180 13971 14182
rect 13905 14179 13971 14180
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 23749 13834 23815 13837
rect 26200 13834 27000 13864
rect 23749 13832 27000 13834
rect 23749 13776 23754 13832
rect 23810 13776 27000 13832
rect 23749 13774 27000 13776
rect 23749 13771 23815 13774
rect 26200 13744 27000 13774
rect 16573 13698 16639 13701
rect 18413 13698 18479 13701
rect 16573 13696 18479 13698
rect 16573 13640 16578 13696
rect 16634 13640 18418 13696
rect 18474 13640 18479 13696
rect 16573 13638 18479 13640
rect 16573 13635 16639 13638
rect 18413 13635 18479 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 17493 13564 17559 13565
rect 17493 13562 17540 13564
rect 17448 13560 17540 13562
rect 17448 13504 17498 13560
rect 17448 13502 17540 13504
rect 17493 13500 17540 13502
rect 17604 13500 17610 13564
rect 17493 13499 17559 13500
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 19425 13018 19491 13021
rect 19793 13018 19859 13021
rect 19425 13016 19859 13018
rect 19425 12960 19430 13016
rect 19486 12960 19798 13016
rect 19854 12960 19859 13016
rect 19425 12958 19859 12960
rect 19425 12955 19491 12958
rect 19793 12955 19859 12958
rect 24761 13018 24827 13021
rect 26200 13018 27000 13048
rect 24761 13016 27000 13018
rect 24761 12960 24766 13016
rect 24822 12960 27000 13016
rect 24761 12958 27000 12960
rect 24761 12955 24827 12958
rect 26200 12928 27000 12958
rect 8753 12882 8819 12885
rect 14641 12882 14707 12885
rect 15469 12882 15535 12885
rect 8753 12880 15535 12882
rect 8753 12824 8758 12880
rect 8814 12824 14646 12880
rect 14702 12824 15474 12880
rect 15530 12824 15535 12880
rect 8753 12822 15535 12824
rect 8753 12819 8819 12822
rect 14641 12819 14707 12822
rect 15469 12819 15535 12822
rect 11789 12746 11855 12749
rect 12617 12746 12683 12749
rect 11789 12744 12683 12746
rect 11789 12688 11794 12744
rect 11850 12688 12622 12744
rect 12678 12688 12683 12744
rect 11789 12686 12683 12688
rect 11789 12683 11855 12686
rect 12617 12683 12683 12686
rect 13077 12746 13143 12749
rect 15929 12746 15995 12749
rect 22829 12746 22895 12749
rect 13077 12744 15995 12746
rect 13077 12688 13082 12744
rect 13138 12688 15934 12744
rect 15990 12688 15995 12744
rect 13077 12686 15995 12688
rect 13077 12683 13143 12686
rect 15929 12683 15995 12686
rect 22694 12744 22895 12746
rect 22694 12688 22834 12744
rect 22890 12688 22895 12744
rect 22694 12686 22895 12688
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22694 12477 22754 12686
rect 22829 12683 22895 12686
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 22645 12472 22754 12477
rect 22645 12416 22650 12472
rect 22706 12416 22754 12472
rect 22645 12414 22754 12416
rect 22645 12411 22711 12414
rect 24945 12202 25011 12205
rect 26200 12202 27000 12232
rect 24945 12200 27000 12202
rect 24945 12144 24950 12200
rect 25006 12144 27000 12200
rect 24945 12142 27000 12144
rect 24945 12139 25011 12142
rect 26200 12112 27000 12142
rect 14365 12066 14431 12069
rect 16113 12066 16179 12069
rect 14365 12064 16179 12066
rect 14365 12008 14370 12064
rect 14426 12008 16118 12064
rect 16174 12008 16179 12064
rect 14365 12006 16179 12008
rect 14365 12003 14431 12006
rect 16113 12003 16179 12006
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 13445 11930 13511 11933
rect 15653 11930 15719 11933
rect 13445 11928 15719 11930
rect 13445 11872 13450 11928
rect 13506 11872 15658 11928
rect 15714 11872 15719 11928
rect 13445 11870 15719 11872
rect 13445 11867 13511 11870
rect 15653 11867 15719 11870
rect 20805 11794 20871 11797
rect 21817 11794 21883 11797
rect 20805 11792 21883 11794
rect 20805 11736 20810 11792
rect 20866 11736 21822 11792
rect 21878 11736 21883 11792
rect 20805 11734 21883 11736
rect 20805 11731 20871 11734
rect 21817 11731 21883 11734
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 24853 11386 24919 11389
rect 26200 11386 27000 11416
rect 24853 11384 27000 11386
rect 24853 11328 24858 11384
rect 24914 11328 27000 11384
rect 24853 11326 27000 11328
rect 24853 11323 24919 11326
rect 26200 11296 27000 11326
rect 16021 11114 16087 11117
rect 16982 11114 16988 11116
rect 16021 11112 16988 11114
rect 16021 11056 16026 11112
rect 16082 11056 16988 11112
rect 16021 11054 16988 11056
rect 16021 11051 16087 11054
rect 16982 11052 16988 11054
rect 17052 11052 17058 11116
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 12709 10842 12775 10845
rect 14273 10842 14339 10845
rect 12709 10840 14339 10842
rect 12709 10784 12714 10840
rect 12770 10784 14278 10840
rect 14334 10784 14339 10840
rect 12709 10782 14339 10784
rect 12709 10779 12775 10782
rect 14273 10779 14339 10782
rect 22553 10842 22619 10845
rect 24117 10842 24183 10845
rect 22553 10840 24183 10842
rect 22553 10784 22558 10840
rect 22614 10784 24122 10840
rect 24178 10784 24183 10840
rect 22553 10782 24183 10784
rect 22553 10779 22619 10782
rect 24117 10779 24183 10782
rect 13997 10708 14063 10709
rect 13997 10706 14044 10708
rect 13956 10704 14044 10706
rect 14108 10706 14114 10708
rect 19977 10706 20043 10709
rect 14108 10704 20043 10706
rect 13956 10648 14002 10704
rect 14108 10648 19982 10704
rect 20038 10648 20043 10704
rect 13956 10646 14044 10648
rect 13997 10644 14044 10646
rect 14108 10646 20043 10648
rect 14108 10644 14114 10646
rect 13997 10643 14063 10644
rect 19977 10643 20043 10646
rect 12525 10570 12591 10573
rect 14457 10570 14523 10573
rect 16481 10570 16547 10573
rect 12525 10568 16547 10570
rect 12525 10512 12530 10568
rect 12586 10512 14462 10568
rect 14518 10512 16486 10568
rect 16542 10512 16547 10568
rect 12525 10510 16547 10512
rect 12525 10507 12591 10510
rect 14457 10507 14523 10510
rect 16481 10507 16547 10510
rect 23289 10570 23355 10573
rect 26200 10570 27000 10600
rect 23289 10568 27000 10570
rect 23289 10512 23294 10568
rect 23350 10512 27000 10568
rect 23289 10510 27000 10512
rect 23289 10507 23355 10510
rect 26200 10480 27000 10510
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 13445 10162 13511 10165
rect 17033 10162 17099 10165
rect 13445 10160 17099 10162
rect 13445 10104 13450 10160
rect 13506 10104 17038 10160
rect 17094 10104 17099 10160
rect 13445 10102 17099 10104
rect 13445 10099 13511 10102
rect 17033 10099 17099 10102
rect 18781 10162 18847 10165
rect 18781 10160 18890 10162
rect 18781 10104 18786 10160
rect 18842 10104 18890 10160
rect 18781 10099 18890 10104
rect 12157 10026 12223 10029
rect 18045 10026 18111 10029
rect 18689 10026 18755 10029
rect 12157 10024 18111 10026
rect 12157 9968 12162 10024
rect 12218 9968 18050 10024
rect 18106 9968 18111 10024
rect 12157 9966 18111 9968
rect 12157 9963 12223 9966
rect 18045 9963 18111 9966
rect 18646 10024 18755 10026
rect 18646 9968 18694 10024
rect 18750 9968 18755 10024
rect 18646 9963 18755 9968
rect 11881 9890 11947 9893
rect 12709 9890 12775 9893
rect 11881 9888 12775 9890
rect 11881 9832 11886 9888
rect 11942 9832 12714 9888
rect 12770 9832 12775 9888
rect 11881 9830 12775 9832
rect 11881 9827 11947 9830
rect 12709 9827 12775 9830
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 18646 9754 18706 9963
rect 18830 9893 18890 10099
rect 18781 9888 18890 9893
rect 18781 9832 18786 9888
rect 18842 9832 18890 9888
rect 18781 9830 18890 9832
rect 18781 9827 18847 9830
rect 18873 9754 18939 9757
rect 18646 9752 18939 9754
rect 18646 9696 18878 9752
rect 18934 9696 18939 9752
rect 18646 9694 18939 9696
rect 18873 9691 18939 9694
rect 24761 9754 24827 9757
rect 26200 9754 27000 9784
rect 24761 9752 27000 9754
rect 24761 9696 24766 9752
rect 24822 9696 27000 9752
rect 24761 9694 27000 9696
rect 24761 9691 24827 9694
rect 26200 9664 27000 9694
rect 18689 9482 18755 9485
rect 21214 9482 21220 9484
rect 18689 9480 21220 9482
rect 18689 9424 18694 9480
rect 18750 9424 21220 9480
rect 18689 9422 21220 9424
rect 18689 9419 18755 9422
rect 21214 9420 21220 9422
rect 21284 9420 21290 9484
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 14273 9074 14339 9077
rect 22645 9074 22711 9077
rect 14273 9072 22711 9074
rect 14273 9016 14278 9072
rect 14334 9016 22650 9072
rect 22706 9016 22711 9072
rect 14273 9014 22711 9016
rect 14273 9011 14339 9014
rect 22645 9011 22711 9014
rect 10133 8938 10199 8941
rect 17953 8938 18019 8941
rect 10133 8936 18019 8938
rect 10133 8880 10138 8936
rect 10194 8880 17958 8936
rect 18014 8880 18019 8936
rect 10133 8878 18019 8880
rect 10133 8875 10199 8878
rect 17953 8875 18019 8878
rect 24945 8938 25011 8941
rect 26200 8938 27000 8968
rect 24945 8936 27000 8938
rect 24945 8880 24950 8936
rect 25006 8880 27000 8936
rect 24945 8878 27000 8880
rect 24945 8875 25011 8878
rect 26200 8848 27000 8878
rect 0 8802 800 8832
rect 2773 8802 2839 8805
rect 0 8800 2839 8802
rect 0 8744 2778 8800
rect 2834 8744 2839 8800
rect 0 8742 2839 8744
rect 0 8712 800 8742
rect 2773 8739 2839 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 13813 8530 13879 8533
rect 17217 8530 17283 8533
rect 13813 8528 17283 8530
rect 13813 8472 13818 8528
rect 13874 8472 17222 8528
rect 17278 8472 17283 8528
rect 13813 8470 17283 8472
rect 13813 8467 13879 8470
rect 17217 8467 17283 8470
rect 11513 8394 11579 8397
rect 19057 8394 19123 8397
rect 11513 8392 19123 8394
rect 11513 8336 11518 8392
rect 11574 8336 19062 8392
rect 19118 8336 19123 8392
rect 11513 8334 19123 8336
rect 11513 8331 11579 8334
rect 19057 8331 19123 8334
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 25129 8122 25195 8125
rect 26200 8122 27000 8152
rect 25129 8120 27000 8122
rect 25129 8064 25134 8120
rect 25190 8064 27000 8120
rect 25129 8062 27000 8064
rect 25129 8059 25195 8062
rect 26200 8032 27000 8062
rect 14641 7986 14707 7989
rect 15101 7986 15167 7989
rect 14641 7984 15167 7986
rect 14641 7928 14646 7984
rect 14702 7928 15106 7984
rect 15162 7928 15167 7984
rect 14641 7926 15167 7928
rect 14641 7923 14707 7926
rect 15101 7923 15167 7926
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 12525 7442 12591 7445
rect 23473 7442 23539 7445
rect 12525 7440 23539 7442
rect 12525 7384 12530 7440
rect 12586 7384 23478 7440
rect 23534 7384 23539 7440
rect 12525 7382 23539 7384
rect 12525 7379 12591 7382
rect 23473 7379 23539 7382
rect 24853 7306 24919 7309
rect 26200 7306 27000 7336
rect 24853 7304 27000 7306
rect 24853 7248 24858 7304
rect 24914 7248 27000 7304
rect 24853 7246 27000 7248
rect 24853 7243 24919 7246
rect 26200 7216 27000 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 19517 7034 19583 7037
rect 20713 7034 20779 7037
rect 19517 7032 20779 7034
rect 19517 6976 19522 7032
rect 19578 6976 20718 7032
rect 20774 6976 20779 7032
rect 19517 6974 20779 6976
rect 19517 6971 19583 6974
rect 20713 6971 20779 6974
rect 19701 6900 19767 6901
rect 19701 6896 19748 6900
rect 19812 6898 19818 6900
rect 19701 6840 19706 6896
rect 19701 6836 19748 6840
rect 19812 6838 19858 6898
rect 19812 6836 19818 6838
rect 19701 6835 19767 6836
rect 13537 6762 13603 6765
rect 23381 6762 23447 6765
rect 13537 6760 23447 6762
rect 13537 6704 13542 6760
rect 13598 6704 23386 6760
rect 23442 6704 23447 6760
rect 13537 6702 23447 6704
rect 13537 6699 13603 6702
rect 23381 6699 23447 6702
rect 19701 6626 19767 6629
rect 20989 6626 21055 6629
rect 19701 6624 21055 6626
rect 19701 6568 19706 6624
rect 19762 6568 20994 6624
rect 21050 6568 21055 6624
rect 19701 6566 21055 6568
rect 19701 6563 19767 6566
rect 20989 6563 21055 6566
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 3417 6490 3483 6493
rect 0 6488 3483 6490
rect 0 6432 3422 6488
rect 3478 6432 3483 6488
rect 0 6430 3483 6432
rect 0 6400 800 6430
rect 3417 6427 3483 6430
rect 25129 6490 25195 6493
rect 26200 6490 27000 6520
rect 25129 6488 27000 6490
rect 25129 6432 25134 6488
rect 25190 6432 27000 6488
rect 25129 6430 27000 6432
rect 25129 6427 25195 6430
rect 26200 6400 27000 6430
rect 14038 6292 14044 6356
rect 14108 6354 14114 6356
rect 14181 6354 14247 6357
rect 14108 6352 14247 6354
rect 14108 6296 14186 6352
rect 14242 6296 14247 6352
rect 14108 6294 14247 6296
rect 14108 6292 14114 6294
rect 14181 6291 14247 6294
rect 15377 6354 15443 6357
rect 20345 6354 20411 6357
rect 15377 6352 20411 6354
rect 15377 6296 15382 6352
rect 15438 6296 20350 6352
rect 20406 6296 20411 6352
rect 15377 6294 20411 6296
rect 15377 6291 15443 6294
rect 20345 6291 20411 6294
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 15193 5810 15259 5813
rect 16430 5810 16436 5812
rect 15193 5808 16436 5810
rect 15193 5752 15198 5808
rect 15254 5752 16436 5808
rect 15193 5750 16436 5752
rect 15193 5747 15259 5750
rect 16430 5748 16436 5750
rect 16500 5810 16506 5812
rect 19977 5810 20043 5813
rect 16500 5808 20043 5810
rect 16500 5752 19982 5808
rect 20038 5752 20043 5808
rect 16500 5750 20043 5752
rect 16500 5748 16506 5750
rect 19977 5747 20043 5750
rect 23289 5674 23355 5677
rect 26200 5674 27000 5704
rect 23289 5672 27000 5674
rect 23289 5616 23294 5672
rect 23350 5616 27000 5672
rect 23289 5614 27000 5616
rect 23289 5611 23355 5614
rect 26200 5584 27000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 19241 5402 19307 5405
rect 20437 5402 20503 5405
rect 19241 5400 20503 5402
rect 19241 5344 19246 5400
rect 19302 5344 20442 5400
rect 20498 5344 20503 5400
rect 19241 5342 20503 5344
rect 19241 5339 19307 5342
rect 20437 5339 20503 5342
rect 10593 5266 10659 5269
rect 18321 5266 18387 5269
rect 10593 5264 18387 5266
rect 10593 5208 10598 5264
rect 10654 5208 18326 5264
rect 18382 5208 18387 5264
rect 10593 5206 18387 5208
rect 10593 5203 10659 5206
rect 18321 5203 18387 5206
rect 22553 5130 22619 5133
rect 22553 5128 23490 5130
rect 22553 5072 22558 5128
rect 22614 5072 23490 5128
rect 22553 5070 23490 5072
rect 22553 5067 22619 5070
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 23430 4858 23490 5070
rect 26200 4858 27000 4888
rect 23430 4798 27000 4858
rect 26200 4768 27000 4798
rect 19701 4588 19767 4589
rect 19701 4586 19748 4588
rect 19656 4584 19748 4586
rect 19656 4528 19706 4584
rect 19656 4526 19748 4528
rect 19701 4524 19748 4526
rect 19812 4524 19818 4588
rect 19701 4523 19767 4524
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 21081 4314 21147 4317
rect 21817 4314 21883 4317
rect 21081 4312 21883 4314
rect 21081 4256 21086 4312
rect 21142 4256 21822 4312
rect 21878 4256 21883 4312
rect 21081 4254 21883 4256
rect 21081 4251 21147 4254
rect 21817 4251 21883 4254
rect 0 4178 800 4208
rect 3417 4178 3483 4181
rect 23749 4178 23815 4181
rect 0 4176 3483 4178
rect 0 4120 3422 4176
rect 3478 4120 3483 4176
rect 0 4118 3483 4120
rect 0 4088 800 4118
rect 3417 4115 3483 4118
rect 20670 4176 23815 4178
rect 20670 4120 23754 4176
rect 23810 4120 23815 4176
rect 20670 4118 23815 4120
rect 12249 4042 12315 4045
rect 20670 4042 20730 4118
rect 23749 4115 23815 4118
rect 12249 4040 20730 4042
rect 12249 3984 12254 4040
rect 12310 3984 20730 4040
rect 12249 3982 20730 3984
rect 21173 4042 21239 4045
rect 26200 4042 27000 4072
rect 21173 4040 27000 4042
rect 21173 3984 21178 4040
rect 21234 3984 27000 4040
rect 21173 3982 27000 3984
rect 12249 3979 12315 3982
rect 21173 3979 21239 3982
rect 26200 3952 27000 3982
rect 18873 3906 18939 3909
rect 22737 3906 22803 3909
rect 18873 3904 22803 3906
rect 18873 3848 18878 3904
rect 18934 3848 22742 3904
rect 22798 3848 22803 3904
rect 18873 3846 22803 3848
rect 18873 3843 18939 3846
rect 22737 3843 22803 3846
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 19926 3770 19932 3772
rect 13494 3710 19932 3770
rect 12617 3634 12683 3637
rect 13494 3634 13554 3710
rect 19926 3708 19932 3710
rect 19996 3708 20002 3772
rect 12617 3632 13554 3634
rect 12617 3576 12622 3632
rect 12678 3576 13554 3632
rect 12617 3574 13554 3576
rect 17493 3634 17559 3637
rect 23381 3634 23447 3637
rect 17493 3632 23447 3634
rect 17493 3576 17498 3632
rect 17554 3576 23386 3632
rect 23442 3576 23447 3632
rect 17493 3574 23447 3576
rect 12617 3571 12683 3574
rect 17493 3571 17559 3574
rect 23381 3571 23447 3574
rect 19006 3436 19012 3500
rect 19076 3498 19082 3500
rect 23933 3498 23999 3501
rect 19076 3496 23999 3498
rect 19076 3440 23938 3496
rect 23994 3440 23999 3496
rect 19076 3438 23999 3440
rect 19076 3436 19082 3438
rect 23933 3435 23999 3438
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 20345 3226 20411 3229
rect 22093 3226 22159 3229
rect 20345 3224 22159 3226
rect 20345 3168 20350 3224
rect 20406 3168 22098 3224
rect 22154 3168 22159 3224
rect 20345 3166 22159 3168
rect 20345 3163 20411 3166
rect 22093 3163 22159 3166
rect 23105 3226 23171 3229
rect 26200 3226 27000 3256
rect 23105 3224 27000 3226
rect 23105 3168 23110 3224
rect 23166 3168 27000 3224
rect 23105 3166 27000 3168
rect 23105 3163 23171 3166
rect 26200 3136 27000 3166
rect 20529 3090 20595 3093
rect 23749 3090 23815 3093
rect 20529 3088 23815 3090
rect 20529 3032 20534 3088
rect 20590 3032 23754 3088
rect 23810 3032 23815 3088
rect 20529 3030 23815 3032
rect 20529 3027 20595 3030
rect 23749 3027 23815 3030
rect 14641 2954 14707 2957
rect 24945 2954 25011 2957
rect 14641 2952 25011 2954
rect 14641 2896 14646 2952
rect 14702 2896 24950 2952
rect 25006 2896 25011 2952
rect 14641 2894 25011 2896
rect 14641 2891 14707 2894
rect 24945 2891 25011 2894
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 5441 2546 5507 2549
rect 13854 2546 13860 2548
rect 5441 2544 13860 2546
rect 5441 2488 5446 2544
rect 5502 2488 13860 2544
rect 5441 2486 13860 2488
rect 5441 2483 5507 2486
rect 13854 2484 13860 2486
rect 13924 2484 13930 2548
rect 21173 2410 21239 2413
rect 26200 2410 27000 2440
rect 21173 2408 27000 2410
rect 21173 2352 21178 2408
rect 21234 2352 27000 2408
rect 21173 2350 27000 2352
rect 21173 2347 21239 2350
rect 26200 2320 27000 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 0 1866 800 1896
rect 3509 1866 3575 1869
rect 0 1864 3575 1866
rect 0 1808 3514 1864
rect 3570 1808 3575 1864
rect 0 1806 3575 1808
rect 0 1776 800 1806
rect 3509 1803 3575 1806
rect 22185 1594 22251 1597
rect 26200 1594 27000 1624
rect 22185 1592 27000 1594
rect 22185 1536 22190 1592
rect 22246 1536 27000 1592
rect 22185 1534 27000 1536
rect 22185 1531 22251 1534
rect 26200 1504 27000 1534
rect 25313 778 25379 781
rect 26200 778 27000 808
rect 25313 776 27000 778
rect 25313 720 25318 776
rect 25374 720 27000 776
rect 25313 718 27000 720
rect 25313 715 25379 718
rect 26200 688 27000 718
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 21404 44236 21468 44300
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 17172 25060 17236 25124
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 19932 24984 19996 24988
rect 19932 24928 19946 24984
rect 19946 24928 19996 24984
rect 19932 24924 19996 24928
rect 16436 24788 16500 24852
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 19012 23428 19076 23492
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 17356 23156 17420 23220
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 14044 20708 14108 20772
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 17540 18668 17604 18732
rect 21404 18668 21468 18732
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 21220 17988 21284 18052
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 17172 17308 17236 17372
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 17356 16220 17420 16284
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 16988 15268 17052 15332
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 13860 14240 13924 14244
rect 13860 14184 13910 14240
rect 13910 14184 13924 14240
rect 13860 14180 13924 14184
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 17540 13560 17604 13564
rect 17540 13504 17554 13560
rect 17554 13504 17604 13560
rect 17540 13500 17604 13504
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 16988 11052 17052 11116
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 14044 10704 14108 10708
rect 14044 10648 14058 10704
rect 14058 10648 14108 10704
rect 14044 10644 14108 10648
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 21220 9420 21284 9484
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 19748 6896 19812 6900
rect 19748 6840 19762 6896
rect 19762 6840 19812 6896
rect 19748 6836 19812 6840
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 14044 6292 14108 6356
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 16436 5748 16500 5812
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 19748 4584 19812 4588
rect 19748 4528 19762 4584
rect 19762 4528 19812 4584
rect 19748 4524 19812 4528
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 19932 3708 19996 3772
rect 19012 3436 19076 3500
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 13860 2484 13924 2548
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 53888 13264 54448
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 17944 53344 18264 54368
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 21403 44300 21469 44301
rect 21403 44236 21404 44300
rect 21468 44236 21469 44300
rect 21403 44235 21469 44236
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17944 38112 18264 39136
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17944 27232 18264 28256
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17171 25124 17237 25125
rect 17171 25060 17172 25124
rect 17236 25060 17237 25124
rect 17171 25059 17237 25060
rect 16435 24852 16501 24853
rect 16435 24788 16436 24852
rect 16500 24788 16501 24852
rect 16435 24787 16501 24788
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 14043 20772 14109 20773
rect 14043 20708 14044 20772
rect 14108 20708 14109 20772
rect 14043 20707 14109 20708
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 13859 14244 13925 14245
rect 13859 14180 13860 14244
rect 13924 14180 13925 14244
rect 13859 14179 13925 14180
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 13862 2549 13922 14179
rect 14046 10709 14106 20707
rect 14043 10708 14109 10709
rect 14043 10644 14044 10708
rect 14108 10644 14109 10708
rect 14043 10643 14109 10644
rect 14046 6357 14106 10643
rect 14043 6356 14109 6357
rect 14043 6292 14044 6356
rect 14108 6292 14109 6356
rect 14043 6291 14109 6292
rect 16438 5813 16498 24787
rect 17174 17373 17234 25059
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 19931 24988 19997 24989
rect 19931 24924 19932 24988
rect 19996 24924 19997 24988
rect 19931 24923 19997 24924
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17355 23220 17421 23221
rect 17355 23156 17356 23220
rect 17420 23156 17421 23220
rect 17355 23155 17421 23156
rect 17171 17372 17237 17373
rect 17171 17308 17172 17372
rect 17236 17308 17237 17372
rect 17171 17307 17237 17308
rect 17358 16285 17418 23155
rect 17944 22880 18264 23904
rect 19011 23492 19077 23493
rect 19011 23428 19012 23492
rect 19076 23428 19077 23492
rect 19011 23427 19077 23428
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17539 18732 17605 18733
rect 17539 18668 17540 18732
rect 17604 18668 17605 18732
rect 17539 18667 17605 18668
rect 17355 16284 17421 16285
rect 17355 16220 17356 16284
rect 17420 16220 17421 16284
rect 17355 16219 17421 16220
rect 16987 15332 17053 15333
rect 16987 15268 16988 15332
rect 17052 15268 17053 15332
rect 16987 15267 17053 15268
rect 16990 11117 17050 15267
rect 17542 13565 17602 18667
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17539 13564 17605 13565
rect 17539 13500 17540 13564
rect 17604 13500 17605 13564
rect 17539 13499 17605 13500
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 16987 11116 17053 11117
rect 16987 11052 16988 11116
rect 17052 11052 17053 11116
rect 16987 11051 17053 11052
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 16435 5812 16501 5813
rect 16435 5748 16436 5812
rect 16500 5748 16501 5812
rect 16435 5747 16501 5748
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 19014 3501 19074 23427
rect 19747 6900 19813 6901
rect 19747 6836 19748 6900
rect 19812 6836 19813 6900
rect 19747 6835 19813 6836
rect 19750 4589 19810 6835
rect 19747 4588 19813 4589
rect 19747 4524 19748 4588
rect 19812 4524 19813 4588
rect 19747 4523 19813 4524
rect 19934 3773 19994 24923
rect 21406 18733 21466 44235
rect 22944 44096 23264 45120
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 21403 18732 21469 18733
rect 21403 18668 21404 18732
rect 21468 18668 21469 18732
rect 21403 18667 21469 18668
rect 21219 18052 21285 18053
rect 21219 17988 21220 18052
rect 21284 17988 21285 18052
rect 21219 17987 21285 17988
rect 21222 9485 21282 17987
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 21219 9484 21285 9485
rect 21219 9420 21220 9484
rect 21284 9420 21285 9484
rect 21219 9419 21285 9420
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 19931 3772 19997 3773
rect 19931 3708 19932 3772
rect 19996 3708 19997 3772
rect 19931 3707 19997 3708
rect 19011 3500 19077 3501
rect 19011 3436 19012 3500
rect 19076 3436 19077 3500
rect 19011 3435 19077 3436
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 13859 2548 13925 2549
rect 13859 2484 13860 2548
rect 13924 2484 13925 2548
rect 13859 2483 13925 2484
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
use sky130_fd_sc_hd__clkbuf_2  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _105_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15456 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _106_
timestamp 1676037725
transform 1 0 11040 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _107_
timestamp 1676037725
transform 1 0 18032 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _108_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _109_
timestamp 1676037725
transform 1 0 21344 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _110_
timestamp 1676037725
transform 1 0 10304 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _111_
timestamp 1676037725
transform 1 0 24472 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _112_
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _113_
timestamp 1676037725
transform 1 0 11868 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _114_
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform 1 0 24564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1676037725
transform 1 0 24564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1676037725
transform 1 0 25024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1676037725
transform 1 0 24840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1676037725
transform 1 0 25024 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1676037725
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1676037725
transform 1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1676037725
transform 1 0 21988 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1676037725
transform 1 0 21988 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1676037725
transform 1 0 22724 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1676037725
transform 1 0 21988 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1676037725
transform 1 0 20792 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1676037725
transform 1 0 21620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1676037725
transform 1 0 23736 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1676037725
transform 1 0 22172 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1676037725
transform 1 0 20792 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1676037725
transform 1 0 21528 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1676037725
transform 1 0 19412 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1676037725
transform 1 0 19688 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform 1 0 16836 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1676037725
transform 1 0 17112 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1676037725
transform 1 0 14260 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 13800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 16744 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 17480 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 17756 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 18492 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 19412 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 19228 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform 1 0 19412 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 18584 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 16008 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform 1 0 14536 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1676037725
transform 1 0 20792 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1676037725
transform 1 0 21896 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1676037725
transform 1 0 20516 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1676037725
transform 1 0 21804 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 20976 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 23092 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1676037725
transform 1 0 23828 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 22724 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1676037725
transform 1 0 21988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1676037725
transform 1 0 24564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1676037725
transform 1 0 23460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform 1 0 23552 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1676037725
transform 1 0 5152 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1676037725
transform 1 0 6532 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1676037725
transform 1 0 7544 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1676037725
transform 1 0 9200 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1676037725
transform 1 0 8280 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1676037725
transform 1 0 9384 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1676037725
transform 1 0 10396 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1676037725
transform 1 0 11408 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15916 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 20516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 11684 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1676037725
transform 1 0 20240 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A
timestamp 1676037725
transform 1 0 18400 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A
timestamp 1676037725
transform 1 0 17480 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1676037725
transform 1 0 12788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1676037725
transform 1 0 20608 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1676037725
transform 1 0 21160 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1676037725
transform 1 0 21344 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A
timestamp 1676037725
transform 1 0 16836 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A
timestamp 1676037725
transform 1 0 14168 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1676037725
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1676037725
transform 1 0 21988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1676037725
transform 1 0 25116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A
timestamp 1676037725
transform 1 0 21896 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1676037725
transform 1 0 25392 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1676037725
transform 1 0 25300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A
timestamp 1676037725
transform 1 0 25300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A
timestamp 1676037725
transform 1 0 25116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A
timestamp 1676037725
transform 1 0 24104 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 7820 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 8556 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10120 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 9292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 8464 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 9568 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12052 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__D
timestamp 1676037725
transform 1 0 11132 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 10948 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 10028 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11868 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__D
timestamp 1676037725
transform 1 0 10120 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 10028 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3__RESET_B
timestamp 1676037725
transform 1 0 10948 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15272 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 12604 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 15272 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16100 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 14352 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2__S
timestamp 1676037725
transform 1 0 14168 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 16008 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 14628 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3__S
timestamp 1676037725
transform 1 0 15456 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 13432 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 12236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4__S
timestamp 1676037725
transform 1 0 12420 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 18124 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16928 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 16284 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2__A1
timestamp 1676037725
transform 1 0 15456 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 16192 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 15272 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 9476 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16744 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15732 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 17112 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 15180 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 14168 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 13156 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0__S
timestamp 1676037725
transform 1 0 11868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1__S
timestamp 1676037725
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 9844 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2__S
timestamp 1676037725
transform 1 0 11224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 15732 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__S
timestamp 1676037725
transform 1 0 14352 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15272 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 15640 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1676037725
transform 1 0 15456 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A0
timestamp 1676037725
transform 1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3__A1
timestamp 1676037725
transform 1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A0
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4__A1
timestamp 1676037725
transform 1 0 13708 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0__S
timestamp 1676037725
transform 1 0 11776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1__S
timestamp 1676037725
transform 1 0 12604 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1676037725
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2__S
timestamp 1676037725
transform 1 0 11040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1676037725
transform 1 0 17296 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__S
timestamp 1676037725
transform 1 0 15272 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 11684 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 11040 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 11684 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 10120 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 11316 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11132 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1676037725
transform 1 0 8280 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1676037725
transform 1 0 8832 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8648 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1676037725
transform 1 0 18860 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1676037725
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1676037725
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1676037725
transform 1 0 20792 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1676037725
transform 1 0 16744 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1676037725
transform 1 0 15732 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1676037725
transform 1 0 15548 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1676037725
transform 1 0 15824 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1676037725
transform 1 0 16928 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1676037725
transform 1 0 19320 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1676037725
transform 1 0 19504 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1676037725
transform 1 0 21528 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold3_A
timestamp 1676037725
transform 1 0 25300 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold4_A
timestamp 1676037725
transform 1 0 2024 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold6_A
timestamp 1676037725
transform 1 0 23920 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1676037725
transform 1 0 24748 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1676037725
transform 1 0 25392 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1676037725
transform 1 0 24748 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1676037725
transform 1 0 25392 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1676037725
transform 1 0 24656 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1676037725
transform 1 0 25392 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1676037725
transform 1 0 24748 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1676037725
transform 1 0 25392 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1676037725
transform 1 0 24748 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1676037725
transform 1 0 25392 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1676037725
transform 1 0 25208 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1676037725
transform 1 0 24656 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1676037725
transform 1 0 25392 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1676037725
transform 1 0 24656 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1676037725
transform 1 0 25392 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1676037725
transform 1 0 24748 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1676037725
transform 1 0 25392 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1676037725
transform 1 0 24748 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1676037725
transform 1 0 25392 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1676037725
transform 1 0 24656 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1676037725
transform 1 0 25392 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1676037725
transform 1 0 24564 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1676037725
transform 1 0 22816 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1676037725
transform 1 0 25392 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1676037725
transform 1 0 25392 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1676037725
transform 1 0 24748 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1676037725
transform 1 0 24748 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1676037725
transform 1 0 24748 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1676037725
transform 1 0 3128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1676037725
transform 1 0 4784 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1676037725
transform 1 0 4140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1676037725
transform 1 0 6900 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1676037725
transform 1 0 7820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1676037725
transform 1 0 7636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1676037725
transform 1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1676037725
transform 1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1676037725
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1676037725
transform 1 0 8924 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1676037725
transform 1 0 9292 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1676037725
transform 1 0 9108 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1676037725
transform 1 0 8924 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1676037725
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1676037725
transform 1 0 9108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1676037725
transform 1 0 9752 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1676037725
transform 1 0 9292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1676037725
transform 1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1676037725
transform 1 0 9936 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1676037725
transform 1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1676037725
transform 1 0 3312 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1676037725
transform 1 0 3772 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1676037725
transform 1 0 4508 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1676037725
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1676037725
transform 1 0 13800 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1676037725
transform 1 0 15364 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1676037725
transform 1 0 17296 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1676037725
transform 1 0 18124 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1676037725
transform 1 0 18952 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1676037725
transform 1 0 9844 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1676037725
transform 1 0 24472 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1676037725
transform 1 0 24472 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1676037725
transform 1 0 24472 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1676037725
transform 1 0 24748 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1676037725
transform 1 0 24104 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1676037725
transform 1 0 24656 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1676037725
transform 1 0 22632 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1676037725
transform 1 0 21252 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1676037725
transform 1 0 22540 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1676037725
transform 1 0 23736 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1676037725
transform 1 0 23920 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output113_A
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output122_A
timestamp 1676037725
transform 1 0 25116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output124_A
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output135_A
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 20608 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25392 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25300 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21436 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 23920 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25208 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25392 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24748 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24748 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25208 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21436 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19964 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18952 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18768 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18768 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19412 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22724 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24472 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25300 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24564 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24104 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24288 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23644 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21068 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 23828 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25392 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22356 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 15456 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15640 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__D
timestamp 1676037725
transform 1 0 11316 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 11132 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13708 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12512 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13156 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13616 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 13432 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15824 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15272 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15456 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12880 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 11408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10120 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1676037725
transform 1 0 8372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10948 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12696 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14536 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 15088 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14536 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 12052 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 10948 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 12788 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 13432 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16744 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16928 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17204 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18124 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18676 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 14720 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 16100 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 17848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 20424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22264 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 22632 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22632 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21252 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 22264 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24012 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25024 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25024 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 25116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 25300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 24104 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 24196 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 21988 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19872 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1676037725
transform 1 0 19320 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1676037725
transform 1 0 18860 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1676037725
transform 1 0 19044 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20332 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 19136 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 25392 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 18860 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22264 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 25024 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 25392 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24012 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19964 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19688 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_31.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21436 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22632 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_35.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24472 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_45.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 22356 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_47.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21804 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_49.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20332 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_51.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 24104 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_bottom_track_51.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 25208 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16928 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16744 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 16560 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 16744 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l2_in_0__S
timestamp 1676037725
transform 1 0 13340 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 7268 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_0.mux_l2_in_1__S
timestamp 1676037725
transform 1 0 8464 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16008 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16192 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16192 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_2.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 9016 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16192 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 16836 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_4.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 10304 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18032 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17848 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 18676 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 18492 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_6.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 11132 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 16192 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 16376 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 17204 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 17020 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_8.mux_l2_in_1__A1
timestamp 1676037725
transform 1 0 8648 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 15088 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15272 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_1__A0
timestamp 1676037725
transform 1 0 16836 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_10.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16652 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_12.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 14352 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_12.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18032 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18216 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_14.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 12052 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19044 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19228 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_16.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 12420 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_18.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 14720 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_18.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_20.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_20.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_22.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_24.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 12696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_26.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_26.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 15272 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18492 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18676 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_28.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 13340 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19044 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_30.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 16192 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18676 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18860 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_32.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 15180 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_34.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 17848 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_34.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18032 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_36.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14352 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_38.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_40.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 17848 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_42.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 17572 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_42.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20424 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21252 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_44.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 17756 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21160 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21344 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_46.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 19964 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21436 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_48.mux_l1_in_1__A1
timestamp 1676037725
transform 1 0 19964 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20976 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 22448 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0__A
timestamp 1676037725
transform 1 0 10580 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_52.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 20148 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_52.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 22448 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_54.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_56.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__A0
timestamp 1676037725
transform 1 0 18768 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__A1
timestamp 1676037725
transform 1 0 18584 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_0__S
timestamp 1676037725
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_0__8_.mux_right_track_58.mux_l1_in_1__S
timestamp 1676037725
transform 1 0 11868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5060 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8188 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6532 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6532 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7636 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9292 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 7268 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6440 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7728 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9936 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 7728 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6900 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 7728 0 -1 20672
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9752 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 8004 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 9108 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14260 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13892 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 14536 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 14996 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11592 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11408 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9016 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__194 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 10396 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10120 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 9108 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 8740 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15824 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 17112 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 15088 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 14260 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12604 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9844 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__195
timestamp 1676037725
transform 1 0 11684 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 12788 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10212 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 9200 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8924 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15916 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 13800 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 11868 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 13340 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12420 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 10212 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__196
timestamp 1676037725
transform 1 0 15640 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 14720 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 12696 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 13064 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 12604 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 13800 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12144 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11592 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__197
timestamp 1676037725
transform 1 0 16008 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 14812 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 9476 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8648 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15640 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 13248 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10580 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10212 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 14812 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 12512 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 10304 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 9568 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 13892 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 11592 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 9384 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 8924 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9108 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 12696 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 10304 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 7544 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 7912 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6624 0 -1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 15916 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10212 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 12604 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 10212 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 12420 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 17296 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 19412 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 17204 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 19228 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 14076 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 14352 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 14628 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 15364 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 20332 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 22172 0 -1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 19872 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 22080 0 -1 32640
box -38 -48 1050 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2484 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35
timestamp 1676037725
transform 1 0 4324 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1676037725
transform 1 0 6900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68
timestamp 1676037725
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1676037725
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1676037725
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_118
timestamp 1676037725
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_143
timestamp 1676037725
transform 1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_161
timestamp 1676037725
transform 1 0 15916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_165
timestamp 1676037725
transform 1 0 16284 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_187
timestamp 1676037725
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_215
timestamp 1676037725
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_243
timestamp 1676037725
transform 1 0 23460 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_263 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1676037725
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_35
timestamp 1676037725
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_42
timestamp 1676037725
transform 1 0 4968 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1676037725
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1676037725
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_83
timestamp 1676037725
transform 1 0 8740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_91
timestamp 1676037725
transform 1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1676037725
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_103
timestamp 1676037725
transform 1 0 10580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1676037725
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1676037725
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1676037725
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1676037725
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_207
timestamp 1676037725
transform 1 0 20148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1676037725
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_231
timestamp 1676037725
transform 1 0 22356 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_239
timestamp 1676037725
transform 1 0 23092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_247
timestamp 1676037725
transform 1 0 23828 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_254
timestamp 1676037725
transform 1 0 24472 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_258
timestamp 1676037725
transform 1 0 24840 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_262
timestamp 1676037725
transform 1 0 25208 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_22
timestamp 1676037725
transform 1 0 3128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_31
timestamp 1676037725
transform 1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1676037725
transform 1 0 4508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_51
timestamp 1676037725
transform 1 0 5796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_55
timestamp 1676037725
transform 1 0 6164 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_60
timestamp 1676037725
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_64
timestamp 1676037725
transform 1 0 6992 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_68
timestamp 1676037725
transform 1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_75
timestamp 1676037725
transform 1 0 8004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1676037725
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_91
timestamp 1676037725
transform 1 0 9476 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_96
timestamp 1676037725
transform 1 0 9936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_100
timestamp 1676037725
transform 1 0 10304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_104
timestamp 1676037725
transform 1 0 10672 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_118
timestamp 1676037725
transform 1 0 11960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1676037725
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1676037725
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_179
timestamp 1676037725
transform 1 0 17572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_183
timestamp 1676037725
transform 1 0 17940 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1676037725
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1676037725
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_235
timestamp 1676037725
transform 1 0 22724 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_239
timestamp 1676037725
transform 1 0 23092 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_243
timestamp 1676037725
transform 1 0 23460 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_250
timestamp 1676037725
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_263
timestamp 1676037725
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1676037725
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_20
timestamp 1676037725
transform 1 0 2944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_24
timestamp 1676037725
transform 1 0 3312 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_28
timestamp 1676037725
transform 1 0 3680 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_31
timestamp 1676037725
transform 1 0 3956 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_36
timestamp 1676037725
transform 1 0 4416 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_41
timestamp 1676037725
transform 1 0 4876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_53
timestamp 1676037725
transform 1 0 5980 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_57 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_65
timestamp 1676037725
transform 1 0 7084 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_77
timestamp 1676037725
transform 1 0 8188 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_87
timestamp 1676037725
transform 1 0 9108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 1676037725
transform 1 0 9568 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_98
timestamp 1676037725
transform 1 0 10120 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1676037725
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_117
timestamp 1676037725
transform 1 0 11868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_135
timestamp 1676037725
transform 1 0 13524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_159
timestamp 1676037725
transform 1 0 15732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1676037725
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1676037725
transform 1 0 18308 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_207
timestamp 1676037725
transform 1 0 20148 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_220
timestamp 1676037725
transform 1 0 21344 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_229
timestamp 1676037725
transform 1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_252
timestamp 1676037725
transform 1 0 24288 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_259
timestamp 1676037725
transform 1 0 24932 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_265
timestamp 1676037725
transform 1 0 25484 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_8
timestamp 1676037725
transform 1 0 1840 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_12
timestamp 1676037725
transform 1 0 2208 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1676037725
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_39
timestamp 1676037725
transform 1 0 4692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1676037725
transform 1 0 7176 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_70
timestamp 1676037725
transform 1 0 7544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1676037725
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_99
timestamp 1676037725
transform 1 0 10212 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_104
timestamp 1676037725
transform 1 0 10672 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_118
timestamp 1676037725
transform 1 0 11960 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1676037725
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_146
timestamp 1676037725
transform 1 0 14536 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_150
timestamp 1676037725
transform 1 0 14904 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_172
timestamp 1676037725
transform 1 0 16928 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_176
timestamp 1676037725
transform 1 0 17296 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1676037725
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_220
timestamp 1676037725
transform 1 0 21344 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_240
timestamp 1676037725
transform 1 0 23184 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_248
timestamp 1676037725
transform 1 0 23920 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_259
timestamp 1676037725
transform 1 0 24932 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1676037725
transform 1 0 10396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1676037725
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_127
timestamp 1676037725
transform 1 0 12788 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_151
timestamp 1676037725
transform 1 0 14996 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_155
timestamp 1676037725
transform 1 0 15364 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1676037725
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_188
timestamp 1676037725
transform 1 0 18400 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_212
timestamp 1676037725
transform 1 0 20608 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_220
timestamp 1676037725
transform 1 0 21344 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1676037725
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_263
timestamp 1676037725
transform 1 0 25300 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_117
timestamp 1676037725
transform 1 0 11868 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_131
timestamp 1676037725
transform 1 0 13156 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1676037725
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_143
timestamp 1676037725
transform 1 0 14260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_146
timestamp 1676037725
transform 1 0 14536 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_157
timestamp 1676037725
transform 1 0 15548 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_181
timestamp 1676037725
transform 1 0 17756 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1676037725
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1676037725
transform 1 0 20884 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_235
timestamp 1676037725
transform 1 0 22724 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_243
timestamp 1676037725
transform 1 0 23460 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1676037725
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_259
timestamp 1676037725
transform 1 0 24932 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1676037725
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_124
timestamp 1676037725
transform 1 0 12512 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_130
timestamp 1676037725
transform 1 0 13064 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_142
timestamp 1676037725
transform 1 0 14168 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_146
timestamp 1676037725
transform 1 0 14536 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1676037725
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_180
timestamp 1676037725
transform 1 0 17664 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_184
timestamp 1676037725
transform 1 0 18032 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_202
timestamp 1676037725
transform 1 0 19688 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1676037725
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_247
timestamp 1676037725
transform 1 0 23828 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_253
timestamp 1676037725
transform 1 0 24380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_258
timestamp 1676037725
transform 1 0 24840 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_125
timestamp 1676037725
transform 1 0 12604 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_129
timestamp 1676037725
transform 1 0 12972 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1676037725
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_144
timestamp 1676037725
transform 1 0 14352 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_150
timestamp 1676037725
transform 1 0 14904 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_170
timestamp 1676037725
transform 1 0 16744 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1676037725
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_208
timestamp 1676037725
transform 1 0 20240 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1676037725
transform 1 0 20608 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_230
timestamp 1676037725
transform 1 0 22264 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1676037725
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_264
timestamp 1676037725
transform 1 0 25392 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_85
timestamp 1676037725
transform 1 0 8924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp 1676037725
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1676037725
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_119
timestamp 1676037725
transform 1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_130
timestamp 1676037725
transform 1 0 13064 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_136
timestamp 1676037725
transform 1 0 13616 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_157
timestamp 1676037725
transform 1 0 15548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1676037725
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_173
timestamp 1676037725
transform 1 0 17020 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_185
timestamp 1676037725
transform 1 0 18124 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_209
timestamp 1676037725
transform 1 0 20332 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1676037725
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_244
timestamp 1676037725
transform 1 0 23552 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1676037725
transform 1 0 25392 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_105
timestamp 1676037725
transform 1 0 10764 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_117
timestamp 1676037725
transform 1 0 11868 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_125
timestamp 1676037725
transform 1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1676037725
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_152
timestamp 1676037725
transform 1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_156
timestamp 1676037725
transform 1 0 15456 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_169
timestamp 1676037725
transform 1 0 16652 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1676037725
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_202
timestamp 1676037725
transform 1 0 19688 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_206
timestamp 1676037725
transform 1 0 20056 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_224
timestamp 1676037725
transform 1 0 21712 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_248
timestamp 1676037725
transform 1 0 23920 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_259
timestamp 1676037725
transform 1 0 24932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_118
timestamp 1676037725
transform 1 0 11960 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_126
timestamp 1676037725
transform 1 0 12696 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_129
timestamp 1676037725
transform 1 0 12972 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_134
timestamp 1676037725
transform 1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_142
timestamp 1676037725
transform 1 0 14168 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_146
timestamp 1676037725
transform 1 0 14536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1676037725
transform 1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1676037725
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_180
timestamp 1676037725
transform 1 0 17664 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_184
timestamp 1676037725
transform 1 0 18032 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_202
timestamp 1676037725
transform 1 0 19688 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1676037725
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_244
timestamp 1676037725
transform 1 0 23552 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_264
timestamp 1676037725
transform 1 0 25392 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_107
timestamp 1676037725
transform 1 0 10948 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_111
timestamp 1676037725
transform 1 0 11316 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_123
timestamp 1676037725
transform 1 0 12420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_127
timestamp 1676037725
transform 1 0 12788 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1676037725
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_152
timestamp 1676037725
transform 1 0 15088 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_158
timestamp 1676037725
transform 1 0 15640 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_170
timestamp 1676037725
transform 1 0 16744 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_183
timestamp 1676037725
transform 1 0 17940 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_187
timestamp 1676037725
transform 1 0 18308 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1676037725
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_228
timestamp 1676037725
transform 1 0 22080 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_232
timestamp 1676037725
transform 1 0 22448 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1676037725
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_258
timestamp 1676037725
transform 1 0 24840 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_109
timestamp 1676037725
transform 1 0 11132 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp 1676037725
transform 1 0 13524 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_148
timestamp 1676037725
transform 1 0 14720 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_174
timestamp 1676037725
transform 1 0 17112 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_196
timestamp 1676037725
transform 1 0 19136 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_200
timestamp 1676037725
transform 1 0 19504 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1676037725
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_230
timestamp 1676037725
transform 1 0 22264 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_254
timestamp 1676037725
transform 1 0 24472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_261
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_265
timestamp 1676037725
transform 1 0 25484 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_110
timestamp 1676037725
transform 1 0 11224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_123
timestamp 1676037725
transform 1 0 12420 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_136
timestamp 1676037725
transform 1 0 13616 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_144
timestamp 1676037725
transform 1 0 14352 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_155
timestamp 1676037725
transform 1 0 15364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_166
timestamp 1676037725
transform 1 0 16376 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_174
timestamp 1676037725
transform 1 0 17112 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_182
timestamp 1676037725
transform 1 0 17848 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_192
timestamp 1676037725
transform 1 0 18768 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_203
timestamp 1676037725
transform 1 0 19780 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_231
timestamp 1676037725
transform 1 0 22356 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_235
timestamp 1676037725
transform 1 0 22724 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_258
timestamp 1676037725
transform 1 0 24840 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_75
timestamp 1676037725
transform 1 0 8004 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_98
timestamp 1676037725
transform 1 0 10120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_102
timestamp 1676037725
transform 1 0 10488 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_106
timestamp 1676037725
transform 1 0 10856 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_109
timestamp 1676037725
transform 1 0 11132 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1676037725
transform 1 0 11960 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_131
timestamp 1676037725
transform 1 0 13156 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 1676037725
transform 1 0 13616 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_147
timestamp 1676037725
transform 1 0 14628 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_155
timestamp 1676037725
transform 1 0 15364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1676037725
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1676037725
transform 1 0 17112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_182
timestamp 1676037725
transform 1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_189
timestamp 1676037725
transform 1 0 18492 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1676037725
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_209
timestamp 1676037725
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1676037725
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_230
timestamp 1676037725
transform 1 0 22264 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_236
timestamp 1676037725
transform 1 0 22816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_259
timestamp 1676037725
transform 1 0 24932 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_263
timestamp 1676037725
transform 1 0 25300 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_107
timestamp 1676037725
transform 1 0 10948 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_111
timestamp 1676037725
transform 1 0 11316 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_134
timestamp 1676037725
transform 1 0 13432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_146
timestamp 1676037725
transform 1 0 14536 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_176
timestamp 1676037725
transform 1 0 17296 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_183
timestamp 1676037725
transform 1 0 17940 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_199
timestamp 1676037725
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1676037725
transform 1 0 20424 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_218
timestamp 1676037725
transform 1 0 21160 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_225
timestamp 1676037725
transform 1 0 21804 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_229
timestamp 1676037725
transform 1 0 22172 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_233
timestamp 1676037725
transform 1 0 22540 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_250
timestamp 1676037725
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_259
timestamp 1676037725
transform 1 0 24932 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_263
timestamp 1676037725
transform 1 0 25300 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_65
timestamp 1676037725
transform 1 0 7084 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_87
timestamp 1676037725
transform 1 0 9108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_104
timestamp 1676037725
transform 1 0 10672 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_115
timestamp 1676037725
transform 1 0 11684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_126
timestamp 1676037725
transform 1 0 12696 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_139
timestamp 1676037725
transform 1 0 13892 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_152
timestamp 1676037725
transform 1 0 15088 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_158
timestamp 1676037725
transform 1 0 15640 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1676037725
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_180
timestamp 1676037725
transform 1 0 17664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_193
timestamp 1676037725
transform 1 0 18860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_201
timestamp 1676037725
transform 1 0 19596 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_209
timestamp 1676037725
transform 1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_216
timestamp 1676037725
transform 1 0 20976 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_244
timestamp 1676037725
transform 1 0 23552 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_264
timestamp 1676037725
transform 1 0 25392 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_71
timestamp 1676037725
transform 1 0 7636 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1676037725
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_87
timestamp 1676037725
transform 1 0 9108 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_108
timestamp 1676037725
transform 1 0 11040 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_134
timestamp 1676037725
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_152
timestamp 1676037725
transform 1 0 15088 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_160
timestamp 1676037725
transform 1 0 15824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_164
timestamp 1676037725
transform 1 0 16192 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1676037725
transform 1 0 16468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_172
timestamp 1676037725
transform 1 0 16928 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_187
timestamp 1676037725
transform 1 0 18308 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1676037725
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_203
timestamp 1676037725
transform 1 0 19780 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_207
timestamp 1676037725
transform 1 0 20148 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_230
timestamp 1676037725
transform 1 0 22264 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1676037725
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_258
timestamp 1676037725
transform 1 0 24840 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_82
timestamp 1676037725
transform 1 0 8648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_95
timestamp 1676037725
transform 1 0 9844 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1676037725
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1676037725
transform 1 0 12420 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_134
timestamp 1676037725
transform 1 0 13432 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_147
timestamp 1676037725
transform 1 0 14628 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_160
timestamp 1676037725
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1676037725
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_180
timestamp 1676037725
transform 1 0 17664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_187
timestamp 1676037725
transform 1 0 18308 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_191
timestamp 1676037725
transform 1 0 18676 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_201
timestamp 1676037725
transform 1 0 19596 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_208
timestamp 1676037725
transform 1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_212
timestamp 1676037725
transform 1 0 20608 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_230
timestamp 1676037725
transform 1 0 22264 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_236
timestamp 1676037725
transform 1 0 22816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_259
timestamp 1676037725
transform 1 0 24932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_263
timestamp 1676037725
transform 1 0 25300 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_79
timestamp 1676037725
transform 1 0 8372 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_136
timestamp 1676037725
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1676037725
transform 1 0 14996 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_162
timestamp 1676037725
transform 1 0 16008 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_166
timestamp 1676037725
transform 1 0 16376 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_174
timestamp 1676037725
transform 1 0 17112 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_179
timestamp 1676037725
transform 1 0 17572 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_185
timestamp 1676037725
transform 1 0 18124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1676037725
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1676037725
transform 1 0 20424 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_218
timestamp 1676037725
transform 1 0 21160 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_230
timestamp 1676037725
transform 1 0 22264 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1676037725
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_258
timestamp 1676037725
transform 1 0 24840 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_262
timestamp 1676037725
transform 1 0 25208 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1676037725
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1676037725
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1676037725
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1676037725
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1676037725
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_95
timestamp 1676037725
transform 1 0 9844 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1676037725
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_118
timestamp 1676037725
transform 1 0 11960 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1676037725
transform 1 0 12420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_134
timestamp 1676037725
transform 1 0 13432 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_158
timestamp 1676037725
transform 1 0 15640 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_162
timestamp 1676037725
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_191
timestamp 1676037725
transform 1 0 18676 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_197
timestamp 1676037725
transform 1 0 19228 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_203
timestamp 1676037725
transform 1 0 19780 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_210
timestamp 1676037725
transform 1 0 20424 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_214
timestamp 1676037725
transform 1 0 20792 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_218
timestamp 1676037725
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_230
timestamp 1676037725
transform 1 0 22264 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1676037725
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_263
timestamp 1676037725
transform 1 0 25300 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_57
timestamp 1676037725
transform 1 0 6348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_78
timestamp 1676037725
transform 1 0 8280 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1676037725
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1676037725
transform 1 0 9476 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_94
timestamp 1676037725
transform 1 0 9752 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_119
timestamp 1676037725
transform 1 0 12052 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1676037725
transform 1 0 13248 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_136
timestamp 1676037725
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_152
timestamp 1676037725
transform 1 0 15088 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_156
timestamp 1676037725
transform 1 0 15456 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_164
timestamp 1676037725
transform 1 0 16192 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_176
timestamp 1676037725
transform 1 0 17296 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_183
timestamp 1676037725
transform 1 0 17940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_205
timestamp 1676037725
transform 1 0 19964 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_211
timestamp 1676037725
transform 1 0 20516 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_219
timestamp 1676037725
transform 1 0 21252 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_230
timestamp 1676037725
transform 1 0 22264 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1676037725
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_257
timestamp 1676037725
transform 1 0 24748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_261
timestamp 1676037725
transform 1 0 25116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_94
timestamp 1676037725
transform 1 0 9752 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_107
timestamp 1676037725
transform 1 0 10948 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_121
timestamp 1676037725
transform 1 0 12236 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_135
timestamp 1676037725
transform 1 0 13524 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_146
timestamp 1676037725
transform 1 0 14536 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_152
timestamp 1676037725
transform 1 0 15088 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1676037725
transform 1 0 15364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1676037725
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_177
timestamp 1676037725
transform 1 0 17388 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_180
timestamp 1676037725
transform 1 0 17664 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_188
timestamp 1676037725
transform 1 0 18400 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_194
timestamp 1676037725
transform 1 0 18952 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_200
timestamp 1676037725
transform 1 0 19504 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_210
timestamp 1676037725
transform 1 0 20424 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_217
timestamp 1676037725
transform 1 0 21068 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_221
timestamp 1676037725
transform 1 0 21436 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_244
timestamp 1676037725
transform 1 0 23552 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_264
timestamp 1676037725
transform 1 0 25392 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_96
timestamp 1676037725
transform 1 0 9936 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_100
timestamp 1676037725
transform 1 0 10304 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_112
timestamp 1676037725
transform 1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_123
timestamp 1676037725
transform 1 0 12420 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_127
timestamp 1676037725
transform 1 0 12788 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_146
timestamp 1676037725
transform 1 0 14536 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_150
timestamp 1676037725
transform 1 0 14904 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_154
timestamp 1676037725
transform 1 0 15272 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_157
timestamp 1676037725
transform 1 0 15548 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_162
timestamp 1676037725
transform 1 0 16008 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_186
timestamp 1676037725
transform 1 0 18216 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_190
timestamp 1676037725
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1676037725
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_226
timestamp 1676037725
transform 1 0 21896 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1676037725
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_258
timestamp 1676037725
transform 1 0 24840 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_262
timestamp 1676037725
transform 1 0 25208 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_79
timestamp 1676037725
transform 1 0 8372 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_83
timestamp 1676037725
transform 1 0 8740 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_95
timestamp 1676037725
transform 1 0 9844 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_107
timestamp 1676037725
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1676037725
transform 1 0 11960 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_129
timestamp 1676037725
transform 1 0 12972 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_142
timestamp 1676037725
transform 1 0 14168 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_155
timestamp 1676037725
transform 1 0 15364 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_162
timestamp 1676037725
transform 1 0 16008 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1676037725
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1676037725
transform 1 0 16928 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1676037725
transform 1 0 17480 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_185
timestamp 1676037725
transform 1 0 18124 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_192
timestamp 1676037725
transform 1 0 18768 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_196
timestamp 1676037725
transform 1 0 19136 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1676037725
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_212
timestamp 1676037725
transform 1 0 20608 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1676037725
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_247
timestamp 1676037725
transform 1 0 23828 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_251
timestamp 1676037725
transform 1 0 24196 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_264
timestamp 1676037725
transform 1 0 25392 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1676037725
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1676037725
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_108
timestamp 1676037725
transform 1 0 11040 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_112
timestamp 1676037725
transform 1 0 11408 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_136
timestamp 1676037725
transform 1 0 13616 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_144
timestamp 1676037725
transform 1 0 14352 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_155
timestamp 1676037725
transform 1 0 15364 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_168
timestamp 1676037725
transform 1 0 16560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_172
timestamp 1676037725
transform 1 0 16928 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_186
timestamp 1676037725
transform 1 0 18216 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_190
timestamp 1676037725
transform 1 0 18584 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1676037725
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_199
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_204
timestamp 1676037725
transform 1 0 19872 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_228
timestamp 1676037725
transform 1 0 22080 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_232
timestamp 1676037725
transform 1 0 22448 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1676037725
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_258
timestamp 1676037725
transform 1 0 24840 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_65
timestamp 1676037725
transform 1 0 7084 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_80
timestamp 1676037725
transform 1 0 8464 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_84
timestamp 1676037725
transform 1 0 8832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_95
timestamp 1676037725
transform 1 0 9844 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1676037725
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_115
timestamp 1676037725
transform 1 0 11684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_121
timestamp 1676037725
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_136
timestamp 1676037725
transform 1 0 13616 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_144
timestamp 1676037725
transform 1 0 14352 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1676037725
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1676037725
transform 1 0 17204 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_179
timestamp 1676037725
transform 1 0 17572 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_186
timestamp 1676037725
transform 1 0 18216 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_210
timestamp 1676037725
transform 1 0 20424 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_214
timestamp 1676037725
transform 1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_218
timestamp 1676037725
transform 1 0 21160 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_228
timestamp 1676037725
transform 1 0 22080 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_239
timestamp 1676037725
transform 1 0 23092 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_264
timestamp 1676037725
transform 1 0 25392 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_69
timestamp 1676037725
transform 1 0 7452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1676037725
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_90
timestamp 1676037725
transform 1 0 9384 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_117
timestamp 1676037725
transform 1 0 11868 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_130
timestamp 1676037725
transform 1 0 13064 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1676037725
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_143
timestamp 1676037725
transform 1 0 14260 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_155
timestamp 1676037725
transform 1 0 15364 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_159
timestamp 1676037725
transform 1 0 15732 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_173
timestamp 1676037725
transform 1 0 17020 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_186
timestamp 1676037725
transform 1 0 18216 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_208
timestamp 1676037725
transform 1 0 20240 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1676037725
transform 1 0 20884 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_222
timestamp 1676037725
transform 1 0 21528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_230
timestamp 1676037725
transform 1 0 22264 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1676037725
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_264
timestamp 1676037725
transform 1 0 25392 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1676037725
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1676037725
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1676037725
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1676037725
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1676037725
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_92
timestamp 1676037725
transform 1 0 9568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_121
timestamp 1676037725
transform 1 0 12236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_134
timestamp 1676037725
transform 1 0 13432 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_147
timestamp 1676037725
transform 1 0 14628 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_151
timestamp 1676037725
transform 1 0 14996 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1676037725
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_191
timestamp 1676037725
transform 1 0 18676 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_195
timestamp 1676037725
transform 1 0 19044 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_207
timestamp 1676037725
transform 1 0 20148 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_215
timestamp 1676037725
transform 1 0 20884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1676037725
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_244
timestamp 1676037725
transform 1 0 23552 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_264
timestamp 1676037725
transform 1 0 25392 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_59
timestamp 1676037725
transform 1 0 6532 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_80
timestamp 1676037725
transform 1 0 8464 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_95
timestamp 1676037725
transform 1 0 9844 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_106
timestamp 1676037725
transform 1 0 10856 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_110
timestamp 1676037725
transform 1 0 11224 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_122
timestamp 1676037725
transform 1 0 12328 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_135
timestamp 1676037725
transform 1 0 13524 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_146
timestamp 1676037725
transform 1 0 14536 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_158
timestamp 1676037725
transform 1 0 15640 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_170
timestamp 1676037725
transform 1 0 16744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_180
timestamp 1676037725
transform 1 0 17664 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_186
timestamp 1676037725
transform 1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1676037725
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_209
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_217
timestamp 1676037725
transform 1 0 21068 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_222
timestamp 1676037725
transform 1 0 21528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_226
timestamp 1676037725
transform 1 0 21896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_230
timestamp 1676037725
transform 1 0 22264 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_259
timestamp 1676037725
transform 1 0 24932 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_263
timestamp 1676037725
transform 1 0 25300 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_79
timestamp 1676037725
transform 1 0 8372 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_92
timestamp 1676037725
transform 1 0 9568 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_104
timestamp 1676037725
transform 1 0 10672 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_118
timestamp 1676037725
transform 1 0 11960 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1676037725
transform 1 0 14352 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_148
timestamp 1676037725
transform 1 0 14720 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_154
timestamp 1676037725
transform 1 0 15272 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_160
timestamp 1676037725
transform 1 0 15824 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1676037725
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_180
timestamp 1676037725
transform 1 0 17664 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_192
timestamp 1676037725
transform 1 0 18768 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_197
timestamp 1676037725
transform 1 0 19228 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_205
timestamp 1676037725
transform 1 0 19964 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1676037725
transform 1 0 20884 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1676037725
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_227
timestamp 1676037725
transform 1 0 21988 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1676037725
transform 1 0 23000 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_262
timestamp 1676037725
transform 1 0 25208 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_77
timestamp 1676037725
transform 1 0 8188 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_81
timestamp 1676037725
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_107
timestamp 1676037725
transform 1 0 10948 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_120
timestamp 1676037725
transform 1 0 12144 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_132
timestamp 1676037725
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_163
timestamp 1676037725
transform 1 0 16100 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_170
timestamp 1676037725
transform 1 0 16744 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_174
timestamp 1676037725
transform 1 0 17112 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_187
timestamp 1676037725
transform 1 0 18308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_203
timestamp 1676037725
transform 1 0 19780 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_224
timestamp 1676037725
transform 1 0 21712 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_248
timestamp 1676037725
transform 1 0 23920 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_255
timestamp 1676037725
transform 1 0 24564 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_263
timestamp 1676037725
transform 1 0 25300 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_95
timestamp 1676037725
transform 1 0 9844 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_99
timestamp 1676037725
transform 1 0 10212 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1676037725
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_146
timestamp 1676037725
transform 1 0 14536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_150
timestamp 1676037725
transform 1 0 14904 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_160
timestamp 1676037725
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1676037725
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_198
timestamp 1676037725
transform 1 0 19320 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1676037725
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_209
timestamp 1676037725
transform 1 0 20332 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_219
timestamp 1676037725
transform 1 0 21252 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_230
timestamp 1676037725
transform 1 0 22264 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_234
timestamp 1676037725
transform 1 0 22632 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_238
timestamp 1676037725
transform 1 0 23000 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_264
timestamp 1676037725
transform 1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1676037725
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_88
timestamp 1676037725
transform 1 0 9200 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_99
timestamp 1676037725
transform 1 0 10212 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_103
timestamp 1676037725
transform 1 0 10580 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_124
timestamp 1676037725
transform 1 0 12512 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_128
timestamp 1676037725
transform 1 0 12880 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1676037725
transform 1 0 14444 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_148
timestamp 1676037725
transform 1 0 14720 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_152
timestamp 1676037725
transform 1 0 15088 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_173
timestamp 1676037725
transform 1 0 17020 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1676037725
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_189
timestamp 1676037725
transform 1 0 18492 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1676037725
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_208
timestamp 1676037725
transform 1 0 20240 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1676037725
transform 1 0 20608 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_217
timestamp 1676037725
transform 1 0 21068 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_223
timestamp 1676037725
transform 1 0 21620 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_230
timestamp 1676037725
transform 1 0 22264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_250
timestamp 1676037725
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_264
timestamp 1676037725
transform 1 0 25392 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1676037725
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1676037725
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1676037725
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_83
timestamp 1676037725
transform 1 0 8740 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_87
timestamp 1676037725
transform 1 0 9108 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_97
timestamp 1676037725
transform 1 0 10028 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1676037725
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_118
timestamp 1676037725
transform 1 0 11960 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_150
timestamp 1676037725
transform 1 0 14904 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_154
timestamp 1676037725
transform 1 0 15272 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1676037725
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1676037725
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_181
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_189
timestamp 1676037725
transform 1 0 18492 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_194
timestamp 1676037725
transform 1 0 18952 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_198
timestamp 1676037725
transform 1 0 19320 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_209
timestamp 1676037725
transform 1 0 20332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_216
timestamp 1676037725
transform 1 0 20976 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_236
timestamp 1676037725
transform 1 0 22816 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_240
timestamp 1676037725
transform 1 0 23184 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_261
timestamp 1676037725
transform 1 0 25116 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_265
timestamp 1676037725
transform 1 0 25484 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1676037725
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1676037725
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_87
timestamp 1676037725
transform 1 0 9108 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_99
timestamp 1676037725
transform 1 0 10212 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_102
timestamp 1676037725
transform 1 0 10488 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_113
timestamp 1676037725
transform 1 0 11500 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_117
timestamp 1676037725
transform 1 0 11868 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_127
timestamp 1676037725
transform 1 0 12788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1676037725
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_158
timestamp 1676037725
transform 1 0 15640 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_162
timestamp 1676037725
transform 1 0 16008 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_183
timestamp 1676037725
transform 1 0 17940 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_187
timestamp 1676037725
transform 1 0 18308 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1676037725
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_201
timestamp 1676037725
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_211
timestamp 1676037725
transform 1 0 20516 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_218
timestamp 1676037725
transform 1 0 21160 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_242
timestamp 1676037725
transform 1 0 23368 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_249
timestamp 1676037725
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_264
timestamp 1676037725
transform 1 0 25392 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1676037725
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1676037725
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_75
timestamp 1676037725
transform 1 0 8004 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_96
timestamp 1676037725
transform 1 0 9936 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_100
timestamp 1676037725
transform 1 0 10304 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_121
timestamp 1676037725
transform 1 0 12236 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_142
timestamp 1676037725
transform 1 0 14168 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_148
timestamp 1676037725
transform 1 0 14720 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_160
timestamp 1676037725
transform 1 0 15824 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_174
timestamp 1676037725
transform 1 0 17112 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_186
timestamp 1676037725
transform 1 0 18216 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_190
timestamp 1676037725
transform 1 0 18584 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_195
timestamp 1676037725
transform 1 0 19044 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_201
timestamp 1676037725
transform 1 0 19596 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_205
timestamp 1676037725
transform 1 0 19964 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_211
timestamp 1676037725
transform 1 0 20516 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_244
timestamp 1676037725
transform 1 0 23552 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_264
timestamp 1676037725
transform 1 0 25392 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1676037725
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1676037725
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_96
timestamp 1676037725
transform 1 0 9936 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_100
timestamp 1676037725
transform 1 0 10304 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_108
timestamp 1676037725
transform 1 0 11040 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_119
timestamp 1676037725
transform 1 0 12052 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_127
timestamp 1676037725
transform 1 0 12788 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_143
timestamp 1676037725
transform 1 0 14260 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_146
timestamp 1676037725
transform 1 0 14536 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_157
timestamp 1676037725
transform 1 0 15548 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_161
timestamp 1676037725
transform 1 0 15916 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_173
timestamp 1676037725
transform 1 0 17020 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_181
timestamp 1676037725
transform 1 0 17756 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_191
timestamp 1676037725
transform 1 0 18676 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1676037725
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_216
timestamp 1676037725
transform 1 0 20976 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_222
timestamp 1676037725
transform 1 0 21528 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_226
timestamp 1676037725
transform 1 0 21896 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1676037725
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1676037725
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_95
timestamp 1676037725
transform 1 0 9844 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_99
timestamp 1676037725
transform 1 0 10212 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1676037725
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_131
timestamp 1676037725
transform 1 0 13156 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_141
timestamp 1676037725
transform 1 0 14076 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_154
timestamp 1676037725
transform 1 0 15272 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1676037725
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1676037725
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1676037725
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_187
timestamp 1676037725
transform 1 0 18308 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_195
timestamp 1676037725
transform 1 0 19044 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_206
timestamp 1676037725
transform 1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_219
timestamp 1676037725
transform 1 0 21252 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1676037725
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_232
timestamp 1676037725
transform 1 0 22448 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_260
timestamp 1676037725
transform 1 0 25024 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1676037725
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1676037725
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_107
timestamp 1676037725
transform 1 0 10948 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_114
timestamp 1676037725
transform 1 0 11592 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1676037725
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_143
timestamp 1676037725
transform 1 0 14260 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_155
timestamp 1676037725
transform 1 0 15364 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_181
timestamp 1676037725
transform 1 0 17756 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1676037725
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_219
timestamp 1676037725
transform 1 0 21252 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_224
timestamp 1676037725
transform 1 0 21712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_246
timestamp 1676037725
transform 1 0 23736 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1676037725
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_258
timestamp 1676037725
transform 1 0 24840 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1676037725
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1676037725
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1676037725
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_81
timestamp 1676037725
transform 1 0 8556 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_89
timestamp 1676037725
transform 1 0 9292 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1676037725
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_124
timestamp 1676037725
transform 1 0 12512 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_128
timestamp 1676037725
transform 1 0 12880 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_149
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_158
timestamp 1676037725
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1676037725
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_180
timestamp 1676037725
transform 1 0 17664 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_193
timestamp 1676037725
transform 1 0 18860 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_199
timestamp 1676037725
transform 1 0 19412 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1676037725
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_237
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1676037725
transform 1 0 23460 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_264
timestamp 1676037725
transform 1 0 25392 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1676037725
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1676037725
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_105
timestamp 1676037725
transform 1 0 10764 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_126
timestamp 1676037725
transform 1 0 12696 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_130
timestamp 1676037725
transform 1 0 13064 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_138
timestamp 1676037725
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_152
timestamp 1676037725
transform 1 0 15088 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_156
timestamp 1676037725
transform 1 0 15456 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_168
timestamp 1676037725
transform 1 0 16560 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_175
timestamp 1676037725
transform 1 0 17204 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_182
timestamp 1676037725
transform 1 0 17848 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_188
timestamp 1676037725
transform 1 0 18400 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1676037725
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_199
timestamp 1676037725
transform 1 0 19412 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_206
timestamp 1676037725
transform 1 0 20056 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_210
timestamp 1676037725
transform 1 0 20424 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_217
timestamp 1676037725
transform 1 0 21068 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_221
timestamp 1676037725
transform 1 0 21436 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_225
timestamp 1676037725
transform 1 0 21804 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_233
timestamp 1676037725
transform 1 0 22540 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1676037725
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_259
timestamp 1676037725
transform 1 0 24932 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_264
timestamp 1676037725
transform 1 0 25392 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1676037725
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1676037725
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1676037725
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1676037725
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1676037725
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_119
timestamp 1676037725
transform 1 0 12052 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_129
timestamp 1676037725
transform 1 0 12972 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_144
timestamp 1676037725
transform 1 0 14352 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_148
timestamp 1676037725
transform 1 0 14720 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_158
timestamp 1676037725
transform 1 0 15640 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1676037725
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_174
timestamp 1676037725
transform 1 0 17112 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_178
timestamp 1676037725
transform 1 0 17480 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_190
timestamp 1676037725
transform 1 0 18584 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_194
timestamp 1676037725
transform 1 0 18952 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_197
timestamp 1676037725
transform 1 0 19228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_209
timestamp 1676037725
transform 1 0 20332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_221
timestamp 1676037725
transform 1 0 21436 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_236
timestamp 1676037725
transform 1 0 22816 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_240
timestamp 1676037725
transform 1 0 23184 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_244
timestamp 1676037725
transform 1 0 23552 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_264
timestamp 1676037725
transform 1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_107
timestamp 1676037725
transform 1 0 10948 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_113
timestamp 1676037725
transform 1 0 11500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_125
timestamp 1676037725
transform 1 0 12604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1676037725
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_152
timestamp 1676037725
transform 1 0 15088 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_156
timestamp 1676037725
transform 1 0 15456 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_167
timestamp 1676037725
transform 1 0 16468 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_177
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_185
timestamp 1676037725
transform 1 0 18124 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1676037725
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_219
timestamp 1676037725
transform 1 0 21252 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_223
timestamp 1676037725
transform 1 0 21620 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_229
timestamp 1676037725
transform 1 0 22172 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_232
timestamp 1676037725
transform 1 0 22448 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_243
timestamp 1676037725
transform 1 0 23460 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1676037725
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_264
timestamp 1676037725
transform 1 0 25392 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1676037725
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1676037725
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1676037725
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_81
timestamp 1676037725
transform 1 0 8556 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp 1676037725
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_115
timestamp 1676037725
transform 1 0 11684 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_127
timestamp 1676037725
transform 1 0 12788 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_150
timestamp 1676037725
transform 1 0 14904 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_163
timestamp 1676037725
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1676037725
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_203
timestamp 1676037725
transform 1 0 19780 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_207
timestamp 1676037725
transform 1 0 20148 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1676037725
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1676037725
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_227
timestamp 1676037725
transform 1 0 21988 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_240
timestamp 1676037725
transform 1 0 23184 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_264
timestamp 1676037725
transform 1 0 25392 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_101
timestamp 1676037725
transform 1 0 10396 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_122
timestamp 1676037725
transform 1 0 12328 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_126
timestamp 1676037725
transform 1 0 12696 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1676037725
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_162
timestamp 1676037725
transform 1 0 16008 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_168
timestamp 1676037725
transform 1 0 16560 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_176
timestamp 1676037725
transform 1 0 17296 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_187
timestamp 1676037725
transform 1 0 18308 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_203
timestamp 1676037725
transform 1 0 19780 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_224
timestamp 1676037725
transform 1 0 21712 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_248
timestamp 1676037725
transform 1 0 23920 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_264
timestamp 1676037725
transform 1 0 25392 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1676037725
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1676037725
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1676037725
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1676037725
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1676037725
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_105
timestamp 1676037725
transform 1 0 10764 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_109
timestamp 1676037725
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_135
timestamp 1676037725
transform 1 0 13524 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_139
timestamp 1676037725
transform 1 0 13892 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_151
timestamp 1676037725
transform 1 0 14996 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_162
timestamp 1676037725
transform 1 0 16008 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_180
timestamp 1676037725
transform 1 0 17664 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_187
timestamp 1676037725
transform 1 0 18308 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_196
timestamp 1676037725
transform 1 0 19136 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_200
timestamp 1676037725
transform 1 0 19504 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_205
timestamp 1676037725
transform 1 0 19964 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_220
timestamp 1676037725
transform 1 0 21344 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_236
timestamp 1676037725
transform 1 0 22816 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_260
timestamp 1676037725
transform 1 0 25024 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_107
timestamp 1676037725
transform 1 0 10948 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_111
timestamp 1676037725
transform 1 0 11316 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_132
timestamp 1676037725
transform 1 0 13248 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1676037725
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_158
timestamp 1676037725
transform 1 0 15640 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_166
timestamp 1676037725
transform 1 0 16376 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_194
timestamp 1676037725
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_208
timestamp 1676037725
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_232
timestamp 1676037725
transform 1 0 22448 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_245
timestamp 1676037725
transform 1 0 23644 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1676037725
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_264
timestamp 1676037725
transform 1 0 25392 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_81
timestamp 1676037725
transform 1 0 8556 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_89
timestamp 1676037725
transform 1 0 9292 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_100
timestamp 1676037725
transform 1 0 10304 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_119
timestamp 1676037725
transform 1 0 12052 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_129
timestamp 1676037725
transform 1 0 12972 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_153
timestamp 1676037725
transform 1 0 15180 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1676037725
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_180
timestamp 1676037725
transform 1 0 17664 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_186
timestamp 1676037725
transform 1 0 18216 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_201
timestamp 1676037725
transform 1 0 19596 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_207
timestamp 1676037725
transform 1 0 20148 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_219
timestamp 1676037725
transform 1 0 21252 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1676037725
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_227
timestamp 1676037725
transform 1 0 21988 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_240
timestamp 1676037725
transform 1 0 23184 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_253
timestamp 1676037725
transform 1 0 24380 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_260
timestamp 1676037725
transform 1 0 25024 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1676037725
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_129
timestamp 1676037725
transform 1 0 12972 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_135
timestamp 1676037725
transform 1 0 13524 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1676037725
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_162
timestamp 1676037725
transform 1 0 16008 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_168
timestamp 1676037725
transform 1 0 16560 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_172
timestamp 1676037725
transform 1 0 16928 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_193
timestamp 1676037725
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_202
timestamp 1676037725
transform 1 0 19688 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_206
timestamp 1676037725
transform 1 0 20056 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_216
timestamp 1676037725
transform 1 0 20976 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_228
timestamp 1676037725
transform 1 0 22080 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_238
timestamp 1676037725
transform 1 0 23000 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_243
timestamp 1676037725
transform 1 0 23460 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_250
timestamp 1676037725
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_255
timestamp 1676037725
transform 1 0 24564 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_259
timestamp 1676037725
transform 1 0 24932 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_264
timestamp 1676037725
transform 1 0 25392 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1676037725
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1676037725
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_81
timestamp 1676037725
transform 1 0 8556 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_88
timestamp 1676037725
transform 1 0 9200 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_100
timestamp 1676037725
transform 1 0 10304 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_136
timestamp 1676037725
transform 1 0 13616 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_140
timestamp 1676037725
transform 1 0 13984 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_152
timestamp 1676037725
transform 1 0 15088 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_51_165
timestamp 1676037725
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_173
timestamp 1676037725
transform 1 0 17020 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_185
timestamp 1676037725
transform 1 0 18124 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_195
timestamp 1676037725
transform 1 0 19044 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_203
timestamp 1676037725
transform 1 0 19780 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_213
timestamp 1676037725
transform 1 0 20700 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_51_222
timestamp 1676037725
transform 1 0 21528 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_236
timestamp 1676037725
transform 1 0 22816 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_240
timestamp 1676037725
transform 1 0 23184 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_261
timestamp 1676037725
transform 1 0 25116 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_265
timestamp 1676037725
transform 1 0 25484 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1676037725
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_90
timestamp 1676037725
transform 1 0 9384 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_102
timestamp 1676037725
transform 1 0 10488 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_114
timestamp 1676037725
transform 1 0 11592 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_126
timestamp 1676037725
transform 1 0 12696 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1676037725
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_155
timestamp 1676037725
transform 1 0 15364 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_161
timestamp 1676037725
transform 1 0 15916 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_169
timestamp 1676037725
transform 1 0 16652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_190
timestamp 1676037725
transform 1 0 18584 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1676037725
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_205
timestamp 1676037725
transform 1 0 19964 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_209
timestamp 1676037725
transform 1 0 20332 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_233
timestamp 1676037725
transform 1 0 22540 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_237
timestamp 1676037725
transform 1 0 22908 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1676037725
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_258
timestamp 1676037725
transform 1 0 24840 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1676037725
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1676037725
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1676037725
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1676037725
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1676037725
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1676037725
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_154
timestamp 1676037725
transform 1 0 15272 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_160
timestamp 1676037725
transform 1 0 15824 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_171
timestamp 1676037725
transform 1 0 16836 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_197
timestamp 1676037725
transform 1 0 19228 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_201
timestamp 1676037725
transform 1 0 19596 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_204
timestamp 1676037725
transform 1 0 19872 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_215
timestamp 1676037725
transform 1 0 20884 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1676037725
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_231
timestamp 1676037725
transform 1 0 22356 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_252
timestamp 1676037725
transform 1 0 24288 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_256
timestamp 1676037725
transform 1 0 24656 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_260
timestamp 1676037725
transform 1 0 25024 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_264
timestamp 1676037725
transform 1 0 25392 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1676037725
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1676037725
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1676037725
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1676037725
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_153
timestamp 1676037725
transform 1 0 15180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_166
timestamp 1676037725
transform 1 0 16376 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_190
timestamp 1676037725
transform 1 0 18584 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_194
timestamp 1676037725
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_219
timestamp 1676037725
transform 1 0 21252 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_232
timestamp 1676037725
transform 1 0 22448 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_236
timestamp 1676037725
transform 1 0 22816 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_247
timestamp 1676037725
transform 1 0 23828 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1676037725
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_259
timestamp 1676037725
transform 1 0 24932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_264
timestamp 1676037725
transform 1 0 25392 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1676037725
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1676037725
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1676037725
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1676037725
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1676037725
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1676037725
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1676037725
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_149
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1676037725
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_174
timestamp 1676037725
transform 1 0 17112 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_186
timestamp 1676037725
transform 1 0 18216 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_194
timestamp 1676037725
transform 1 0 18952 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_215
timestamp 1676037725
transform 1 0 20884 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_219
timestamp 1676037725
transform 1 0 21252 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_239
timestamp 1676037725
transform 1 0 23092 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_55_263
timestamp 1676037725
transform 1 0 25300 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1676037725
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1676037725
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1676037725
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1676037725
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1676037725
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1676037725
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1676037725
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_166
timestamp 1676037725
transform 1 0 16376 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_174
timestamp 1676037725
transform 1 0 17112 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_186
timestamp 1676037725
transform 1 0 18216 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1676037725
transform 1 0 18952 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_202
timestamp 1676037725
transform 1 0 19688 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_215
timestamp 1676037725
transform 1 0 20884 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_227
timestamp 1676037725
transform 1 0 21988 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1676037725
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_264
timestamp 1676037725
transform 1 0 25392 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1676037725
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1676037725
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1676037725
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1676037725
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1676037725
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1676037725
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1676037725
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1676037725
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1676037725
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_193
timestamp 1676037725
transform 1 0 18860 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_199
timestamp 1676037725
transform 1 0 19412 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_220
timestamp 1676037725
transform 1 0 21344 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_247
timestamp 1676037725
transform 1 0 23828 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_57_256
timestamp 1676037725
transform 1 0 24656 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_259
timestamp 1676037725
transform 1 0 24932 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_264
timestamp 1676037725
transform 1 0 25392 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1676037725
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1676037725
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1676037725
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1676037725
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_90
timestamp 1676037725
transform 1 0 9384 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_102
timestamp 1676037725
transform 1 0 10488 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_114
timestamp 1676037725
transform 1 0 11592 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_126
timestamp 1676037725
transform 1 0 12696 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_138
timestamp 1676037725
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_158
timestamp 1676037725
transform 1 0 15640 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_162
timestamp 1676037725
transform 1 0 16008 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_174
timestamp 1676037725
transform 1 0 17112 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_186
timestamp 1676037725
transform 1 0 18216 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_194
timestamp 1676037725
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_219
timestamp 1676037725
transform 1 0 21252 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_243
timestamp 1676037725
transform 1 0 23460 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_247
timestamp 1676037725
transform 1 0 23828 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1676037725
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_259
timestamp 1676037725
transform 1 0 24932 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_264
timestamp 1676037725
transform 1 0 25392 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1676037725
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1676037725
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1676037725
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1676037725
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1676037725
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1676037725
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1676037725
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1676037725
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1676037725
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1676037725
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1676037725
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1676037725
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1676037725
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1676037725
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1676037725
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_217
timestamp 1676037725
transform 1 0 21068 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_221
timestamp 1676037725
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1676037725
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_249
timestamp 1676037725
transform 1 0 24012 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_259
timestamp 1676037725
transform 1 0 24932 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_264
timestamp 1676037725
transform 1 0 25392 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1676037725
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1676037725
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1676037725
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1676037725
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1676037725
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1676037725
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1676037725
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1676037725
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1676037725
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1676037725
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1676037725
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_221
timestamp 1676037725
transform 1 0 21436 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_227
timestamp 1676037725
transform 1 0 21988 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_233
timestamp 1676037725
transform 1 0 22540 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_244
timestamp 1676037725
transform 1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_264
timestamp 1676037725
transform 1 0 25392 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1676037725
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1676037725
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1676037725
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1676037725
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_81
timestamp 1676037725
transform 1 0 8556 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_89
timestamp 1676037725
transform 1 0 9292 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1676037725
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_117
timestamp 1676037725
transform 1 0 11868 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_129
timestamp 1676037725
transform 1 0 12972 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_141
timestamp 1676037725
transform 1 0 14076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_153
timestamp 1676037725
transform 1 0 15180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_165
timestamp 1676037725
transform 1 0 16284 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1676037725
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1676037725
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_205
timestamp 1676037725
transform 1 0 19964 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_211
timestamp 1676037725
transform 1 0 20516 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1676037725
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_236
timestamp 1676037725
transform 1 0 22816 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_248
timestamp 1676037725
transform 1 0 23920 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_260
timestamp 1676037725
transform 1 0 25024 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1676037725
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1676037725
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1676037725
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1676037725
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1676037725
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1676037725
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1676037725
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1676037725
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1676037725
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1676037725
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1676037725
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1676037725
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1676037725
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1676037725
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1676037725
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1676037725
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1676037725
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1676037725
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_259
timestamp 1676037725
transform 1 0 24932 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_264
timestamp 1676037725
transform 1 0 25392 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1676037725
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1676037725
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1676037725
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1676037725
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1676037725
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1676037725
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1676037725
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1676037725
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1676037725
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1676037725
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1676037725
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1676037725
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1676037725
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1676037725
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1676037725
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1676037725
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1676037725
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1676037725
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1676037725
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_249
timestamp 1676037725
transform 1 0 24012 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_257
timestamp 1676037725
transform 1 0 24748 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_264
timestamp 1676037725
transform 1 0 25392 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1676037725
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1676037725
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1676037725
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1676037725
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1676037725
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1676037725
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1676037725
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1676037725
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1676037725
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1676037725
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1676037725
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1676037725
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1676037725
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1676037725
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1676037725
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1676037725
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1676037725
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1676037725
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_261
timestamp 1676037725
transform 1 0 25116 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1676037725
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1676037725
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1676037725
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1676037725
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1676037725
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_81
timestamp 1676037725
transform 1 0 8556 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_85
timestamp 1676037725
transform 1 0 8924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_97
timestamp 1676037725
transform 1 0 10028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_109
timestamp 1676037725
transform 1 0 11132 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1676037725
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1676037725
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1676037725
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1676037725
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1676037725
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1676037725
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1676037725
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1676037725
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1676037725
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1676037725
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_249
timestamp 1676037725
transform 1 0 24012 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_255
timestamp 1676037725
transform 1 0 24564 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_258
timestamp 1676037725
transform 1 0 24840 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_264
timestamp 1676037725
transform 1 0 25392 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1676037725
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1676037725
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1676037725
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1676037725
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1676037725
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1676037725
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1676037725
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1676037725
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1676037725
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1676037725
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1676037725
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1676037725
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1676037725
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1676037725
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1676037725
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1676037725
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1676037725
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1676037725
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1676037725
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_264
timestamp 1676037725
transform 1 0 25392 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1676037725
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1676037725
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1676037725
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1676037725
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1676037725
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1676037725
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1676037725
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1676037725
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1676037725
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1676037725
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1676037725
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1676037725
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1676037725
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1676037725
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1676037725
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1676037725
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1676037725
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1676037725
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_261
timestamp 1676037725
transform 1 0 25116 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1676037725
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1676037725
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1676037725
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1676037725
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1676037725
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1676037725
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1676037725
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1676037725
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1676037725
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1676037725
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1676037725
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1676037725
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1676037725
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1676037725
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1676037725
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1676037725
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1676037725
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_259
timestamp 1676037725
transform 1 0 24932 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_264
timestamp 1676037725
transform 1 0 25392 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1676037725
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1676037725
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1676037725
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1676037725
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1676037725
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1676037725
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1676037725
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1676037725
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1676037725
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1676037725
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1676037725
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1676037725
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1676037725
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1676037725
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1676037725
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1676037725
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1676037725
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1676037725
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1676037725
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1676037725
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1676037725
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_264
timestamp 1676037725
transform 1 0 25392 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1676037725
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1676037725
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1676037725
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1676037725
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1676037725
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1676037725
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1676037725
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1676037725
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1676037725
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1676037725
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1676037725
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1676037725
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1676037725
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1676037725
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1676037725
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1676037725
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_253
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_261
timestamp 1676037725
transform 1 0 25116 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1676037725
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1676037725
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1676037725
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1676037725
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1676037725
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1676037725
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1676037725
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1676037725
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1676037725
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1676037725
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1676037725
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1676037725
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1676037725
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1676037725
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1676037725
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1676037725
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1676037725
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1676037725
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1676037725
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1676037725
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_249
timestamp 1676037725
transform 1 0 24012 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_259
timestamp 1676037725
transform 1 0 24932 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_264
timestamp 1676037725
transform 1 0 25392 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1676037725
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1676037725
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1676037725
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1676037725
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1676037725
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_107
timestamp 1676037725
transform 1 0 10948 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_119
timestamp 1676037725
transform 1 0 12052 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_131
timestamp 1676037725
transform 1 0 13156 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1676037725
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1676037725
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1676037725
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1676037725
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1676037725
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1676037725
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1676037725
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1676037725
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1676037725
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1676037725
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_259
timestamp 1676037725
transform 1 0 24932 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_264
timestamp 1676037725
transform 1 0 25392 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1676037725
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1676037725
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1676037725
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1676037725
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1676037725
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_81
timestamp 1676037725
transform 1 0 8556 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_89
timestamp 1676037725
transform 1 0 9292 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_110
timestamp 1676037725
transform 1 0 11224 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_117
timestamp 1676037725
transform 1 0 11868 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_129
timestamp 1676037725
transform 1 0 12972 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_141
timestamp 1676037725
transform 1 0 14076 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_153
timestamp 1676037725
transform 1 0 15180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_165
timestamp 1676037725
transform 1 0 16284 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1676037725
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1676037725
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1676037725
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1676037725
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1676037725
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1676037725
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1676037725
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_261
timestamp 1676037725
transform 1 0 25116 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1676037725
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1676037725
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1676037725
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1676037725
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1676037725
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1676037725
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_85
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_91
timestamp 1676037725
transform 1 0 9476 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_100
timestamp 1676037725
transform 1 0 10304 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_112
timestamp 1676037725
transform 1 0 11408 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_124
timestamp 1676037725
transform 1 0 12512 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_136
timestamp 1676037725
transform 1 0 13616 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1676037725
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1676037725
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1676037725
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1676037725
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1676037725
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1676037725
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1676037725
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1676037725
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1676037725
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1676037725
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_253
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_258
timestamp 1676037725
transform 1 0 24840 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_264
timestamp 1676037725
transform 1 0 25392 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1676037725
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1676037725
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1676037725
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1676037725
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1676037725
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1676037725
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1676037725
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1676037725
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1676037725
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1676037725
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1676037725
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1676037725
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1676037725
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1676037725
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1676037725
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1676037725
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1676037725
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1676037725
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1676037725
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1676037725
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_249
timestamp 1676037725
transform 1 0 24012 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_257
timestamp 1676037725
transform 1 0 24748 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_264
timestamp 1676037725
transform 1 0 25392 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1676037725
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1676037725
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1676037725
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1676037725
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1676037725
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1676037725
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1676037725
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1676037725
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1676037725
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1676037725
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1676037725
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1676037725
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1676037725
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1676037725
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1676037725
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1676037725
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_229
timestamp 1676037725
transform 1 0 22172 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1676037725
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1676037725
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1676037725
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_261
timestamp 1676037725
transform 1 0 25116 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1676037725
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1676037725
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1676037725
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1676037725
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1676037725
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1676037725
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_81
timestamp 1676037725
transform 1 0 8556 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_93
timestamp 1676037725
transform 1 0 9660 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_101
timestamp 1676037725
transform 1 0 10396 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_77_109
timestamp 1676037725
transform 1 0 11132 0 -1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_77_115
timestamp 1676037725
transform 1 0 11684 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_127
timestamp 1676037725
transform 1 0 12788 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_139
timestamp 1676037725
transform 1 0 13892 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_151
timestamp 1676037725
transform 1 0 14996 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_163
timestamp 1676037725
transform 1 0 16100 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1676037725
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1676037725
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1676037725
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1676037725
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1676037725
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1676037725
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1676037725
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_249
timestamp 1676037725
transform 1 0 24012 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_255
timestamp 1676037725
transform 1 0 24564 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_258
timestamp 1676037725
transform 1 0 24840 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_264
timestamp 1676037725
transform 1 0 25392 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1676037725
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1676037725
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1676037725
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_107
timestamp 1676037725
transform 1 0 10948 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_113
timestamp 1676037725
transform 1 0 11500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_125
timestamp 1676037725
transform 1 0 12604 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_137
timestamp 1676037725
transform 1 0 13708 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_153
timestamp 1676037725
transform 1 0 15180 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_157
timestamp 1676037725
transform 1 0 15548 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_179
timestamp 1676037725
transform 1 0 17572 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_191
timestamp 1676037725
transform 1 0 18676 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1676037725
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1676037725
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1676037725
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1676037725
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1676037725
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1676037725
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_253
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_264
timestamp 1676037725
transform 1 0 25392 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1676037725
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1676037725
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1676037725
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1676037725
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1676037725
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1676037725
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1676037725
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1676037725
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1676037725
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1676037725
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_125
timestamp 1676037725
transform 1 0 12604 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_147
timestamp 1676037725
transform 1 0 14628 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_159
timestamp 1676037725
transform 1 0 15732 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1676037725
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1676037725
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1676037725
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1676037725
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1676037725
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1676037725
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1676037725
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1676037725
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_261
timestamp 1676037725
transform 1 0 25116 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1676037725
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_73
timestamp 1676037725
transform 1 0 7820 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_82
timestamp 1676037725
transform 1 0 8648 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1676037725
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_121
timestamp 1676037725
transform 1 0 12236 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_129
timestamp 1676037725
transform 1 0 12972 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_135
timestamp 1676037725
transform 1 0 13524 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1676037725
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_141
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_170
timestamp 1676037725
transform 1 0 16744 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_182
timestamp 1676037725
transform 1 0 17848 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_194
timestamp 1676037725
transform 1 0 18952 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1676037725
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1676037725
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1676037725
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1676037725
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1676037725
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_253
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_259
timestamp 1676037725
transform 1 0 24932 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_264
timestamp 1676037725
transform 1 0 25392 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1676037725
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1676037725
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1676037725
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1676037725
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1676037725
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1676037725
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1676037725
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_93
timestamp 1676037725
transform 1 0 9660 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_99
timestamp 1676037725
transform 1 0 10212 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_106
timestamp 1676037725
transform 1 0 10856 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_110
timestamp 1676037725
transform 1 0 11224 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_121
timestamp 1676037725
transform 1 0 12236 0 -1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_127
timestamp 1676037725
transform 1 0 12788 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_160
timestamp 1676037725
transform 1 0 15824 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1676037725
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1676037725
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1676037725
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1676037725
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1676037725
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1676037725
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1676037725
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_264
timestamp 1676037725
transform 1 0 25392 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1676037725
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1676037725
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_109
timestamp 1676037725
transform 1 0 11132 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_113
timestamp 1676037725
transform 1 0 11500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_117
timestamp 1676037725
transform 1 0 11868 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_129
timestamp 1676037725
transform 1 0 12972 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_137
timestamp 1676037725
transform 1 0 13708 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1676037725
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1676037725
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1676037725
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1676037725
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1676037725
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1676037725
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1676037725
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1676037725
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1676037725
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1676037725
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_261
timestamp 1676037725
transform 1 0 25116 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1676037725
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1676037725
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1676037725
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1676037725
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1676037725
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_89
timestamp 1676037725
transform 1 0 9292 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_96
timestamp 1676037725
transform 1 0 9936 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_100
timestamp 1676037725
transform 1 0 10304 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1676037725
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1676037725
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1676037725
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1676037725
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1676037725
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1676037725
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1676037725
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1676037725
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1676037725
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1676037725
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1676037725
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_249
timestamp 1676037725
transform 1 0 24012 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_259
timestamp 1676037725
transform 1 0 24932 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_264
timestamp 1676037725
transform 1 0 25392 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1676037725
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1676037725
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_84_103
timestamp 1676037725
transform 1 0 10580 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_115
timestamp 1676037725
transform 1 0 11684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_127
timestamp 1676037725
transform 1 0 12788 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1676037725
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1676037725
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1676037725
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1676037725
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1676037725
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1676037725
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1676037725
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1676037725
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_233
timestamp 1676037725
transform 1 0 22540 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_241
timestamp 1676037725
transform 1 0 23276 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_250
timestamp 1676037725
transform 1 0 24104 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_84_253
timestamp 1676037725
transform 1 0 24380 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_259
timestamp 1676037725
transform 1 0 24932 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_264
timestamp 1676037725
transform 1 0 25392 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1676037725
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1676037725
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1676037725
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1676037725
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1676037725
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_85_80
timestamp 1676037725
transform 1 0 8464 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_86
timestamp 1676037725
transform 1 0 9016 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_98
timestamp 1676037725
transform 1 0 10120 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_110
timestamp 1676037725
transform 1 0 11224 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1676037725
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1676037725
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1676037725
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1676037725
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1676037725
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1676037725
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1676037725
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1676037725
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1676037725
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_261
timestamp 1676037725
transform 1 0 25116 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1676037725
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1676037725
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1676037725
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1676037725
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1676037725
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1676037725
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_97
timestamp 1676037725
transform 1 0 10028 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_105
timestamp 1676037725
transform 1 0 10764 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_111
timestamp 1676037725
transform 1 0 11316 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_116
timestamp 1676037725
transform 1 0 11776 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_128
timestamp 1676037725
transform 1 0 12880 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1676037725
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1676037725
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1676037725
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1676037725
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1676037725
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1676037725
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1676037725
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1676037725
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1676037725
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1676037725
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_86_253
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_86_258
timestamp 1676037725
transform 1 0 24840 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_264
timestamp 1676037725
transform 1 0 25392 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1676037725
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1676037725
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1676037725
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1676037725
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1676037725
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1676037725
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1676037725
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1676037725
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1676037725
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1676037725
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1676037725
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1676037725
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1676037725
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1676037725
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1676037725
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1676037725
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1676037725
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1676037725
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1676037725
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1676037725
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1676037725
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_249
timestamp 1676037725
transform 1 0 24012 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_253
timestamp 1676037725
transform 1 0 24380 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_264
timestamp 1676037725
transform 1 0 25392 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1676037725
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1676037725
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1676037725
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1676037725
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1676037725
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_65
timestamp 1676037725
transform 1 0 7084 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_69
timestamp 1676037725
transform 1 0 7452 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_88_76
timestamp 1676037725
transform 1 0 8096 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_80
timestamp 1676037725
transform 1 0 8464 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_89
timestamp 1676037725
transform 1 0 9292 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_94
timestamp 1676037725
transform 1 0 9752 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_106
timestamp 1676037725
transform 1 0 10856 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_118
timestamp 1676037725
transform 1 0 11960 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_130
timestamp 1676037725
transform 1 0 13064 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_138
timestamp 1676037725
transform 1 0 13800 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1676037725
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1676037725
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1676037725
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1676037725
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1676037725
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1676037725
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1676037725
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1676037725
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1676037725
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1676037725
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_88_261
timestamp 1676037725
transform 1 0 25116 0 1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1676037725
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1676037725
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1676037725
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1676037725
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1676037725
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1676037725
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1676037725
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1676037725
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1676037725
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1676037725
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1676037725
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1676037725
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1676037725
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1676037725
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1676037725
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1676037725
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1676037725
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1676037725
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1676037725
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1676037725
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_249
timestamp 1676037725
transform 1 0 24012 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_253
timestamp 1676037725
transform 1 0 24380 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_256
timestamp 1676037725
transform 1 0 24656 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_264
timestamp 1676037725
transform 1 0 25392 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1676037725
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1676037725
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1676037725
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1676037725
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_65
timestamp 1676037725
transform 1 0 7084 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_69
timestamp 1676037725
transform 1 0 7452 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_74
timestamp 1676037725
transform 1 0 7912 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_90_81
timestamp 1676037725
transform 1 0 8556 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_91
timestamp 1676037725
transform 1 0 9476 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_103
timestamp 1676037725
transform 1 0 10580 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_115
timestamp 1676037725
transform 1 0 11684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_127
timestamp 1676037725
transform 1 0 12788 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1676037725
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1676037725
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1676037725
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1676037725
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1676037725
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1676037725
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1676037725
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1676037725
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1676037725
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1676037725
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_90_253
timestamp 1676037725
transform 1 0 24380 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_90_256
timestamp 1676037725
transform 1 0 24656 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_264
timestamp 1676037725
transform 1 0 25392 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1676037725
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1676037725
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1676037725
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1676037725
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1676037725
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1676037725
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1676037725
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1676037725
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1676037725
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1676037725
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1676037725
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1676037725
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1676037725
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1676037725
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1676037725
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1676037725
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1676037725
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1676037725
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1676037725
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_249
timestamp 1676037725
transform 1 0 24012 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_259
timestamp 1676037725
transform 1 0 24932 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_264
timestamp 1676037725
transform 1 0 25392 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1676037725
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1676037725
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1676037725
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_53
timestamp 1676037725
transform 1 0 5980 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_62
timestamp 1676037725
transform 1 0 6808 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_74
timestamp 1676037725
transform 1 0 7912 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_82
timestamp 1676037725
transform 1 0 8648 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1676037725
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1676037725
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1676037725
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1676037725
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1676037725
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1676037725
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1676037725
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1676037725
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1676037725
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1676037725
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1676037725
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1676037725
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1676037725
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_92_245
timestamp 1676037725
transform 1 0 23644 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_92_250
timestamp 1676037725
transform 1 0 24104 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_92_253
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_256
timestamp 1676037725
transform 1 0 24656 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_264
timestamp 1676037725
transform 1 0 25392 0 1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1676037725
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1676037725
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_39
timestamp 1676037725
transform 1 0 4692 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_43
timestamp 1676037725
transform 1 0 5060 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_47
timestamp 1676037725
transform 1 0 5428 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1676037725
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1676037725
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1676037725
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1676037725
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1676037725
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1676037725
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1676037725
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1676037725
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1676037725
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1676037725
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1676037725
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1676037725
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1676037725
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1676037725
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1676037725
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1676037725
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1676037725
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_237
timestamp 1676037725
transform 1 0 22908 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_243
timestamp 1676037725
transform 1 0 23460 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_248
timestamp 1676037725
transform 1 0 23920 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_256
timestamp 1676037725
transform 1 0 24656 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_264
timestamp 1676037725
transform 1 0 25392 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_21
timestamp 1676037725
transform 1 0 3036 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1676037725
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_29
timestamp 1676037725
transform 1 0 3772 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_47
timestamp 1676037725
transform 1 0 5428 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_59
timestamp 1676037725
transform 1 0 6532 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_76
timestamp 1676037725
transform 1 0 8096 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_97
timestamp 1676037725
transform 1 0 10028 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1676037725
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1676037725
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1676037725
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1676037725
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1676037725
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1676037725
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1676037725
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1676037725
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1676037725
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1676037725
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_233
timestamp 1676037725
transform 1 0 22540 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_236
timestamp 1676037725
transform 1 0 22816 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_242
timestamp 1676037725
transform 1 0 23368 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_250
timestamp 1676037725
transform 1 0 24104 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_94_255
timestamp 1676037725
transform 1 0 24564 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_258
timestamp 1676037725
transform 1 0 24840 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_264
timestamp 1676037725
transform 1 0 25392 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1676037725
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1676037725
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_29
timestamp 1676037725
transform 1 0 3772 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_37
timestamp 1676037725
transform 1 0 4508 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1676037725
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_65
timestamp 1676037725
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_82
timestamp 1676037725
transform 1 0 8648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_85
timestamp 1676037725
transform 1 0 8924 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_89
timestamp 1676037725
transform 1 0 9292 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_95_106
timestamp 1676037725
transform 1 0 10856 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_119
timestamp 1676037725
transform 1 0 12052 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_136
timestamp 1676037725
transform 1 0 13616 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_141
timestamp 1676037725
transform 1 0 14076 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_146
timestamp 1676037725
transform 1 0 14536 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_153
timestamp 1676037725
transform 1 0 15180 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_157
timestamp 1676037725
transform 1 0 15548 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_165
timestamp 1676037725
transform 1 0 16284 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_174
timestamp 1676037725
transform 1 0 17112 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_178
timestamp 1676037725
transform 1 0 17480 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_183
timestamp 1676037725
transform 1 0 17940 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_187
timestamp 1676037725
transform 1 0 18308 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_193
timestamp 1676037725
transform 1 0 18860 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_197
timestamp 1676037725
transform 1 0 19228 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_209
timestamp 1676037725
transform 1 0 20332 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_217
timestamp 1676037725
transform 1 0 21068 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_221
timestamp 1676037725
transform 1 0 21436 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_231
timestamp 1676037725
transform 1 0 22356 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_235
timestamp 1676037725
transform 1 0 22724 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_239
timestamp 1676037725
transform 1 0 23092 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_244
timestamp 1676037725
transform 1 0 23552 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_253
timestamp 1676037725
transform 1 0 24380 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_264
timestamp 1676037725
transform 1 0 25392 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24564 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  hold2
timestamp 1676037725
transform 1 0 22448 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1676037725
transform 1 0 24564 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1676037725
transform 1 0 3956 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1676037725
transform 1 0 24656 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1676037725
transform 1 0 23368 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 25116 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 1564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 23276 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1676037725
transform 1 0 25116 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 25116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 25116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1676037725
transform 1 0 25024 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1676037725
transform 1 0 25024 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 25116 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 25116 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1676037725
transform 1 0 25116 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 25116 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1676037725
transform 1 0 25024 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1676037725
transform 1 0 25116 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1676037725
transform 1 0 25024 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1676037725
transform 1 0 25024 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1676037725
transform 1 0 25024 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1676037725
transform 1 0 25116 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1676037725
transform 1 0 25116 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1676037725
transform 1 0 25116 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1676037725
transform 1 0 25116 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1676037725
transform 1 0 25024 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1676037725
transform 1 0 25024 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1676037725
transform 1 0 24472 0 -1 50048
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1676037725
transform 1 0 23828 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1676037725
transform 1 0 23828 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 23184 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 25116 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 25116 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1676037725
transform 1 0 25116 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1676037725
transform 1 0 25116 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1676037725
transform 1 0 5152 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1676037725
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 6348 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1676037725
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1676037725
transform 1 0 7176 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1676037725
transform 1 0 7820 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1676037725
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1676037725
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1676037725
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1676037725
transform 1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1676037725
transform 1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1676037725
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1676037725
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1676037725
transform 1 0 11684 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1676037725
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1676037725
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1676037725
transform 1 0 11040 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1676037725
transform 1 0 2116 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1676037725
transform 1 0 3404 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1676037725
transform 1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1676037725
transform 1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input61
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1676037725
transform 1 0 5152 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 14260 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1676037725
transform 1 0 14904 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1676037725
transform 1 0 16836 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 17664 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1676037725
transform 1 0 19412 0 -1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1676037725
transform 1 0 10396 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input69 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24840 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1676037725
transform 1 0 24840 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input71
timestamp 1676037725
transform 1 0 24840 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input72 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25024 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1676037725
transform 1 0 25024 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1676037725
transform 1 0 23736 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1676037725
transform 1 0 24288 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1676037725
transform 1 0 23000 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1676037725
transform 1 0 20700 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1676037725
transform 1 0 21988 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input79
timestamp 1676037725
transform 1 0 23184 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input80
timestamp 1676037725
transform 1 0 23552 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output81 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17480 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1676037725
transform 1 0 1564 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1676037725
transform 1 0 14904 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1676037725
transform 1 0 23920 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1676037725
transform 1 0 22632 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1676037725
transform 1 0 22080 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1676037725
transform 1 0 22632 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1676037725
transform 1 0 23920 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1676037725
transform 1 0 22632 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1676037725
transform 1 0 22632 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1676037725
transform 1 0 22080 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1676037725
transform 1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1676037725
transform 1 0 22632 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1676037725
transform 1 0 9752 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1676037725
transform 1 0 22632 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1676037725
transform 1 0 22080 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1676037725
transform 1 0 22632 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1676037725
transform 1 0 23920 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1676037725
transform 1 0 22632 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1676037725
transform 1 0 22080 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1676037725
transform 1 0 22632 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1676037725
transform 1 0 23920 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1676037725
transform 1 0 22632 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1676037725
transform 1 0 23920 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1676037725
transform 1 0 18216 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1676037725
transform 1 0 20056 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1676037725
transform 1 0 18216 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1676037725
transform 1 0 20792 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1676037725
transform 1 0 22632 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1676037725
transform 1 0 22080 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1676037725
transform 1 0 23920 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 22632 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 12328 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 18676 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 19412 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 18676 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 12328 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 21252 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 19412 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 21988 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 21712 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 12328 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 21988 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 21252 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 15272 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 23828 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 20056 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 16928 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 22080 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 20240 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 20056 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 12052 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 12972 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 14260 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 14444 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 16836 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 16100 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 16836 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 2024 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 3956 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 4600 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 6624 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 7176 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 9384 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 10764 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 12144 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 25852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 25852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 25852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 25852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 25852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 25852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 25852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 25852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 25852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 25852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 25852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 25852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 25852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 25852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 25852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 25852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 25852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 25852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 25852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 25852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 25852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 25852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 25852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 25852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 25852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 25852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 25852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 25852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 25852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 25852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 25852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 25852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 25852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 25852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 25852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 25852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 25852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 25852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 25852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 25852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 25852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 25852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 25852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 25852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 25852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 25852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 25852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 25852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 25852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 25852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 25852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 25852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 25852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 25852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 25852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 25852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 25852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 25852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 25852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 25852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 25852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 25852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 25852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 25852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 25852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 25852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 25852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 25852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 25852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 25852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 25852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 25852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 25852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 25852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 25852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 25852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 25852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 25852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 25852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 25852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 25852 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 25852 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 25852 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 25852 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 25852 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 25852 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 25852 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 25852 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 25852 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18584 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19872 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22080 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23368 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23552 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23276 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21528 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_9.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21896 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23184 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23552 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23552 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23184 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22080 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_15.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19872 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_17.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17940 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_19.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17020 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16744 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16744 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17388 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_31.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20700 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_33.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22448 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23276 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_35.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23460 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21620 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_47.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19504 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19412 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_49.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19044 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20608 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_bottom_track_51.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23460 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20332 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13340 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9108 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10488 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9292 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11132 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11776 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 11408 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13340 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13064 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12972 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10856 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 9108 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9384 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 8096 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6532 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6624 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10672 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12328 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13064 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12696 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12512 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11776 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10396 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9108 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9016 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10764 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13800 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16100 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16836 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16376 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14904 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 13156 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13892 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15088 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15916 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19596 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20516 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20424 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20240 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21988 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22816 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23092 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 23092 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22632 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22080 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19504 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18768 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 18492 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17296 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__8_.mem_right_track_58.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16836 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_1__198
timestamp 1676037725
transform 1 0 20700 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19504 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20056 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18584 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_3.mux_l2_in_0__153
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21988 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_5.mux_l2_in_0__160
timestamp 1676037725
transform 1 0 21252 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22172 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19228 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_7.mux_l1_in_1__162
timestamp 1676037725
transform 1 0 19688 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19504 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17848 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_9.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22632 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_9.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_9.mux_l2_in_0__163
timestamp 1676037725
transform 1 0 21988 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20240 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_11.mux_l2_in_0__199
timestamp 1676037725
transform 1 0 20884 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22080 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_13.mux_l2_in_0__200
timestamp 1676037725
transform 1 0 24564 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19596 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_15.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_15.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20424 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_15.mux_l2_in_0__201
timestamp 1676037725
transform 1 0 20700 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18492 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_17.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_17.mux_l2_in_0__202
timestamp 1676037725
transform 1 0 18676 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_17.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17848 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_19.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20148 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_19.mux_l2_in_0__151
timestamp 1676037725
transform 1 0 18216 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_19.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20056 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17480 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_29.mux_l2_in_0__152
timestamp 1676037725
transform 1 0 18032 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15916 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_31.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21620 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_31.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_31.mux_l2_in_0__154
timestamp 1676037725
transform 1 0 19688 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_33.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23000 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_33.mux_l2_in_0__155
timestamp 1676037725
transform 1 0 24564 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_33.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22356 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21068 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_35.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_35.mux_l2_in_0__156
timestamp 1676037725
transform 1 0 24748 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_35.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22724 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_45.mux_l2_in_0__157
timestamp 1676037725
transform 1 0 21252 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19688 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_47.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_47.mux_l2_in_0__158
timestamp 1676037725
transform 1 0 20056 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_47.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19872 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19044 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_49.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_49.mux_l2_in_0__159
timestamp 1676037725
transform 1 0 19412 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_49.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18768 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15548 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_51.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23552 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_bottom_track_51.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22264 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_bottom_track_51.mux_l2_in_0__161
timestamp 1676037725
transform 1 0 21252 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12144 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_0.mux_l2_in_1__164
timestamp 1676037725
transform 1 0 7176 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 7636 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16928 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14812 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15180 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9200 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_2.mux_l2_in_1__170
timestamp 1676037725
transform 1 0 9936 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 12144 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15180 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15456 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 10672 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_4.mux_l2_in_1__181
timestamp 1676037725
transform 1 0 11684 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 13524 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17572 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 16836 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15272 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11316 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_6.mux_l2_in_1__192
timestamp 1676037725
transform 1 0 11684 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 14444 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18032 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15640 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13248 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_8.mux_l2_in_1__193
timestamp 1676037725
transform 1 0 9108 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9016 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 11960 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11224 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6624 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_10.mux_l2_in_1__165
timestamp 1676037725
transform 1 0 7360 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9936 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14996 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 7820 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_12.mux_l1_in_1__166
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11500 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16468 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15732 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_14.mux_l1_in_1__167
timestamp 1676037725
transform 1 0 14260 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14812 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_16.mux_l1_in_1__168
timestamp 1676037725
transform 1 0 13432 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12788 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14996 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18952 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14536 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14536 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_18.mux_l2_in_0__169
timestamp 1676037725
transform 1 0 15732 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11408 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_20.mux_l2_in_0__171
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12328 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18032 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_22.mux_l2_in_0__172
timestamp 1676037725
transform 1 0 12328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12236 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_24.mux_l2_in_0__173
timestamp 1676037725
transform 1 0 16100 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18216 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 13800 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_26.mux_l2_in_0__174
timestamp 1676037725
transform 1 0 17664 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16468 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20148 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_28.mux_l1_in_1__175
timestamp 1676037725
transform 1 0 14260 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20608 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_30.mux_l1_in_1__176
timestamp 1676037725
transform 1 0 15456 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15732 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17480 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17848 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_32.mux_l1_in_1__177
timestamp 1676037725
transform 1 0 15732 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21620 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_34.mux_l1_in_1__178
timestamp 1676037725
transform 1 0 13156 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21528 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 13340 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_36.mux_l2_in_0__179
timestamp 1676037725
transform 1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_38.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14720 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_38.mux_l2_in_0__180
timestamp 1676037725
transform 1 0 19412 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_38.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_40.mux_l2_in_0__182
timestamp 1676037725
transform 1 0 16100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24196 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_42.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_42.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_42.mux_l2_in_0__183
timestamp 1676037725
transform 1 0 21988 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_44.mux_l1_in_1__184
timestamp 1676037725
transform 1 0 16652 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18032 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19596 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19688 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l1_in_1_
timestamp 1676037725
transform 1 0 18768 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_46.mux_l1_in_1__185
timestamp 1676037725
transform 1 0 18676 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20424 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_48.mux_l1_in_1__186
timestamp 1676037725
transform 1 0 20700 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l1_in_1_
timestamp 1676037725
transform 1 0 19596 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21436 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 23828 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22816 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_50.mux_l2_in_0__187
timestamp 1676037725
transform 1 0 24656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10948 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19504 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_52.mux_l2_in_0__188
timestamp 1676037725
transform 1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_54.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_54.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20516 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_54.mux_l2_in_0__189
timestamp 1676037725
transform 1 0 21252 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21252 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_56.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17940 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_56.mux_l2_in_0_
timestamp 1676037725
transform 1 0 17296 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_56.mux_l2_in_0__190
timestamp 1676037725
transform 1 0 23184 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__8_.mux_right_track_58.mux_l1_in_1__191
timestamp 1676037725
transform 1 0 11684 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l1_in_1_
timestamp 1676037725
transform 1 0 11040 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__8_.mux_right_track_58.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 25870 56200 25926 57000 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 26200 688 27000 808 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1030 56200 1086 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 26200 25984 27000 26104 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 26200 34144 27000 34264 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 26200 34960 27000 35080 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 26200 35776 27000 35896 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 26200 36592 27000 36712 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 26200 37408 27000 37528 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 26200 38224 27000 38344 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 26200 39040 27000 39160 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 26200 39856 27000 39976 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 26200 40672 27000 40792 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 26200 41488 27000 41608 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 26200 26800 27000 26920 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 26200 42304 27000 42424 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 26200 43120 27000 43240 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 26200 43936 27000 44056 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 26200 44752 27000 44872 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 26200 45568 27000 45688 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 26200 46384 27000 46504 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 26200 47200 27000 47320 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 26200 48016 27000 48136 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 26200 48832 27000 48952 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 26200 49648 27000 49768 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 26200 27616 27000 27736 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 26200 28432 27000 28552 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 26200 29248 27000 29368 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 26200 30064 27000 30184 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 26200 30880 27000 31000 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 26200 31696 27000 31816 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 26200 32512 27000 32632 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 26200 33328 27000 33448 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 26200 1504 27000 1624 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 26200 9664 27000 9784 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 26200 10480 27000 10600 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 26200 11296 27000 11416 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 26200 12112 27000 12232 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 26200 12928 27000 13048 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 26200 13744 27000 13864 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 26200 14560 27000 14680 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 26200 15376 27000 15496 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 26200 16192 27000 16312 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 26200 17008 27000 17128 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 26200 2320 27000 2440 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 26200 17824 27000 17944 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 26200 18640 27000 18760 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 26200 19456 27000 19576 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 26200 20272 27000 20392 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 26200 21088 27000 21208 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 26200 21904 27000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 26200 22720 27000 22840 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 26200 23536 27000 23656 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 26200 24352 27000 24472 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 26200 25168 27000 25288 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 26200 3136 27000 3256 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 26200 3952 27000 4072 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 26200 4768 27000 4888 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 26200 5584 27000 5704 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 26200 6400 27000 6520 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 26200 7216 27000 7336 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 26200 8032 27000 8152 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 26200 8848 27000 8968 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 1858 0 1914 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[0]
port 66 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[10]
port 67 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[11]
port 68 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[12]
port 69 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[13]
port 70 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[14]
port 71 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[15]
port 72 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[16]
port 73 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[17]
port 74 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[18]
port 75 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[19]
port 76 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[1]
port 77 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[20]
port 78 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[21]
port 79 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[22]
port 80 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[23]
port 81 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[24]
port 82 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[25]
port 83 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[26]
port 84 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[27]
port 85 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[28]
port 86 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[29]
port 87 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[2]
port 88 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[3]
port 89 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[4]
port 90 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[5]
port 91 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[6]
port 92 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[7]
port 93 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[8]
port 94 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in_0[9]
port 95 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[0]
port 96 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[10]
port 97 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[11]
port 98 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[12]
port 99 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[13]
port 100 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[14]
port 101 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[15]
port 102 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[16]
port 103 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[17]
port 104 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[18]
port 105 nsew signal tristate
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[19]
port 106 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[1]
port 107 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[20]
port 108 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[21]
port 109 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[22]
port 110 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[23]
port 111 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[24]
port 112 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[25]
port 113 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[26]
port 114 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[27]
port 115 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[28]
port 116 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[29]
port 117 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[2]
port 118 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[3]
port 119 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[4]
port 120 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[5]
port 121 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[6]
port 122 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[7]
port 123 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[8]
port 124 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_out_0[9]
port 125 nsew signal tristate
flabel metal2 s 2410 56200 2466 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 126 nsew signal tristate
flabel metal2 s 3790 56200 3846 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 127 nsew signal tristate
flabel metal2 s 5170 56200 5226 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 128 nsew signal tristate
flabel metal2 s 6550 56200 6606 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 129 nsew signal tristate
flabel metal2 s 13450 56200 13506 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 130 nsew signal input
flabel metal2 s 14830 56200 14886 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 131 nsew signal input
flabel metal2 s 16210 56200 16266 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 132 nsew signal input
flabel metal2 s 17590 56200 17646 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 133 nsew signal input
flabel metal2 s 7930 56200 7986 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 134 nsew signal tristate
flabel metal2 s 9310 56200 9366 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 135 nsew signal tristate
flabel metal2 s 10690 56200 10746 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 136 nsew signal tristate
flabel metal2 s 12070 56200 12126 57000 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 137 nsew signal tristate
flabel metal2 s 18970 56200 19026 57000 0 FreeSans 224 90 0 0 isol_n
port 138 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 prog_clk
port 139 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 prog_reset
port 140 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 reset
port 141 nsew signal input
flabel metal3 s 26200 50464 27000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 142 nsew signal input
flabel metal3 s 26200 51280 27000 51400 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 143 nsew signal input
flabel metal3 s 26200 52096 27000 52216 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 144 nsew signal input
flabel metal3 s 26200 52912 27000 53032 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 145 nsew signal input
flabel metal3 s 26200 53728 27000 53848 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 146 nsew signal input
flabel metal3 s 26200 54544 27000 54664 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 147 nsew signal input
flabel metal3 s 26200 55360 27000 55480 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 148 nsew signal input
flabel metal3 s 26200 56176 27000 56296 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 149 nsew signal input
flabel metal2 s 20350 56200 20406 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
port 150 nsew signal input
flabel metal2 s 21730 56200 21786 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
port 151 nsew signal input
flabel metal2 s 23110 56200 23166 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
port 152 nsew signal input
flabel metal2 s 24490 56200 24546 57000 0 FreeSans 224 90 0 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
port 153 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 154 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 155 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 156 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 157 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 test_enable
port 158 nsew signal input
rlabel metal1 13478 54400 13478 54400 0 VGND
rlabel metal1 13478 53856 13478 53856 0 VPWR
rlabel metal1 10074 29138 10074 29138 0 cby_0__8_.cby_0__1_.ccff_tail
rlabel metal1 9706 30906 9706 30906 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 9292 42670 9292 42670 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal1 9016 44302 9016 44302 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 8280 37978 8280 37978 0 cby_0__8_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 8832 16218 8832 16218 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal1 7498 10438 7498 10438 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal1 11546 12274 11546 12274 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal1 9660 15538 9660 15538 0 cby_0__8_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal1 8050 14586 8050 14586 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal1 9384 10098 9384 10098 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal1 10442 11628 10442 11628 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal1 9200 11866 9200 11866 0 cby_0__8_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal1 8510 21318 8510 21318 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal1 16376 10574 16376 10574 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal1 14306 23018 14306 23018 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal1 10994 20332 10994 20332 0 cby_0__8_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal1 9890 20366 9890 20366 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel metal1 12742 15980 12742 15980 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal1 9752 23834 9752 23834 0 cby_0__8_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal1 13570 9146 13570 9146 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9108 15674 9108 15674 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9062 30702 9062 30702 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 12374 9724 12374 9724 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14352 10234 14352 10234 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12121 12206 12121 12206 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 12650 13294 12650 13294 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 11132 14858 11132 14858 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 10994 15062 10994 15062 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9154 12954 9154 12954 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 10258 12954 10258 12954 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 10166 17238 10166 17238 0 cby_0__8_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 15870 8500 15870 8500 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9062 13498 9062 13498 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 7774 17850 7774 17850 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 15272 8874 15272 8874 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14444 9350 14444 9350 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15272 13158 15272 13158 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 14214 11849 14214 11849 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13202 9078 13202 9078 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 10626 11696 10626 11696 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9798 11866 9798 11866 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 12466 10234 12466 10234 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 8924 12410 8924 12410 0 cby_0__8_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 15824 8806 15824 8806 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9982 23018 9982 23018 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9292 33966 9292 33966 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13432 12614 13432 12614 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13294 14314 13294 14314 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12788 14246 12788 14246 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 11638 16456 11638 16456 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12834 12614 12834 12614 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 12558 14586 12558 14586 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 10258 18394 10258 18394 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 12650 21063 12650 21063 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 11776 18938 11776 18938 0 cby_0__8_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 13662 15878 13662 15878 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 10442 26554 10442 26554 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 9200 29274 9200 29274 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 13340 15334 13340 15334 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13386 14433 13386 14433 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12604 12410 12604 12410 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 10902 18360 10902 18360 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 12144 15946 12144 15946 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 11408 15674 11408 15674 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10488 23630 10488 23630 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 14214 24888 14214 24888 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10350 21658 10350 21658 0 cby_0__8_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 9752 42126 9752 42126 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 11040 44166 11040 44166 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 11224 49130 11224 49130 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 15502 44778 15502 44778 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 9568 44778 9568 44778 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 10212 42670 10212 42670 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 10396 49130 10396 49130 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal2 15042 46172 15042 46172 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 10212 45050 10212 45050 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 9200 44370 9200 44370 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal1 9568 50218 9568 50218 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal1 13938 46614 13938 46614 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 7912 50422 7912 50422 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal2 8510 48756 8510 48756 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 12788 45526 12788 45526 0 cby_0__8_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 25300 54162 25300 54162 0 ccff_head
rlabel metal1 1564 4114 1564 4114 0 ccff_head_0
rlabel metal3 25860 748 25860 748 0 ccff_tail
rlabel metal1 1564 53618 1564 53618 0 ccff_tail_0
rlabel metal1 24702 25398 24702 25398 0 chanx_right_in[0]
rlabel metal2 25346 34391 25346 34391 0 chanx_right_in[10]
rlabel via2 25346 35037 25346 35037 0 chanx_right_in[11]
rlabel metal1 25116 36142 25116 36142 0 chanx_right_in[12]
rlabel metal2 25530 36873 25530 36873 0 chanx_right_in[13]
rlabel metal2 25162 37655 25162 37655 0 chanx_right_in[14]
rlabel via2 25346 38301 25346 38301 0 chanx_right_in[15]
rlabel metal2 25346 39253 25346 39253 0 chanx_right_in[16]
rlabel metal2 25530 40137 25530 40137 0 chanx_right_in[17]
rlabel metal2 25346 40919 25346 40919 0 chanx_right_in[18]
rlabel via2 25162 41565 25162 41565 0 chanx_right_in[19]
rlabel metal2 25346 24820 25346 24820 0 chanx_right_in[1]
rlabel metal2 25162 42483 25162 42483 0 chanx_right_in[20]
rlabel metal2 25530 43401 25530 43401 0 chanx_right_in[21]
rlabel metal2 24794 44183 24794 44183 0 chanx_right_in[22]
rlabel via2 25346 44829 25346 44829 0 chanx_right_in[23]
rlabel metal2 25346 45781 25346 45781 0 chanx_right_in[24]
rlabel metal2 25346 46495 25346 46495 0 chanx_right_in[25]
rlabel metal2 25346 47447 25346 47447 0 chanx_right_in[26]
rlabel via2 25162 48093 25162 48093 0 chanx_right_in[27]
rlabel metal2 25162 49011 25162 49011 0 chanx_right_in[28]
rlabel metal2 25530 49929 25530 49929 0 chanx_right_in[29]
rlabel metal1 24334 25466 24334 25466 0 chanx_right_in[2]
rlabel metal2 24518 28985 24518 28985 0 chanx_right_in[3]
rlabel metal1 23414 29580 23414 29580 0 chanx_right_in[4]
rlabel metal2 25346 29869 25346 29869 0 chanx_right_in[5]
rlabel via2 25530 30923 25530 30923 0 chanx_right_in[6]
rlabel via2 25346 31773 25346 31773 0 chanx_right_in[7]
rlabel metal1 24840 33286 24840 33286 0 chanx_right_in[8]
rlabel metal2 25346 33677 25346 33677 0 chanx_right_in[9]
rlabel metal1 18538 2516 18538 2516 0 chanx_right_out[0]
rlabel metal2 24794 9061 24794 9061 0 chanx_right_out[10]
rlabel metal3 24848 10540 24848 10540 0 chanx_right_out[11]
rlabel metal1 24104 11798 24104 11798 0 chanx_right_out[12]
rlabel metal3 25676 12172 25676 12172 0 chanx_right_out[13]
rlabel metal3 25584 12988 25584 12988 0 chanx_right_out[14]
rlabel metal2 23782 13583 23782 13583 0 chanx_right_out[15]
rlabel metal1 24380 14450 24380 14450 0 chanx_right_out[16]
rlabel metal2 23322 15249 23322 15249 0 chanx_right_out[17]
rlabel metal2 25162 15657 25162 15657 0 chanx_right_out[18]
rlabel metal1 23506 16558 23506 16558 0 chanx_right_out[19]
rlabel metal2 21206 2329 21206 2329 0 chanx_right_out[1]
rlabel metal1 24380 17714 24380 17714 0 chanx_right_out[20]
rlabel metal1 24104 18326 24104 18326 0 chanx_right_out[21]
rlabel metal2 23874 19159 23874 19159 0 chanx_right_out[22]
rlabel metal2 24702 19261 24702 19261 0 chanx_right_out[23]
rlabel metal1 24380 20978 24380 20978 0 chanx_right_out[24]
rlabel metal3 24848 21964 24848 21964 0 chanx_right_out[25]
rlabel metal3 26136 22780 26136 22780 0 chanx_right_out[26]
rlabel metal2 24794 23069 24794 23069 0 chanx_right_out[27]
rlabel metal3 25124 24412 25124 24412 0 chanx_right_out[28]
rlabel metal2 25162 25517 25162 25517 0 chanx_right_out[29]
rlabel metal2 20562 5882 20562 5882 0 chanx_right_out[2]
rlabel metal2 21206 6749 21206 6749 0 chanx_right_out[3]
rlabel metal1 20654 6290 20654 6290 0 chanx_right_out[4]
rlabel metal3 24848 5644 24848 5644 0 chanx_right_out[5]
rlabel metal3 25768 6460 25768 6460 0 chanx_right_out[6]
rlabel metal1 24104 7310 24104 7310 0 chanx_right_out[7]
rlabel metal2 25162 7769 25162 7769 0 chanx_right_out[8]
rlabel metal3 25676 8908 25676 8908 0 chanx_right_out[9]
rlabel metal1 2392 4114 2392 4114 0 chany_bottom_in_0[0]
rlabel metal1 5382 2414 5382 2414 0 chany_bottom_in_0[10]
rlabel metal1 4738 2380 4738 2380 0 chany_bottom_in_0[11]
rlabel metal1 6210 3366 6210 3366 0 chany_bottom_in_0[12]
rlabel metal1 6578 2278 6578 2278 0 chany_bottom_in_0[13]
rlabel metal1 7176 3502 7176 3502 0 chany_bottom_in_0[14]
rlabel metal2 7406 1894 7406 1894 0 chany_bottom_in_0[15]
rlabel metal1 7820 2958 7820 2958 0 chany_bottom_in_0[16]
rlabel metal1 8464 2414 8464 2414 0 chany_bottom_in_0[17]
rlabel metal1 8556 3502 8556 3502 0 chany_bottom_in_0[18]
rlabel metal1 7314 2380 7314 2380 0 chany_bottom_in_0[19]
rlabel metal1 2668 3502 2668 3502 0 chany_bottom_in_0[1]
rlabel metal1 9154 3910 9154 3910 0 chany_bottom_in_0[20]
rlabel metal1 9522 3366 9522 3366 0 chany_bottom_in_0[21]
rlabel metal1 9338 2380 9338 2380 0 chany_bottom_in_0[22]
rlabel metal1 10120 3026 10120 3026 0 chany_bottom_in_0[23]
rlabel metal1 10672 3502 10672 3502 0 chany_bottom_in_0[24]
rlabel metal1 10810 3026 10810 3026 0 chany_bottom_in_0[25]
rlabel metal2 11730 3468 11730 3468 0 chany_bottom_in_0[26]
rlabel metal1 11500 3026 11500 3026 0 chany_bottom_in_0[27]
rlabel metal1 12052 2414 12052 2414 0 chany_bottom_in_0[28]
rlabel metal2 10074 3740 10074 3740 0 chany_bottom_in_0[29]
rlabel metal1 2392 2958 2392 2958 0 chany_bottom_in_0[2]
rlabel metal1 2806 2414 2806 2414 0 chany_bottom_in_0[3]
rlabel metal1 3404 2958 3404 2958 0 chany_bottom_in_0[4]
rlabel metal2 3818 3145 3818 3145 0 chany_bottom_in_0[5]
rlabel metal1 4002 3910 4002 3910 0 chany_bottom_in_0[6]
rlabel metal1 4508 2822 4508 2822 0 chany_bottom_in_0[7]
rlabel metal1 4876 3502 4876 3502 0 chany_bottom_in_0[8]
rlabel metal2 5198 1860 5198 1860 0 chany_bottom_in_0[9]
rlabel metal2 12926 1231 12926 1231 0 chany_bottom_out_0[0]
rlabel metal1 17894 3094 17894 3094 0 chany_bottom_out_0[10]
rlabel metal1 18446 2822 18446 2822 0 chany_bottom_out_0[11]
rlabel metal2 17342 1503 17342 1503 0 chany_bottom_out_0[12]
rlabel metal1 18814 3434 18814 3434 0 chany_bottom_out_0[13]
rlabel metal2 18078 823 18078 823 0 chany_bottom_out_0[14]
rlabel metal2 18446 891 18446 891 0 chany_bottom_out_0[15]
rlabel metal1 20286 3638 20286 3638 0 chany_bottom_out_0[16]
rlabel metal1 19550 3910 19550 3910 0 chany_bottom_out_0[17]
rlabel metal1 22310 2482 22310 2482 0 chany_bottom_out_0[18]
rlabel metal2 19918 1503 19918 1503 0 chany_bottom_out_0[19]
rlabel metal2 13294 1554 13294 1554 0 chany_bottom_out_0[1]
rlabel metal1 20930 3706 20930 3706 0 chany_bottom_out_0[20]
rlabel metal1 20654 5712 20654 5712 0 chany_bottom_out_0[21]
rlabel metal1 16514 6664 16514 6664 0 chany_bottom_out_0[22]
rlabel metal2 21390 1860 21390 1860 0 chany_bottom_out_0[23]
rlabel metal1 21528 6222 21528 6222 0 chany_bottom_out_0[24]
rlabel metal2 22126 1503 22126 1503 0 chany_bottom_out_0[25]
rlabel metal1 22540 8398 22540 8398 0 chany_bottom_out_0[26]
rlabel metal2 21666 5610 21666 5610 0 chany_bottom_out_0[27]
rlabel metal2 23230 1690 23230 1690 0 chany_bottom_out_0[28]
rlabel metal2 17526 3757 17526 3757 0 chany_bottom_out_0[29]
rlabel metal2 13662 1860 13662 1860 0 chany_bottom_out_0[2]
rlabel metal1 14398 3570 14398 3570 0 chany_bottom_out_0[3]
rlabel metal2 14398 1622 14398 1622 0 chany_bottom_out_0[4]
rlabel metal1 15042 2958 15042 2958 0 chany_bottom_out_0[5]
rlabel metal2 17342 2621 17342 2621 0 chany_bottom_out_0[6]
rlabel metal1 16054 3570 16054 3570 0 chany_bottom_out_0[7]
rlabel metal1 16606 2958 16606 2958 0 chany_bottom_out_0[8]
rlabel metal1 16790 4046 16790 4046 0 chany_bottom_out_0[9]
rlabel metal1 21758 32198 21758 32198 0 clknet_0_prog_clk
rlabel metal1 9844 5678 9844 5678 0 clknet_4_0_0_prog_clk
rlabel metal1 6670 48790 6670 48790 0 clknet_4_10_0_prog_clk
rlabel metal2 16790 32062 16790 32062 0 clknet_4_11_0_prog_clk
rlabel metal1 18170 20570 18170 20570 0 clknet_4_12_0_prog_clk
rlabel metal1 23460 24786 23460 24786 0 clknet_4_13_0_prog_clk
rlabel metal1 19090 32266 19090 32266 0 clknet_4_14_0_prog_clk
rlabel metal1 19964 43758 19964 43758 0 clknet_4_15_0_prog_clk
rlabel metal1 11270 6834 11270 6834 0 clknet_4_1_0_prog_clk
rlabel metal2 9798 17442 9798 17442 0 clknet_4_2_0_prog_clk
rlabel metal1 13018 18190 13018 18190 0 clknet_4_3_0_prog_clk
rlabel metal2 16882 13129 16882 13129 0 clknet_4_4_0_prog_clk
rlabel metal2 18538 7106 18538 7106 0 clknet_4_5_0_prog_clk
rlabel metal1 15916 20978 15916 20978 0 clknet_4_6_0_prog_clk
rlabel metal2 20286 18258 20286 18258 0 clknet_4_7_0_prog_clk
rlabel metal2 13386 29648 13386 29648 0 clknet_4_8_0_prog_clk
rlabel metal1 16146 28526 16146 28526 0 clknet_4_9_0_prog_clk
rlabel metal1 2484 54094 2484 54094 0 gfpga_pad_io_soc_dir[0]
rlabel metal1 4140 53618 4140 53618 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 5198 55158 5198 55158 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 6578 54920 6578 54920 0 gfpga_pad_io_soc_dir[3]
rlabel metal2 13662 56236 13662 56236 0 gfpga_pad_io_soc_in[0]
rlabel metal1 14996 54162 14996 54162 0 gfpga_pad_io_soc_in[1]
rlabel metal1 16836 54162 16836 54162 0 gfpga_pad_io_soc_in[2]
rlabel metal1 17756 54162 17756 54162 0 gfpga_pad_io_soc_in[3]
rlabel metal2 7958 55711 7958 55711 0 gfpga_pad_io_soc_out[0]
rlabel metal1 9614 54094 9614 54094 0 gfpga_pad_io_soc_out[1]
rlabel metal1 10718 53652 10718 53652 0 gfpga_pad_io_soc_out[2]
rlabel metal2 12282 56236 12282 56236 0 gfpga_pad_io_soc_out[3]
rlabel metal1 19228 54162 19228 54162 0 isol_n
rlabel metal2 23414 49946 23414 49946 0 net1
rlabel metal1 23552 39270 23552 39270 0 net10
rlabel metal2 22126 22780 22126 22780 0 net100
rlabel metal2 23782 22644 23782 22644 0 net101
rlabel metal2 23966 23052 23966 23052 0 net102
rlabel metal1 22678 25228 22678 25228 0 net103
rlabel metal2 23966 25670 23966 25670 0 net104
rlabel metal2 14950 4862 14950 4862 0 net105
rlabel metal1 18768 3502 18768 3502 0 net106
rlabel metal1 13800 5882 13800 5882 0 net107
rlabel metal1 21620 13294 21620 13294 0 net108
rlabel metal2 10626 4675 10626 4675 0 net109
rlabel metal1 24242 40154 24242 40154 0 net11
rlabel metal2 23552 12614 23552 12614 0 net110
rlabel metal2 12558 6545 12558 6545 0 net111
rlabel metal1 12144 5134 12144 5134 0 net112
rlabel metal2 19642 14178 19642 14178 0 net113
rlabel metal1 18952 3026 18952 3026 0 net114
rlabel metal2 19458 6970 19458 6970 0 net115
rlabel metal1 18078 4590 18078 4590 0 net116
rlabel metal1 19412 3502 19412 3502 0 net117
rlabel metal1 18262 4114 18262 4114 0 net118
rlabel metal1 13432 4590 13432 4590 0 net119
rlabel metal1 25116 40902 25116 40902 0 net12
rlabel metal2 21390 7514 21390 7514 0 net120
rlabel metal1 19918 5678 19918 5678 0 net121
rlabel metal1 23690 2346 23690 2346 0 net122
rlabel metal2 21850 5865 21850 5865 0 net123
rlabel metal2 12650 3825 12650 3825 0 net124
rlabel metal1 21390 3094 21390 3094 0 net125
rlabel metal2 21482 7242 21482 7242 0 net126
rlabel metal2 15502 5882 15502 5882 0 net127
rlabel metal1 23828 5202 23828 5202 0 net128
rlabel metal1 23276 3706 23276 3706 0 net129
rlabel metal1 23368 41514 23368 41514 0 net13
rlabel metal1 17802 5202 17802 5202 0 net130
rlabel metal2 22218 5814 22218 5814 0 net131
rlabel metal1 20792 7854 20792 7854 0 net132
rlabel metal1 20286 8500 20286 8500 0 net133
rlabel metal2 12282 4063 12282 4063 0 net134
rlabel metal1 16882 16966 16882 16966 0 net135
rlabel metal3 17181 15300 17181 15300 0 net136
rlabel metal1 14398 4454 14398 4454 0 net137
rlabel metal1 14490 3026 14490 3026 0 net138
rlabel metal1 16836 2414 16836 2414 0 net139
rlabel metal2 22402 24038 22402 24038 0 net14
rlabel metal1 17020 3502 17020 3502 0 net140
rlabel metal1 18216 13226 18216 13226 0 net141
rlabel metal1 17388 4114 17388 4114 0 net142
rlabel metal1 4646 53210 4646 53210 0 net143
rlabel metal1 5382 52666 5382 52666 0 net144
rlabel metal2 4830 52768 4830 52768 0 net145
rlabel metal1 8556 51510 8556 51510 0 net146
rlabel metal1 7866 51578 7866 51578 0 net147
rlabel metal2 9614 52326 9614 52326 0 net148
rlabel metal2 10718 51442 10718 51442 0 net149
rlabel metal1 24794 42534 24794 42534 0 net15
rlabel metal2 11730 51748 11730 51748 0 net150
rlabel metal1 18262 26010 18262 26010 0 net151
rlabel metal1 17940 27438 17940 27438 0 net152
rlabel metal1 24656 15538 24656 15538 0 net153
rlabel metal2 19734 28288 19734 28288 0 net154
rlabel metal1 22724 26962 22724 26962 0 net155
rlabel metal2 24978 28798 24978 28798 0 net156
rlabel metal1 21850 30226 21850 30226 0 net157
rlabel metal1 20194 30362 20194 30362 0 net158
rlabel metal2 19182 29376 19182 29376 0 net159
rlabel metal1 24748 43078 24748 43078 0 net16
rlabel metal1 21942 19346 21942 19346 0 net160
rlabel metal1 21988 17170 21988 17170 0 net161
rlabel metal1 19688 22746 19688 22746 0 net162
rlabel metal2 22034 21250 22034 21250 0 net163
rlabel metal1 7636 17306 7636 17306 0 net164
rlabel metal1 7222 12274 7222 12274 0 net165
rlabel metal2 8234 12546 8234 12546 0 net166
rlabel metal1 13478 17646 13478 17646 0 net167
rlabel metal2 13202 17374 13202 17374 0 net168
rlabel metal1 15732 16218 15732 16218 0 net169
rlabel metal3 23161 44268 23161 44268 0 net17
rlabel metal2 9982 21250 9982 21250 0 net170
rlabel via2 12742 10795 12742 10795 0 net171
rlabel metal2 12650 7616 12650 7616 0 net172
rlabel metal2 14674 7905 14674 7905 0 net173
rlabel metal1 17296 14314 17296 14314 0 net174
rlabel metal1 14214 15130 14214 15130 0 net175
rlabel metal1 15824 16558 15824 16558 0 net176
rlabel metal1 15870 15130 15870 15130 0 net177
rlabel metal2 13386 8126 13386 8126 0 net178
rlabel metal1 16698 4250 16698 4250 0 net179
rlabel metal1 25208 44710 25208 44710 0 net18
rlabel metal1 18676 5678 18676 5678 0 net180
rlabel metal1 11408 21658 11408 21658 0 net181
rlabel metal1 16100 9894 16100 9894 0 net182
rlabel metal1 21574 9690 21574 9690 0 net183
rlabel metal2 18446 11968 18446 11968 0 net184
rlabel metal1 18768 12274 18768 12274 0 net185
rlabel metal2 20010 11390 20010 11390 0 net186
rlabel metal2 24702 7072 24702 7072 0 net187
rlabel metal1 24380 2482 24380 2482 0 net188
rlabel metal1 21114 3162 21114 3162 0 net189
rlabel metal1 24288 35802 24288 35802 0 net19
rlabel metal2 18906 5661 18906 5661 0 net190
rlabel metal2 11454 8126 11454 8126 0 net191
rlabel metal2 11730 19584 11730 19584 0 net192
rlabel metal2 9430 17408 9430 17408 0 net193
rlabel metal1 10948 12954 10948 12954 0 net194
rlabel metal1 12972 10030 12972 10030 0 net195
rlabel metal1 15410 23086 15410 23086 0 net196
rlabel metal1 15640 25874 15640 25874 0 net197
rlabel metal1 20332 21522 20332 21522 0 net198
rlabel metal1 24978 22066 24978 22066 0 net199
rlabel metal1 4002 4556 4002 4556 0 net2
rlabel metal1 23460 35734 23460 35734 0 net20
rlabel metal1 24380 24242 24380 24242 0 net200
rlabel metal1 20792 23154 20792 23154 0 net201
rlabel metal2 18538 24650 18538 24650 0 net202
rlabel metal2 25254 2040 25254 2040 0 net203
rlabel metal1 25484 25194 25484 25194 0 net204
rlabel metal1 24932 3366 24932 3366 0 net205
rlabel metal1 2024 4250 2024 4250 0 net206
rlabel metal1 5014 4522 5014 4522 0 net207
rlabel metal2 25346 52972 25346 52972 0 net208
rlabel metal1 22356 43826 22356 43826 0 net209
rlabel metal1 25392 29138 25392 29138 0 net21
rlabel metal1 21482 48042 21482 48042 0 net22
rlabel metal2 20010 34204 20010 34204 0 net23
rlabel metal1 22494 41446 22494 41446 0 net24
rlabel metal2 24932 24956 24932 24956 0 net25
rlabel metal1 25070 23188 25070 23188 0 net26
rlabel metal1 22862 29478 22862 29478 0 net27
rlabel metal1 23276 26350 23276 26350 0 net28
rlabel metal1 25070 26384 25070 26384 0 net29
rlabel metal1 22908 25670 22908 25670 0 net3
rlabel metal2 25070 29716 25070 29716 0 net30
rlabel metal1 24656 28458 24656 28458 0 net31
rlabel metal1 24380 28186 24380 28186 0 net32
rlabel metal2 2714 5066 2714 5066 0 net33
rlabel via2 5474 2499 5474 2499 0 net34
rlabel metal2 4554 2176 4554 2176 0 net35
rlabel metal2 6394 4964 6394 4964 0 net36
rlabel metal2 11178 4590 11178 4590 0 net37
rlabel metal1 8004 3638 8004 3638 0 net38
rlabel metal1 8188 3162 8188 3162 0 net39
rlabel metal1 23000 34714 23000 34714 0 net4
rlabel metal2 16238 16320 16238 16320 0 net40
rlabel metal1 8510 2618 8510 2618 0 net41
rlabel metal1 10028 7922 10028 7922 0 net42
rlabel metal2 7130 2074 7130 2074 0 net43
rlabel metal1 3128 3706 3128 3706 0 net44
rlabel metal1 12374 4148 12374 4148 0 net45
rlabel metal1 14168 10574 14168 10574 0 net46
rlabel metal1 9844 2278 9844 2278 0 net47
rlabel metal1 11914 10132 11914 10132 0 net48
rlabel metal1 10488 3706 10488 3706 0 net49
rlabel metal1 25438 34918 25438 34918 0 net5
rlabel metal1 19918 9894 19918 9894 0 net50
rlabel metal1 12006 3060 12006 3060 0 net51
rlabel metal2 20194 9792 20194 9792 0 net52
rlabel metal1 13708 2278 13708 2278 0 net53
rlabel metal1 11362 3468 11362 3468 0 net54
rlabel metal2 2438 5916 2438 5916 0 net55
rlabel metal1 2898 2516 2898 2516 0 net56
rlabel metal2 3726 7446 3726 7446 0 net57
rlabel metal1 5290 3604 5290 3604 0 net58
rlabel metal1 5750 3978 5750 3978 0 net59
rlabel metal1 25530 31246 25530 31246 0 net6
rlabel metal1 6072 3706 6072 3706 0 net60
rlabel metal1 14076 18394 14076 18394 0 net61
rlabel metal1 12926 17102 12926 17102 0 net62
rlabel metal1 13524 53958 13524 53958 0 net63
rlabel metal2 13938 50286 13938 50286 0 net64
rlabel metal2 15594 50014 15594 50014 0 net65
rlabel metal2 15686 49470 15686 49470 0 net66
rlabel metal1 18262 54196 18262 54196 0 net67
rlabel metal1 15226 4692 15226 4692 0 net68
rlabel metal1 21850 50694 21850 50694 0 net69
rlabel metal1 25484 36618 25484 36618 0 net7
rlabel metal1 25990 51306 25990 51306 0 net70
rlabel metal2 16606 31994 16606 31994 0 net71
rlabel metal1 21988 52938 21988 52938 0 net72
rlabel metal1 22218 30090 22218 30090 0 net73
rlabel metal1 17756 32470 17756 32470 0 net74
rlabel metal2 24518 47464 24518 47464 0 net75
rlabel metal1 19872 44166 19872 44166 0 net76
rlabel metal2 16790 32980 16790 32980 0 net77
rlabel metal2 20148 34068 20148 34068 0 net78
rlabel metal1 22770 53958 22770 53958 0 net79
rlabel metal1 25576 37706 25576 37706 0 net8
rlabel metal1 19504 32946 19504 32946 0 net80
rlabel metal1 17848 7854 17848 7854 0 net81
rlabel metal1 1794 53516 1794 53516 0 net82
rlabel metal1 16146 6290 16146 6290 0 net83
rlabel metal1 23966 8534 23966 8534 0 net84
rlabel metal1 24978 7990 24978 7990 0 net85
rlabel metal1 24196 6426 24196 6426 0 net86
rlabel metal1 24334 11322 24334 11322 0 net87
rlabel metal1 24564 11730 24564 11730 0 net88
rlabel metal1 23322 13294 23322 13294 0 net89
rlabel metal1 25300 38182 25300 38182 0 net9
rlabel metal1 24564 13498 24564 13498 0 net90
rlabel metal2 22034 13838 22034 13838 0 net91
rlabel metal1 24380 12410 24380 12410 0 net92
rlabel metal1 22034 13804 22034 13804 0 net93
rlabel metal1 9890 2516 9890 2516 0 net94
rlabel metal1 23736 16422 23736 16422 0 net95
rlabel metal2 22126 18428 22126 18428 0 net96
rlabel metal2 22770 19482 22770 19482 0 net97
rlabel metal2 23506 19278 23506 19278 0 net98
rlabel metal1 22678 20978 22678 20978 0 net99
rlabel metal2 18906 23970 18906 23970 0 prog_clk
rlabel metal2 24610 4522 24610 4522 0 prog_reset
rlabel metal2 24978 50711 24978 50711 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel via2 24978 51323 24978 51323 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal2 24978 52275 24978 52275 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal2 25070 53023 25070 53023 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 25070 53669 25070 53669 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal2 24518 54179 24518 54179 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal3 25584 55420 25584 55420 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel via2 23437 56100 23437 56100 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel metal2 20562 56236 20562 56236 0 right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal1 21896 54162 21896 54162 0 right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal1 23184 54162 23184 54162 0 right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 24518 55711 24518 55711 0 right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal3 2108 1836 2108 1836 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 2062 4148 2062 4148 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 2062 6460 2062 6460 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 1740 8772 1740 8772 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 18768 13838 18768 13838 0 sb_0__8_.mem_bottom_track_1.ccff_head
rlabel metal2 21666 19482 21666 19482 0 sb_0__8_.mem_bottom_track_1.ccff_tail
rlabel metal2 20194 18530 20194 18530 0 sb_0__8_.mem_bottom_track_1.mem_out\[0\]
rlabel metal1 23552 23630 23552 23630 0 sb_0__8_.mem_bottom_track_11.ccff_head
rlabel metal1 25300 24582 25300 24582 0 sb_0__8_.mem_bottom_track_11.ccff_tail
rlabel metal1 25070 23834 25070 23834 0 sb_0__8_.mem_bottom_track_11.mem_out\[0\]
rlabel metal2 22402 27608 22402 27608 0 sb_0__8_.mem_bottom_track_13.ccff_tail
rlabel metal1 25162 27540 25162 27540 0 sb_0__8_.mem_bottom_track_13.mem_out\[0\]
rlabel metal1 20700 26418 20700 26418 0 sb_0__8_.mem_bottom_track_15.ccff_tail
rlabel metal1 23552 28594 23552 28594 0 sb_0__8_.mem_bottom_track_15.mem_out\[0\]
rlabel metal1 19366 26758 19366 26758 0 sb_0__8_.mem_bottom_track_17.ccff_tail
rlabel metal2 22126 27234 22126 27234 0 sb_0__8_.mem_bottom_track_17.mem_out\[0\]
rlabel metal2 18814 30022 18814 30022 0 sb_0__8_.mem_bottom_track_19.ccff_tail
rlabel metal2 18906 29172 18906 29172 0 sb_0__8_.mem_bottom_track_19.mem_out\[0\]
rlabel metal1 18124 31858 18124 31858 0 sb_0__8_.mem_bottom_track_29.ccff_tail
rlabel metal1 17795 31994 17795 31994 0 sb_0__8_.mem_bottom_track_29.mem_out\[0\]
rlabel metal2 25162 19924 25162 19924 0 sb_0__8_.mem_bottom_track_3.ccff_tail
rlabel metal1 23920 20026 23920 20026 0 sb_0__8_.mem_bottom_track_3.mem_out\[0\]
rlabel metal2 21022 29614 21022 29614 0 sb_0__8_.mem_bottom_track_31.ccff_tail
rlabel metal1 20240 31858 20240 31858 0 sb_0__8_.mem_bottom_track_31.mem_out\[0\]
rlabel metal2 23598 28781 23598 28781 0 sb_0__8_.mem_bottom_track_33.ccff_tail
rlabel metal1 22908 31382 22908 31382 0 sb_0__8_.mem_bottom_track_33.mem_out\[0\]
rlabel metal1 25300 32538 25300 32538 0 sb_0__8_.mem_bottom_track_35.ccff_tail
rlabel metal2 25254 31552 25254 31552 0 sb_0__8_.mem_bottom_track_35.mem_out\[0\]
rlabel metal1 23368 33422 23368 33422 0 sb_0__8_.mem_bottom_track_45.ccff_tail
rlabel metal1 22356 33422 22356 33422 0 sb_0__8_.mem_bottom_track_45.mem_out\[0\]
rlabel via1 20562 33422 20562 33422 0 sb_0__8_.mem_bottom_track_47.ccff_tail
rlabel metal1 23322 33830 23322 33830 0 sb_0__8_.mem_bottom_track_47.mem_out\[0\]
rlabel metal1 20884 32198 20884 32198 0 sb_0__8_.mem_bottom_track_49.ccff_tail
rlabel metal2 21206 33082 21206 33082 0 sb_0__8_.mem_bottom_track_49.mem_out\[0\]
rlabel metal2 22126 21522 22126 21522 0 sb_0__8_.mem_bottom_track_5.ccff_tail
rlabel metal1 25300 23154 25300 23154 0 sb_0__8_.mem_bottom_track_5.mem_out\[0\]
rlabel metal1 23966 29070 23966 29070 0 sb_0__8_.mem_bottom_track_51.mem_out\[0\]
rlabel metal1 20838 24378 20838 24378 0 sb_0__8_.mem_bottom_track_7.ccff_tail
rlabel metal1 23046 25806 23046 25806 0 sb_0__8_.mem_bottom_track_7.mem_out\[0\]
rlabel metal1 22264 24106 22264 24106 0 sb_0__8_.mem_bottom_track_9.mem_out\[0\]
rlabel metal1 10994 26418 10994 26418 0 sb_0__8_.mem_right_track_0.ccff_tail
rlabel metal1 19366 43962 19366 43962 0 sb_0__8_.mem_right_track_0.mem_out\[0\]
rlabel metal1 13662 29818 13662 29818 0 sb_0__8_.mem_right_track_0.mem_out\[1\]
rlabel metal2 10902 23766 10902 23766 0 sb_0__8_.mem_right_track_10.ccff_head
rlabel metal1 8740 19142 8740 19142 0 sb_0__8_.mem_right_track_10.ccff_tail
rlabel metal2 11178 23562 11178 23562 0 sb_0__8_.mem_right_track_10.mem_out\[0\]
rlabel metal1 6900 19278 6900 19278 0 sb_0__8_.mem_right_track_10.mem_out\[1\]
rlabel metal2 10902 19244 10902 19244 0 sb_0__8_.mem_right_track_12.ccff_tail
rlabel metal1 8464 18598 8464 18598 0 sb_0__8_.mem_right_track_12.mem_out\[0\]
rlabel metal1 13754 21454 13754 21454 0 sb_0__8_.mem_right_track_14.ccff_tail
rlabel metal1 12926 21046 12926 21046 0 sb_0__8_.mem_right_track_14.mem_out\[0\]
rlabel metal1 14030 20230 14030 20230 0 sb_0__8_.mem_right_track_16.ccff_tail
rlabel metal1 13248 20366 13248 20366 0 sb_0__8_.mem_right_track_16.mem_out\[0\]
rlabel metal2 13570 14960 13570 14960 0 sb_0__8_.mem_right_track_18.ccff_tail
rlabel metal1 15134 16082 15134 16082 0 sb_0__8_.mem_right_track_18.mem_out\[0\]
rlabel metal1 12558 25772 12558 25772 0 sb_0__8_.mem_right_track_2.ccff_tail
rlabel metal1 15778 27948 15778 27948 0 sb_0__8_.mem_right_track_2.mem_out\[0\]
rlabel metal1 9568 21454 9568 21454 0 sb_0__8_.mem_right_track_2.mem_out\[1\]
rlabel metal1 10304 10982 10304 10982 0 sb_0__8_.mem_right_track_20.ccff_tail
rlabel metal1 12144 11186 12144 11186 0 sb_0__8_.mem_right_track_20.mem_out\[0\]
rlabel metal1 10580 5746 10580 5746 0 sb_0__8_.mem_right_track_22.ccff_tail
rlabel metal1 10948 8806 10948 8806 0 sb_0__8_.mem_right_track_22.mem_out\[0\]
rlabel metal1 12466 6970 12466 6970 0 sb_0__8_.mem_right_track_24.ccff_tail
rlabel metal1 11454 5882 11454 5882 0 sb_0__8_.mem_right_track_24.mem_out\[0\]
rlabel metal2 15594 15572 15594 15572 0 sb_0__8_.mem_right_track_26.ccff_tail
rlabel via1 14122 12750 14122 12750 0 sb_0__8_.mem_right_track_26.mem_out\[0\]
rlabel metal1 15916 20026 15916 20026 0 sb_0__8_.mem_right_track_28.ccff_tail
rlabel metal1 15226 19890 15226 19890 0 sb_0__8_.mem_right_track_28.mem_out\[0\]
rlabel metal2 17158 21182 17158 21182 0 sb_0__8_.mem_right_track_30.ccff_tail
rlabel metal1 16744 20774 16744 20774 0 sb_0__8_.mem_right_track_30.mem_out\[0\]
rlabel metal1 18492 18054 18492 18054 0 sb_0__8_.mem_right_track_32.ccff_tail
rlabel metal1 16928 18190 16928 18190 0 sb_0__8_.mem_right_track_32.mem_out\[0\]
rlabel metal2 16698 9282 16698 9282 0 sb_0__8_.mem_right_track_34.ccff_tail
rlabel metal1 17480 15334 17480 15334 0 sb_0__8_.mem_right_track_34.mem_out\[0\]
rlabel metal1 16146 5338 16146 5338 0 sb_0__8_.mem_right_track_36.ccff_tail
rlabel metal1 13800 6222 13800 6222 0 sb_0__8_.mem_right_track_36.mem_out\[0\]
rlabel metal1 16238 5576 16238 5576 0 sb_0__8_.mem_right_track_38.ccff_tail
rlabel metal2 15410 5134 15410 5134 0 sb_0__8_.mem_right_track_38.mem_out\[0\]
rlabel metal1 13662 28594 13662 28594 0 sb_0__8_.mem_right_track_4.ccff_tail
rlabel metal1 15962 29682 15962 29682 0 sb_0__8_.mem_right_track_4.mem_out\[0\]
rlabel metal1 13616 30022 13616 30022 0 sb_0__8_.mem_right_track_4.mem_out\[1\]
rlabel metal1 20562 7310 20562 7310 0 sb_0__8_.mem_right_track_40.ccff_tail
rlabel metal2 17434 7616 17434 7616 0 sb_0__8_.mem_right_track_40.mem_out\[0\]
rlabel metal2 21298 11424 21298 11424 0 sb_0__8_.mem_right_track_42.ccff_tail
rlabel metal1 20792 9962 20792 9962 0 sb_0__8_.mem_right_track_42.mem_out\[0\]
rlabel metal1 20838 15674 20838 15674 0 sb_0__8_.mem_right_track_44.ccff_tail
rlabel metal2 19734 18190 19734 18190 0 sb_0__8_.mem_right_track_44.mem_out\[0\]
rlabel metal2 21390 15810 21390 15810 0 sb_0__8_.mem_right_track_46.ccff_tail
rlabel metal1 22080 16422 22080 16422 0 sb_0__8_.mem_right_track_46.mem_out\[0\]
rlabel metal1 23368 12886 23368 12886 0 sb_0__8_.mem_right_track_48.ccff_tail
rlabel metal1 21712 20366 21712 20366 0 sb_0__8_.mem_right_track_48.mem_out\[0\]
rlabel metal2 23414 10268 23414 10268 0 sb_0__8_.mem_right_track_50.ccff_tail
rlabel metal1 24150 12614 24150 12614 0 sb_0__8_.mem_right_track_50.mem_out\[0\]
rlabel metal2 23874 6970 23874 6970 0 sb_0__8_.mem_right_track_52.ccff_tail
rlabel metal1 20194 10540 20194 10540 0 sb_0__8_.mem_right_track_52.mem_out\[0\]
rlabel metal2 21298 4964 21298 4964 0 sb_0__8_.mem_right_track_54.ccff_tail
rlabel metal2 19826 5304 19826 5304 0 sb_0__8_.mem_right_track_54.mem_out\[0\]
rlabel metal1 17756 7310 17756 7310 0 sb_0__8_.mem_right_track_56.ccff_tail
rlabel metal1 19044 7310 19044 7310 0 sb_0__8_.mem_right_track_56.mem_out\[0\]
rlabel metal1 11868 7922 11868 7922 0 sb_0__8_.mem_right_track_58.mem_out\[0\]
rlabel metal1 13846 24038 13846 24038 0 sb_0__8_.mem_right_track_6.ccff_tail
rlabel metal1 14536 29274 14536 29274 0 sb_0__8_.mem_right_track_6.mem_out\[0\]
rlabel metal1 15870 26860 15870 26860 0 sb_0__8_.mem_right_track_6.mem_out\[1\]
rlabel metal1 14674 24718 14674 24718 0 sb_0__8_.mem_right_track_8.mem_out\[0\]
rlabel metal2 12926 23970 12926 23970 0 sb_0__8_.mem_right_track_8.mem_out\[1\]
rlabel metal1 15640 7786 15640 7786 0 sb_0__8_.mux_bottom_track_1.out
rlabel metal1 20654 19482 20654 19482 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20010 19482 20010 19482 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18998 15062 18998 15062 0 sb_0__8_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21482 14824 21482 14824 0 sb_0__8_.mux_bottom_track_11.out
rlabel metal1 24840 26486 24840 26486 0 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21022 15028 21022 15028 0 sb_0__8_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19964 15334 19964 15334 0 sb_0__8_.mux_bottom_track_13.out
rlabel metal1 22586 24684 22586 24684 0 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22356 22100 22356 22100 0 sb_0__8_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16928 9418 16928 9418 0 sb_0__8_.mux_bottom_track_15.out
rlabel metal1 22471 28662 22471 28662 0 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19412 19380 19412 19380 0 sb_0__8_.mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19504 8806 19504 8806 0 sb_0__8_.mux_bottom_track_17.out
rlabel metal1 18952 24174 18952 24174 0 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18998 20434 18998 20434 0 sb_0__8_.mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20608 3094 20608 3094 0 sb_0__8_.mux_bottom_track_19.out
rlabel metal1 18354 25942 18354 25942 0 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16146 17748 16146 17748 0 sb_0__8_.mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11960 11730 11960 11730 0 sb_0__8_.mux_bottom_track_29.out
rlabel metal1 17802 27302 17802 27302 0 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16836 27574 16836 27574 0 sb_0__8_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20746 7582 20746 7582 0 sb_0__8_.mux_bottom_track_3.out
rlabel metal1 25024 17714 25024 17714 0 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 23736 15980 23736 15980 0 sb_0__8_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 17526 13668 17526 13668 0 sb_0__8_.mux_bottom_track_31.out
rlabel metal2 21666 30022 21666 30022 0 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18768 19822 18768 19822 0 sb_0__8_.mux_bottom_track_31.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 21183 18020 21183 18020 0 sb_0__8_.mux_bottom_track_33.out
rlabel metal1 22816 27098 22816 27098 0 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22632 25738 22632 25738 0 sb_0__8_.mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20930 18598 20930 18598 0 sb_0__8_.mux_bottom_track_35.out
rlabel metal1 24978 28594 24978 28594 0 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 24518 28390 24518 28390 0 sb_0__8_.mux_bottom_track_35.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18814 16694 18814 16694 0 sb_0__8_.mux_bottom_track_45.out
rlabel metal2 22494 32606 22494 32606 0 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20884 20434 20884 20434 0 sb_0__8_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17986 9962 17986 9962 0 sb_0__8_.mux_bottom_track_47.out
rlabel metal2 22034 33601 22034 33601 0 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19550 20434 19550 20434 0 sb_0__8_.mux_bottom_track_47.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15226 21386 15226 21386 0 sb_0__8_.mux_bottom_track_49.out
rlabel metal1 20700 35462 20700 35462 0 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15548 21590 15548 21590 0 sb_0__8_.mux_bottom_track_49.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 20884 10574 20884 10574 0 sb_0__8_.mux_bottom_track_5.out
rlabel metal1 23644 19482 23644 19482 0 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21942 17170 21942 17170 0 sb_0__8_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19734 12614 19734 12614 0 sb_0__8_.mux_bottom_track_51.out
rlabel metal2 24610 23052 24610 23052 0 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20516 12818 20516 12818 0 sb_0__8_.mux_bottom_track_51.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17112 17034 17112 17034 0 sb_0__8_.mux_bottom_track_7.out
rlabel metal1 20838 23086 20838 23086 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19596 23086 19596 23086 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18492 17238 18492 17238 0 sb_0__8_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20102 14246 20102 14246 0 sb_0__8_.mux_bottom_track_9.out
rlabel metal1 22632 26486 22632 26486 0 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21068 14382 21068 14382 0 sb_0__8_.mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21758 25330 21758 25330 0 sb_0__8_.mux_right_track_0.out
rlabel metal1 14122 32742 14122 32742 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14076 31926 14076 31926 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12190 26894 12190 26894 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7636 17034 7636 17034 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 14766 24616 14766 24616 0 sb_0__8_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15088 19142 15088 19142 0 sb_0__8_.mux_right_track_10.out
rlabel metal2 11730 24310 11730 24310 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11638 24786 11638 24786 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10488 18394 10488 18394 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 8556 12682 8556 12682 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 15226 19414 15226 19414 0 sb_0__8_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 22218 20230 22218 20230 0 sb_0__8_.mux_right_track_12.out
rlabel metal1 12098 18734 12098 18734 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7820 12954 7820 12954 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16698 19346 16698 19346 0 sb_0__8_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22494 20910 22494 20910 0 sb_0__8_.mux_right_track_14.out
rlabel metal1 15548 22134 15548 22134 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15226 19856 15226 19856 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14858 21692 14858 21692 0 sb_0__8_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18998 19448 18998 19448 0 sb_0__8_.mux_right_track_16.out
rlabel metal1 15548 20570 15548 20570 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13248 17034 13248 17034 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 19182 19822 19182 19822 0 sb_0__8_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 18722 16320 18722 16320 0 sb_0__8_.mux_right_track_18.out
rlabel metal1 14812 16218 14812 16218 0 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17572 16558 17572 16558 0 sb_0__8_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21022 25296 21022 25296 0 sb_0__8_.mux_right_track_2.out
rlabel metal1 14168 27438 14168 27438 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13616 27370 13616 27370 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12650 26656 12650 26656 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12558 23596 12558 23596 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12834 25772 12834 25772 0 sb_0__8_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 18400 12954 18400 12954 0 sb_0__8_.mux_right_track_20.out
rlabel metal2 12834 10948 12834 10948 0 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12466 12699 12466 12699 0 sb_0__8_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16882 10540 16882 10540 0 sb_0__8_.mux_right_track_22.out
rlabel metal1 10810 6426 10810 6426 0 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12880 7174 12880 7174 0 sb_0__8_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21482 10472 21482 10472 0 sb_0__8_.mux_right_track_24.out
rlabel metal2 13386 6936 13386 6936 0 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14812 8058 14812 8058 0 sb_0__8_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20194 13804 20194 13804 0 sb_0__8_.mux_right_track_26.out
rlabel metal1 14122 12614 14122 12614 0 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20378 13974 20378 13974 0 sb_0__8_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21574 15878 21574 15878 0 sb_0__8_.mux_right_track_28.out
rlabel metal1 17112 23494 17112 23494 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13754 15096 13754 15096 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20102 17646 20102 17646 0 sb_0__8_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23598 17544 23598 17544 0 sb_0__8_.mux_right_track_30.out
rlabel metal1 17940 19890 17940 19890 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15824 16422 15824 16422 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21482 18666 21482 18666 0 sb_0__8_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 22816 15334 22816 15334 0 sb_0__8_.mux_right_track_32.out
rlabel metal1 19412 17714 19412 17714 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16652 14858 16652 14858 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21482 15470 21482 15470 0 sb_0__8_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24472 6290 24472 6290 0 sb_0__8_.mux_right_track_34.out
rlabel metal1 16974 18598 16974 18598 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16928 11730 16928 11730 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21758 11356 21758 11356 0 sb_0__8_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 13570 6681 13570 6681 0 sb_0__8_.mux_right_track_36.out
rlabel metal1 15364 6426 15364 6426 0 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15318 6154 15318 6154 0 sb_0__8_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 24978 2907 24978 2907 0 sb_0__8_.mux_right_track_38.out
rlabel metal1 17940 5746 17940 5746 0 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20562 5712 20562 5712 0 sb_0__8_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22402 23732 22402 23732 0 sb_0__8_.mux_right_track_4.out
rlabel metal1 15640 29274 15640 29274 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15962 29614 15962 29614 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14352 26010 14352 26010 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 10718 23902 10718 23902 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 17802 25500 17802 25500 0 sb_0__8_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 11914 4964 11914 4964 0 sb_0__8_.mux_right_track_40.out
rlabel metal1 20148 7514 20148 7514 0 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22862 7021 22862 7021 0 sb_0__8_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12236 5746 12236 5746 0 sb_0__8_.mux_right_track_42.out
rlabel metal1 20930 10574 20930 10574 0 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19090 10676 19090 10676 0 sb_0__8_.mux_right_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24564 16014 24564 16014 0 sb_0__8_.mux_right_track_44.out
rlabel metal1 19872 15130 19872 15130 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18078 11832 18078 11832 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20746 14892 20746 14892 0 sb_0__8_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20930 9044 20930 9044 0 sb_0__8_.mux_right_track_46.out
rlabel metal1 19734 21896 19734 21896 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 19458 12971 19458 12971 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21114 15878 21114 15878 0 sb_0__8_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21528 13158 21528 13158 0 sb_0__8_.mux_right_track_48.out
rlabel metal1 21298 14450 21298 14450 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19642 11016 19642 11016 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 22770 14586 22770 14586 0 sb_0__8_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11316 5338 11316 5338 0 sb_0__8_.mux_right_track_50.out
rlabel metal1 21344 12614 21344 12614 0 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 20654 9758 20654 9758 0 sb_0__8_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18400 3570 18400 3570 0 sb_0__8_.mux_right_track_52.out
rlabel metal1 21850 10200 21850 10200 0 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22724 2278 22724 2278 0 sb_0__8_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 19964 2550 19964 2550 0 sb_0__8_.mux_right_track_54.out
rlabel metal2 21022 5355 21022 5355 0 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21022 3910 21022 3910 0 sb_0__8_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8096 2278 8096 2278 0 sb_0__8_.mux_right_track_56.out
rlabel metal1 18078 7514 18078 7514 0 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 7866 2176 7866 2176 0 sb_0__8_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24656 5678 24656 5678 0 sb_0__8_.mux_right_track_58.out
rlabel metal1 17388 12954 17388 12954 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11454 8058 11454 8058 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17020 12682 17020 12682 0 sb_0__8_.mux_right_track_58.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 22034 22950 22034 22950 0 sb_0__8_.mux_right_track_6.out
rlabel metal2 15778 28016 15778 28016 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16284 27098 16284 27098 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14950 25296 14950 25296 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14444 23698 14444 23698 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18262 23630 18262 23630 0 sb_0__8_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 16882 22882 16882 22882 0 sb_0__8_.mux_right_track_8.out
rlabel metal2 13754 25534 13754 25534 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13662 25160 13662 25160 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12466 22066 12466 22066 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9154 17306 9154 17306 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 12972 22202 12972 22202 0 sb_0__8_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
<< properties >>
string FIXED_BBOX 0 0 27000 57000
<< end >>
