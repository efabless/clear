VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__0_
  CLASS BLOCK ;
  FOREIGN sb_1__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 115.000 BY 115.000 ;
  PIN SC_IN_TOP
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 111.000 8.650 115.000 ;
    END
  END SC_IN_TOP
  PIN SC_OUT_TOP
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 111.000 106.170 115.000 ;
    END
  END SC_OUT_TOP
  PIN Test_en_N_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 111.000 27.050 115.000 ;
    END
  END Test_en_N_out
  PIN Test_en_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END Test_en_S_in
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 30.710 10.640 32.310 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.700 10.640 58.300 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.690 10.640 84.290 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.680 10.640 110.280 103.600 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 17.715 10.640 19.315 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 43.705 10.640 45.305 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.695 10.640 71.295 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 95.685 10.640 97.285 103.600 ;
    END
  END VPWR
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.680 4.000 84.280 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 26.560 115.000 27.160 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 46.960 115.000 47.560 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 49.000 115.000 49.600 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 51.040 115.000 51.640 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 53.080 115.000 53.680 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 55.120 115.000 55.720 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 57.160 115.000 57.760 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 59.200 115.000 59.800 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 61.240 115.000 61.840 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 63.280 115.000 63.880 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 65.320 115.000 65.920 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 28.600 115.000 29.200 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 30.640 115.000 31.240 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 32.680 115.000 33.280 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 34.720 115.000 35.320 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 36.760 115.000 37.360 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 38.800 115.000 39.400 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 40.840 115.000 41.440 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 42.880 115.000 43.480 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 44.920 115.000 45.520 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 67.360 115.000 67.960 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 87.760 115.000 88.360 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 89.800 115.000 90.400 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 91.840 115.000 92.440 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 93.880 115.000 94.480 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 95.920 115.000 96.520 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 97.960 115.000 98.560 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 100.000 115.000 100.600 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 102.040 115.000 102.640 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 104.080 115.000 104.680 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 106.120 115.000 106.720 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 69.400 115.000 70.000 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 71.440 115.000 72.040 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 73.480 115.000 74.080 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 75.520 115.000 76.120 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 77.560 115.000 78.160 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 79.600 115.000 80.200 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 81.640 115.000 82.240 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 83.680 115.000 84.280 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 85.720 115.000 86.320 ;
    END
  END chanx_right_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 111.000 32.570 115.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 111.000 50.970 115.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 111.000 52.810 115.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 111.000 54.650 115.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 111.000 56.490 115.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 111.000 58.330 115.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 111.000 60.170 115.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 111.000 62.010 115.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 111.000 63.850 115.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 111.000 65.690 115.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 111.000 67.530 115.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 111.000 34.410 115.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 111.000 36.250 115.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 111.000 38.090 115.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 111.000 39.930 115.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 111.000 41.770 115.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 111.000 43.610 115.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 111.000 45.450 115.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 111.000 47.290 115.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 111.000 49.130 115.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 111.000 69.370 115.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 111.000 87.770 115.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 111.000 89.610 115.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 111.000 91.450 115.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 111.000 93.290 115.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 111.000 95.130 115.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 111.000 96.970 115.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 111.000 98.810 115.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 111.000 100.650 115.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 111.000 102.490 115.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 111.000 104.330 115.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 111.000 71.210 115.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 111.000 73.050 115.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 111.000 74.890 115.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 111.000 76.730 115.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 111.000 78.570 115.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 111.000 80.410 115.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 111.000 82.250 115.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 111.000 84.090 115.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 111.000 85.930 115.000 ;
    END
  END chany_top_out[9]
  PIN clk_3_N_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 111.000 28.890 115.000 ;
    END
  END clk_3_N_out
  PIN clk_3_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END clk_3_S_in
  PIN left_bottom_grid_pin_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 18.400 4.000 19.000 ;
    END
  END left_bottom_grid_pin_11_
  PIN left_bottom_grid_pin_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END left_bottom_grid_pin_13_
  PIN left_bottom_grid_pin_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END left_bottom_grid_pin_15_
  PIN left_bottom_grid_pin_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END left_bottom_grid_pin_17_
  PIN left_bottom_grid_pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END left_bottom_grid_pin_1_
  PIN left_bottom_grid_pin_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END left_bottom_grid_pin_3_
  PIN left_bottom_grid_pin_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END left_bottom_grid_pin_5_
  PIN left_bottom_grid_pin_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END left_bottom_grid_pin_7_
  PIN left_bottom_grid_pin_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END left_bottom_grid_pin_9_
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 111.000 25.210 115.000 ;
    END
  END prog_clk_0_N_in
  PIN prog_clk_3_N_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 111.000 30.730 115.000 ;
    END
  END prog_clk_3_N_out
  PIN prog_clk_3_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END prog_clk_3_S_in
  PIN right_bottom_grid_pin_11_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 18.400 115.000 19.000 ;
    END
  END right_bottom_grid_pin_11_
  PIN right_bottom_grid_pin_13_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 20.440 115.000 21.040 ;
    END
  END right_bottom_grid_pin_13_
  PIN right_bottom_grid_pin_15_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 22.480 115.000 23.080 ;
    END
  END right_bottom_grid_pin_15_
  PIN right_bottom_grid_pin_17_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 24.520 115.000 25.120 ;
    END
  END right_bottom_grid_pin_17_
  PIN right_bottom_grid_pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 8.200 115.000 8.800 ;
    END
  END right_bottom_grid_pin_1_
  PIN right_bottom_grid_pin_3_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 10.240 115.000 10.840 ;
    END
  END right_bottom_grid_pin_3_
  PIN right_bottom_grid_pin_5_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 12.280 115.000 12.880 ;
    END
  END right_bottom_grid_pin_5_
  PIN right_bottom_grid_pin_7_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 14.320 115.000 14.920 ;
    END
  END right_bottom_grid_pin_7_
  PIN right_bottom_grid_pin_9_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 16.360 115.000 16.960 ;
    END
  END right_bottom_grid_pin_9_
  PIN top_left_grid_pin_42_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 111.000 10.490 115.000 ;
    END
  END top_left_grid_pin_42_
  PIN top_left_grid_pin_43_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 111.000 12.330 115.000 ;
    END
  END top_left_grid_pin_43_
  PIN top_left_grid_pin_44_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 111.000 14.170 115.000 ;
    END
  END top_left_grid_pin_44_
  PIN top_left_grid_pin_45_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 111.000 16.010 115.000 ;
    END
  END top_left_grid_pin_45_
  PIN top_left_grid_pin_46_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 111.000 17.850 115.000 ;
    END
  END top_left_grid_pin_46_
  PIN top_left_grid_pin_47_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 111.000 19.690 115.000 ;
    END
  END top_left_grid_pin_47_
  PIN top_left_grid_pin_48_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 111.000 21.530 115.000 ;
    END
  END top_left_grid_pin_48_
  PIN top_left_grid_pin_49_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 111.000 23.370 115.000 ;
    END
  END top_left_grid_pin_49_
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 109.480 103.445 ;
      LAYER met1 ;
        RECT 5.520 10.640 112.170 104.340 ;
      LAYER met2 ;
        RECT 6.530 110.720 8.090 111.250 ;
        RECT 8.930 110.720 9.930 111.250 ;
        RECT 10.770 110.720 11.770 111.250 ;
        RECT 12.610 110.720 13.610 111.250 ;
        RECT 14.450 110.720 15.450 111.250 ;
        RECT 16.290 110.720 17.290 111.250 ;
        RECT 18.130 110.720 19.130 111.250 ;
        RECT 19.970 110.720 20.970 111.250 ;
        RECT 21.810 110.720 22.810 111.250 ;
        RECT 23.650 110.720 24.650 111.250 ;
        RECT 25.490 110.720 26.490 111.250 ;
        RECT 27.330 110.720 28.330 111.250 ;
        RECT 29.170 110.720 30.170 111.250 ;
        RECT 31.010 110.720 32.010 111.250 ;
        RECT 32.850 110.720 33.850 111.250 ;
        RECT 34.690 110.720 35.690 111.250 ;
        RECT 36.530 110.720 37.530 111.250 ;
        RECT 38.370 110.720 39.370 111.250 ;
        RECT 40.210 110.720 41.210 111.250 ;
        RECT 42.050 110.720 43.050 111.250 ;
        RECT 43.890 110.720 44.890 111.250 ;
        RECT 45.730 110.720 46.730 111.250 ;
        RECT 47.570 110.720 48.570 111.250 ;
        RECT 49.410 110.720 50.410 111.250 ;
        RECT 51.250 110.720 52.250 111.250 ;
        RECT 53.090 110.720 54.090 111.250 ;
        RECT 54.930 110.720 55.930 111.250 ;
        RECT 56.770 110.720 57.770 111.250 ;
        RECT 58.610 110.720 59.610 111.250 ;
        RECT 60.450 110.720 61.450 111.250 ;
        RECT 62.290 110.720 63.290 111.250 ;
        RECT 64.130 110.720 65.130 111.250 ;
        RECT 65.970 110.720 66.970 111.250 ;
        RECT 67.810 110.720 68.810 111.250 ;
        RECT 69.650 110.720 70.650 111.250 ;
        RECT 71.490 110.720 72.490 111.250 ;
        RECT 73.330 110.720 74.330 111.250 ;
        RECT 75.170 110.720 76.170 111.250 ;
        RECT 77.010 110.720 78.010 111.250 ;
        RECT 78.850 110.720 79.850 111.250 ;
        RECT 80.690 110.720 81.690 111.250 ;
        RECT 82.530 110.720 83.530 111.250 ;
        RECT 84.370 110.720 85.370 111.250 ;
        RECT 86.210 110.720 87.210 111.250 ;
        RECT 88.050 110.720 89.050 111.250 ;
        RECT 89.890 110.720 90.890 111.250 ;
        RECT 91.730 110.720 92.730 111.250 ;
        RECT 93.570 110.720 94.570 111.250 ;
        RECT 95.410 110.720 96.410 111.250 ;
        RECT 97.250 110.720 98.250 111.250 ;
        RECT 99.090 110.720 100.090 111.250 ;
        RECT 100.930 110.720 101.930 111.250 ;
        RECT 102.770 110.720 103.770 111.250 ;
        RECT 104.610 110.720 105.610 111.250 ;
        RECT 106.450 110.720 112.140 111.250 ;
        RECT 6.530 4.280 112.140 110.720 ;
        RECT 6.530 3.670 10.850 4.280 ;
        RECT 11.690 3.670 33.850 4.280 ;
        RECT 34.690 3.670 56.850 4.280 ;
        RECT 57.690 3.670 79.850 4.280 ;
        RECT 80.690 3.670 102.850 4.280 ;
        RECT 103.690 3.670 112.140 4.280 ;
      LAYER met3 ;
        RECT 4.400 105.720 110.600 106.585 ;
        RECT 4.000 105.080 111.010 105.720 ;
        RECT 4.400 103.680 110.600 105.080 ;
        RECT 4.000 103.040 111.010 103.680 ;
        RECT 4.400 101.640 110.600 103.040 ;
        RECT 4.000 101.000 111.010 101.640 ;
        RECT 4.400 99.600 110.600 101.000 ;
        RECT 4.000 98.960 111.010 99.600 ;
        RECT 4.400 97.560 110.600 98.960 ;
        RECT 4.000 96.920 111.010 97.560 ;
        RECT 4.400 95.520 110.600 96.920 ;
        RECT 4.000 94.880 111.010 95.520 ;
        RECT 4.400 93.480 110.600 94.880 ;
        RECT 4.000 92.840 111.010 93.480 ;
        RECT 4.400 91.440 110.600 92.840 ;
        RECT 4.000 90.800 111.010 91.440 ;
        RECT 4.400 89.400 110.600 90.800 ;
        RECT 4.000 88.760 111.010 89.400 ;
        RECT 4.400 87.360 110.600 88.760 ;
        RECT 4.000 86.720 111.010 87.360 ;
        RECT 4.400 85.320 110.600 86.720 ;
        RECT 4.000 84.680 111.010 85.320 ;
        RECT 4.400 83.280 110.600 84.680 ;
        RECT 4.000 82.640 111.010 83.280 ;
        RECT 4.400 81.240 110.600 82.640 ;
        RECT 4.000 80.600 111.010 81.240 ;
        RECT 4.400 79.200 110.600 80.600 ;
        RECT 4.000 78.560 111.010 79.200 ;
        RECT 4.400 77.160 110.600 78.560 ;
        RECT 4.000 76.520 111.010 77.160 ;
        RECT 4.400 75.120 110.600 76.520 ;
        RECT 4.000 74.480 111.010 75.120 ;
        RECT 4.400 73.080 110.600 74.480 ;
        RECT 4.000 72.440 111.010 73.080 ;
        RECT 4.400 71.040 110.600 72.440 ;
        RECT 4.000 70.400 111.010 71.040 ;
        RECT 4.400 69.000 110.600 70.400 ;
        RECT 4.000 68.360 111.010 69.000 ;
        RECT 4.400 66.960 110.600 68.360 ;
        RECT 4.000 66.320 111.010 66.960 ;
        RECT 4.400 64.920 110.600 66.320 ;
        RECT 4.000 64.280 111.010 64.920 ;
        RECT 4.400 62.880 110.600 64.280 ;
        RECT 4.000 62.240 111.010 62.880 ;
        RECT 4.400 60.840 110.600 62.240 ;
        RECT 4.000 60.200 111.010 60.840 ;
        RECT 4.400 58.800 110.600 60.200 ;
        RECT 4.000 58.160 111.010 58.800 ;
        RECT 4.400 56.760 110.600 58.160 ;
        RECT 4.000 56.120 111.010 56.760 ;
        RECT 4.400 54.720 110.600 56.120 ;
        RECT 4.000 54.080 111.010 54.720 ;
        RECT 4.400 52.680 110.600 54.080 ;
        RECT 4.000 52.040 111.010 52.680 ;
        RECT 4.400 50.640 110.600 52.040 ;
        RECT 4.000 50.000 111.010 50.640 ;
        RECT 4.400 48.600 110.600 50.000 ;
        RECT 4.000 47.960 111.010 48.600 ;
        RECT 4.400 46.560 110.600 47.960 ;
        RECT 4.000 45.920 111.010 46.560 ;
        RECT 4.400 44.520 110.600 45.920 ;
        RECT 4.000 43.880 111.010 44.520 ;
        RECT 4.400 42.480 110.600 43.880 ;
        RECT 4.000 41.840 111.010 42.480 ;
        RECT 4.400 40.440 110.600 41.840 ;
        RECT 4.000 39.800 111.010 40.440 ;
        RECT 4.400 38.400 110.600 39.800 ;
        RECT 4.000 37.760 111.010 38.400 ;
        RECT 4.400 36.360 110.600 37.760 ;
        RECT 4.000 35.720 111.010 36.360 ;
        RECT 4.400 34.320 110.600 35.720 ;
        RECT 4.000 33.680 111.010 34.320 ;
        RECT 4.400 32.280 110.600 33.680 ;
        RECT 4.000 31.640 111.010 32.280 ;
        RECT 4.400 30.240 110.600 31.640 ;
        RECT 4.000 29.600 111.010 30.240 ;
        RECT 4.400 28.200 110.600 29.600 ;
        RECT 4.000 27.560 111.010 28.200 ;
        RECT 4.400 26.160 110.600 27.560 ;
        RECT 4.000 25.520 111.010 26.160 ;
        RECT 4.400 24.120 110.600 25.520 ;
        RECT 4.000 23.480 111.010 24.120 ;
        RECT 4.400 22.080 110.600 23.480 ;
        RECT 4.000 21.440 111.010 22.080 ;
        RECT 4.400 20.040 110.600 21.440 ;
        RECT 4.000 19.400 111.010 20.040 ;
        RECT 4.400 18.000 110.600 19.400 ;
        RECT 4.000 17.360 111.010 18.000 ;
        RECT 4.400 15.960 110.600 17.360 ;
        RECT 4.000 15.320 111.010 15.960 ;
        RECT 4.400 13.920 110.600 15.320 ;
        RECT 4.000 13.280 111.010 13.920 ;
        RECT 4.400 11.880 110.600 13.280 ;
        RECT 4.000 11.240 111.010 11.880 ;
        RECT 4.400 9.840 110.600 11.240 ;
        RECT 4.000 9.200 111.010 9.840 ;
        RECT 4.400 8.335 110.600 9.200 ;
      LAYER met4 ;
        RECT 19.715 14.455 30.310 101.145 ;
        RECT 32.710 14.455 43.305 101.145 ;
        RECT 45.705 14.455 56.300 101.145 ;
        RECT 58.700 14.455 69.295 101.145 ;
        RECT 71.695 14.455 82.290 101.145 ;
        RECT 84.690 14.455 95.285 101.145 ;
        RECT 97.685 14.455 102.745 101.145 ;
  END
END sb_1__0_
END LIBRARY

