magic
tech sky130A
magscale 1 2
timestamp 1656943348
<< viali >>
rect 7941 20553 7975 20587
rect 8493 20553 8527 20587
rect 9321 20553 9355 20587
rect 11621 20553 11655 20587
rect 14289 20553 14323 20587
rect 18705 20553 18739 20587
rect 19441 20553 19475 20587
rect 13001 20485 13035 20519
rect 6653 20417 6687 20451
rect 7205 20417 7239 20451
rect 7757 20417 7791 20451
rect 8309 20417 8343 20451
rect 10517 20417 10551 20451
rect 14105 20417 14139 20451
rect 15025 20417 15059 20451
rect 15669 20417 15703 20451
rect 16681 20417 16715 20451
rect 17693 20417 17727 20451
rect 18245 20417 18279 20451
rect 18521 20417 18555 20451
rect 19257 20417 19291 20451
rect 21106 20417 21140 20451
rect 9413 20349 9447 20383
rect 9597 20349 9631 20383
rect 10333 20349 10367 20383
rect 21373 20349 21407 20383
rect 13737 20281 13771 20315
rect 15853 20281 15887 20315
rect 16865 20281 16899 20315
rect 18061 20281 18095 20315
rect 5641 20213 5675 20247
rect 6009 20213 6043 20247
rect 6837 20213 6871 20247
rect 7389 20213 7423 20247
rect 8953 20213 8987 20247
rect 10885 20213 10919 20247
rect 12173 20213 12207 20247
rect 12633 20213 12667 20247
rect 13369 20213 13403 20247
rect 14657 20213 14691 20247
rect 15209 20213 15243 20247
rect 16221 20213 16255 20247
rect 17509 20213 17543 20247
rect 19993 20213 20027 20247
rect 7941 20009 7975 20043
rect 18613 20009 18647 20043
rect 6745 19873 6779 19907
rect 16221 19873 16255 19907
rect 16957 19873 16991 19907
rect 19441 19873 19475 19907
rect 21373 19873 21407 19907
rect 4445 19805 4479 19839
rect 6285 19805 6319 19839
rect 7021 19805 7055 19839
rect 7757 19805 7791 19839
rect 8309 19805 8343 19839
rect 10609 19805 10643 19839
rect 10885 19805 10919 19839
rect 12909 19805 12943 19839
rect 13277 19805 13311 19839
rect 15485 19805 15519 19839
rect 15945 19805 15979 19839
rect 17141 19805 17175 19839
rect 17417 19805 17451 19839
rect 18245 19805 18279 19839
rect 18797 19805 18831 19839
rect 19257 19805 19291 19839
rect 10342 19737 10376 19771
rect 11152 19737 11186 19771
rect 15218 19737 15252 19771
rect 21106 19737 21140 19771
rect 4629 19669 4663 19703
rect 5089 19669 5123 19703
rect 5733 19669 5767 19703
rect 6101 19669 6135 19703
rect 7389 19669 7423 19703
rect 8493 19669 8527 19703
rect 9229 19669 9263 19703
rect 12265 19669 12299 19703
rect 12541 19669 12575 19703
rect 13461 19669 13495 19703
rect 14105 19669 14139 19703
rect 17601 19669 17635 19703
rect 18061 19669 18095 19703
rect 19993 19669 20027 19703
rect 6377 19465 6411 19499
rect 6745 19465 6779 19499
rect 8125 19465 8159 19499
rect 11161 19465 11195 19499
rect 13001 19465 13035 19499
rect 14657 19465 14691 19499
rect 18705 19465 18739 19499
rect 7573 19397 7607 19431
rect 10026 19397 10060 19431
rect 12357 19397 12391 19431
rect 12725 19397 12759 19431
rect 15770 19397 15804 19431
rect 17316 19397 17350 19431
rect 21189 19397 21223 19431
rect 5641 19329 5675 19363
rect 5733 19329 5767 19363
rect 7849 19329 7883 19363
rect 9238 19329 9272 19363
rect 14114 19329 14148 19363
rect 14381 19329 14415 19363
rect 19818 19329 19852 19363
rect 20085 19329 20119 19363
rect 20545 19329 20579 19363
rect 4905 19261 4939 19295
rect 5917 19261 5951 19295
rect 6837 19261 6871 19295
rect 7021 19261 7055 19295
rect 9505 19261 9539 19295
rect 9781 19261 9815 19295
rect 16037 19261 16071 19295
rect 17049 19261 17083 19295
rect 11529 19193 11563 19227
rect 5273 19125 5307 19159
rect 11897 19125 11931 19159
rect 16681 19125 16715 19159
rect 18429 19125 18463 19159
rect 18705 18921 18739 18955
rect 11437 18853 11471 18887
rect 16497 18853 16531 18887
rect 6745 18785 6779 18819
rect 20637 18785 20671 18819
rect 6929 18717 6963 18751
rect 8585 18717 8619 18751
rect 10333 18717 10367 18751
rect 12817 18717 12851 18751
rect 13185 18717 13219 18751
rect 13737 18717 13771 18751
rect 14197 18717 14231 18751
rect 14473 18717 14507 18751
rect 16313 18717 16347 18751
rect 18245 18717 18279 18751
rect 18889 18717 18923 18751
rect 20370 18717 20404 18751
rect 20913 18717 20947 18751
rect 8340 18649 8374 18683
rect 10066 18649 10100 18683
rect 12572 18649 12606 18683
rect 14718 18649 14752 18683
rect 18000 18649 18034 18683
rect 21189 18649 21223 18683
rect 5733 18581 5767 18615
rect 6101 18581 6135 18615
rect 7205 18581 7239 18615
rect 8953 18581 8987 18615
rect 10701 18581 10735 18615
rect 10977 18581 11011 18615
rect 15853 18581 15887 18615
rect 16865 18581 16899 18615
rect 19257 18581 19291 18615
rect 6745 18377 6779 18411
rect 7849 18377 7883 18411
rect 8585 18377 8619 18411
rect 16037 18377 16071 18411
rect 19717 18377 19751 18411
rect 13654 18309 13688 18343
rect 14534 18309 14568 18343
rect 7113 18241 7147 18275
rect 7941 18241 7975 18275
rect 10158 18241 10192 18275
rect 10425 18241 10459 18275
rect 13921 18241 13955 18275
rect 14289 18241 14323 18275
rect 16937 18241 16971 18275
rect 18337 18241 18371 18275
rect 18593 18241 18627 18275
rect 19993 18241 20027 18275
rect 20249 18241 20283 18275
rect 8125 18173 8159 18207
rect 16681 18173 16715 18207
rect 9045 18105 9079 18139
rect 12541 18105 12575 18139
rect 7481 18037 7515 18071
rect 10701 18037 10735 18071
rect 11069 18037 11103 18071
rect 11805 18037 11839 18071
rect 12173 18037 12207 18071
rect 15669 18037 15703 18071
rect 18061 18037 18095 18071
rect 21373 18037 21407 18071
rect 13185 17833 13219 17867
rect 17141 17833 17175 17867
rect 19993 17833 20027 17867
rect 19625 17765 19659 17799
rect 7205 17697 7239 17731
rect 7481 17629 7515 17663
rect 9045 17629 9079 17663
rect 9781 17629 9815 17663
rect 10037 17629 10071 17663
rect 11805 17629 11839 17663
rect 13553 17629 13587 17663
rect 14197 17629 14231 17663
rect 14841 17629 14875 17663
rect 15117 17629 15151 17663
rect 16865 17629 16899 17663
rect 18521 17629 18555 17663
rect 19441 17629 19475 17663
rect 21373 17629 21407 17663
rect 12050 17561 12084 17595
rect 15362 17561 15396 17595
rect 18254 17561 18288 17595
rect 21128 17561 21162 17595
rect 11161 17493 11195 17527
rect 11437 17493 11471 17527
rect 16497 17493 16531 17527
rect 18797 17493 18831 17527
rect 4537 17289 4571 17323
rect 4905 17289 4939 17323
rect 5549 17289 5583 17323
rect 7665 17289 7699 17323
rect 8033 17289 8067 17323
rect 11989 17289 12023 17323
rect 5641 17221 5675 17255
rect 12633 17221 12667 17255
rect 13001 17221 13035 17255
rect 10158 17153 10192 17187
rect 14850 17153 14884 17187
rect 18061 17153 18095 17187
rect 18337 17153 18371 17187
rect 20002 17153 20036 17187
rect 20269 17153 20303 17187
rect 20637 17153 20671 17187
rect 5457 17085 5491 17119
rect 8125 17085 8159 17119
rect 8217 17085 8251 17119
rect 10425 17085 10459 17119
rect 15117 17085 15151 17119
rect 15577 17085 15611 17119
rect 15945 17085 15979 17119
rect 20821 17085 20855 17119
rect 8769 17017 8803 17051
rect 13737 17017 13771 17051
rect 18521 17017 18555 17051
rect 6009 16949 6043 16983
rect 9045 16949 9079 16983
rect 10701 16949 10735 16983
rect 11069 16949 11103 16983
rect 11529 16949 11563 16983
rect 12265 16949 12299 16983
rect 13461 16949 13495 16983
rect 16773 16949 16807 16983
rect 17233 16949 17267 16983
rect 17877 16949 17911 16983
rect 18889 16949 18923 16983
rect 17509 16677 17543 16711
rect 14105 16609 14139 16643
rect 8585 16541 8619 16575
rect 9045 16541 9079 16575
rect 10701 16541 10735 16575
rect 15761 16541 15795 16575
rect 16028 16541 16062 16575
rect 18889 16541 18923 16575
rect 19257 16541 19291 16575
rect 20913 16541 20947 16575
rect 8318 16473 8352 16507
rect 9290 16473 9324 16507
rect 10968 16473 11002 16507
rect 14350 16473 14384 16507
rect 18622 16473 18656 16507
rect 19502 16473 19536 16507
rect 4537 16405 4571 16439
rect 6469 16405 6503 16439
rect 7205 16405 7239 16439
rect 10425 16405 10459 16439
rect 12081 16405 12115 16439
rect 12449 16405 12483 16439
rect 13001 16405 13035 16439
rect 13369 16405 13403 16439
rect 15485 16405 15519 16439
rect 17141 16405 17175 16439
rect 20637 16405 20671 16439
rect 21097 16405 21131 16439
rect 4169 16201 4203 16235
rect 5273 16201 5307 16235
rect 6653 16201 6687 16235
rect 11897 16201 11931 16235
rect 18061 16201 18095 16235
rect 20361 16201 20395 16235
rect 20913 16201 20947 16235
rect 16948 16133 16982 16167
rect 18766 16133 18800 16167
rect 5181 16065 5215 16099
rect 6745 16065 6779 16099
rect 8686 16065 8720 16099
rect 10353 16065 10387 16099
rect 13010 16065 13044 16099
rect 13820 16065 13854 16099
rect 20177 16065 20211 16099
rect 20729 16065 20763 16099
rect 3985 15997 4019 16031
rect 4077 15997 4111 16031
rect 5457 15997 5491 16031
rect 6561 15997 6595 16031
rect 8953 15997 8987 16031
rect 10609 15997 10643 16031
rect 13277 15997 13311 16031
rect 13553 15997 13587 16031
rect 16681 15997 16715 16031
rect 18521 15997 18555 16031
rect 14933 15929 14967 15963
rect 4537 15861 4571 15895
rect 4813 15861 4847 15895
rect 5825 15861 5859 15895
rect 7113 15861 7147 15895
rect 7573 15861 7607 15895
rect 9229 15861 9263 15895
rect 10977 15861 11011 15895
rect 15209 15861 15243 15895
rect 15669 15861 15703 15895
rect 16221 15861 16255 15895
rect 19901 15861 19935 15895
rect 21281 15861 21315 15895
rect 9781 15589 9815 15623
rect 5733 15521 5767 15555
rect 6745 15521 6779 15555
rect 6837 15521 6871 15555
rect 5917 15453 5951 15487
rect 11161 15453 11195 15487
rect 13102 15453 13136 15487
rect 13369 15453 13403 15487
rect 15577 15453 15611 15487
rect 15853 15453 15887 15487
rect 17509 15453 17543 15487
rect 18153 15453 18187 15487
rect 18797 15453 18831 15487
rect 19257 15453 19291 15487
rect 21373 15453 21407 15487
rect 5825 15385 5859 15419
rect 6929 15385 6963 15419
rect 7941 15385 7975 15419
rect 10894 15385 10928 15419
rect 15310 15385 15344 15419
rect 16098 15385 16132 15419
rect 21106 15385 21140 15419
rect 4629 15317 4663 15351
rect 6285 15317 6319 15351
rect 7297 15317 7331 15351
rect 7665 15317 7699 15351
rect 9137 15317 9171 15351
rect 11437 15317 11471 15351
rect 11989 15317 12023 15351
rect 13737 15317 13771 15351
rect 14197 15317 14231 15351
rect 17233 15317 17267 15351
rect 19717 15317 19751 15351
rect 19993 15317 20027 15351
rect 4629 15113 4663 15147
rect 6837 15113 6871 15147
rect 14933 15113 14967 15147
rect 5733 15045 5767 15079
rect 7297 15045 7331 15079
rect 4537 14977 4571 15011
rect 5641 14977 5675 15011
rect 6377 14977 6411 15011
rect 7205 14977 7239 15011
rect 10037 14977 10071 15011
rect 16046 14977 16080 15011
rect 16313 14977 16347 15011
rect 19973 14977 20007 15011
rect 4445 14909 4479 14943
rect 5917 14909 5951 14943
rect 7481 14909 7515 14943
rect 9781 14909 9815 14943
rect 16773 14909 16807 14943
rect 17141 14909 17175 14943
rect 17693 14909 17727 14943
rect 18061 14909 18095 14943
rect 18705 14909 18739 14943
rect 19441 14909 19475 14943
rect 19717 14909 19751 14943
rect 11529 14841 11563 14875
rect 4997 14773 5031 14807
rect 5273 14773 5307 14807
rect 11161 14773 11195 14807
rect 14197 14773 14231 14807
rect 14565 14773 14599 14807
rect 19073 14773 19107 14807
rect 21097 14773 21131 14807
rect 3341 14569 3375 14603
rect 6193 14569 6227 14603
rect 7665 14569 7699 14603
rect 16221 14569 16255 14603
rect 4169 14433 4203 14467
rect 4261 14433 4295 14467
rect 5089 14433 5123 14467
rect 7113 14433 7147 14467
rect 5273 14365 5307 14399
rect 5365 14365 5399 14399
rect 10609 14365 10643 14399
rect 14841 14365 14875 14399
rect 16497 14365 16531 14399
rect 18153 14365 18187 14399
rect 18521 14365 18555 14399
rect 19717 14365 19751 14399
rect 21373 14365 21407 14399
rect 10342 14297 10376 14331
rect 15086 14297 15120 14331
rect 16742 14297 16776 14331
rect 21106 14297 21140 14331
rect 4353 14229 4387 14263
rect 4721 14229 4755 14263
rect 5733 14229 5767 14263
rect 7205 14229 7239 14263
rect 7297 14229 7331 14263
rect 9229 14229 9263 14263
rect 10977 14229 11011 14263
rect 14105 14229 14139 14263
rect 14473 14229 14507 14263
rect 17877 14229 17911 14263
rect 19349 14229 19383 14263
rect 19993 14229 20027 14263
rect 3709 14025 3743 14059
rect 4813 14025 4847 14059
rect 5273 14025 5307 14059
rect 14289 14025 14323 14059
rect 10342 13957 10376 13991
rect 15402 13957 15436 13991
rect 16948 13957 16982 13991
rect 12889 13889 12923 13923
rect 19450 13889 19484 13923
rect 19717 13889 19751 13923
rect 21106 13889 21140 13923
rect 21373 13889 21407 13923
rect 10609 13821 10643 13855
rect 10885 13821 10919 13855
rect 12633 13821 12667 13855
rect 15669 13821 15703 13855
rect 15945 13821 15979 13855
rect 16681 13821 16715 13855
rect 8861 13753 8895 13787
rect 18061 13753 18095 13787
rect 18337 13753 18371 13787
rect 7849 13685 7883 13719
rect 8217 13685 8251 13719
rect 8493 13685 8527 13719
rect 9229 13685 9263 13719
rect 14013 13685 14047 13719
rect 19993 13685 20027 13719
rect 10701 13481 10735 13515
rect 12357 13481 12391 13515
rect 19257 13481 19291 13515
rect 21097 13481 21131 13515
rect 8585 13413 8619 13447
rect 18245 13413 18279 13447
rect 18797 13413 18831 13447
rect 5089 13345 5123 13379
rect 5273 13345 5307 13379
rect 9045 13345 9079 13379
rect 20637 13345 20671 13379
rect 7205 13277 7239 13311
rect 7472 13277 7506 13311
rect 12081 13277 12115 13311
rect 13737 13277 13771 13311
rect 15218 13277 15252 13311
rect 15485 13277 15519 13311
rect 15761 13277 15795 13311
rect 16221 13277 16255 13311
rect 18061 13277 18095 13311
rect 18613 13277 18647 13311
rect 20913 13277 20947 13311
rect 5365 13209 5399 13243
rect 9290 13209 9324 13243
rect 11836 13209 11870 13243
rect 13492 13209 13526 13243
rect 16488 13209 16522 13243
rect 20370 13209 20404 13243
rect 5733 13141 5767 13175
rect 6101 13141 6135 13175
rect 10425 13141 10459 13175
rect 14105 13141 14139 13175
rect 17601 13141 17635 13175
rect 5273 12937 5307 12971
rect 7849 12937 7883 12971
rect 5365 12869 5399 12903
rect 11529 12869 11563 12903
rect 12173 12869 12207 12903
rect 12541 12869 12575 12903
rect 16221 12869 16255 12903
rect 21128 12869 21162 12903
rect 6469 12801 6503 12835
rect 6736 12801 6770 12835
rect 8125 12801 8159 12835
rect 8392 12801 8426 12835
rect 9781 12801 9815 12835
rect 10048 12801 10082 12835
rect 14022 12801 14056 12835
rect 14289 12801 14323 12835
rect 15678 12801 15712 12835
rect 15945 12801 15979 12835
rect 17794 12801 17828 12835
rect 18604 12801 18638 12835
rect 21373 12801 21407 12835
rect 5089 12733 5123 12767
rect 18061 12733 18095 12767
rect 18337 12733 18371 12767
rect 9505 12665 9539 12699
rect 12909 12665 12943 12699
rect 16681 12665 16715 12699
rect 19993 12665 20027 12699
rect 5733 12597 5767 12631
rect 11161 12597 11195 12631
rect 14565 12597 14599 12631
rect 19717 12597 19751 12631
rect 12909 12393 12943 12427
rect 13277 12393 13311 12427
rect 13645 12393 13679 12427
rect 14105 12393 14139 12427
rect 19625 12393 19659 12427
rect 5457 12257 5491 12291
rect 6837 12257 6871 12291
rect 15485 12257 15519 12291
rect 7205 12189 7239 12223
rect 9137 12189 9171 12223
rect 11253 12189 11287 12223
rect 11509 12189 11543 12223
rect 17141 12189 17175 12223
rect 18797 12189 18831 12223
rect 19441 12189 19475 12223
rect 21373 12189 21407 12223
rect 6653 12121 6687 12155
rect 7472 12121 7506 12155
rect 9404 12121 9438 12155
rect 15240 12121 15274 12155
rect 16896 12121 16930 12155
rect 18552 12121 18586 12155
rect 21128 12121 21162 12155
rect 4997 12053 5031 12087
rect 5917 12053 5951 12087
rect 6193 12053 6227 12087
rect 6561 12053 6595 12087
rect 8585 12053 8619 12087
rect 10517 12053 10551 12087
rect 10885 12053 10919 12087
rect 12633 12053 12667 12087
rect 15761 12053 15795 12087
rect 17417 12053 17451 12087
rect 19993 12053 20027 12087
rect 7021 11849 7055 11883
rect 7481 11849 7515 11883
rect 8125 11849 8159 11883
rect 12909 11849 12943 11883
rect 14381 11849 14415 11883
rect 15577 11849 15611 11883
rect 16313 11849 16347 11883
rect 6745 11781 6779 11815
rect 8493 11781 8527 11815
rect 12265 11781 12299 11815
rect 18236 11781 18270 11815
rect 5549 11713 5583 11747
rect 5641 11713 5675 11747
rect 7389 11713 7423 11747
rect 10353 11713 10387 11747
rect 11897 11713 11931 11747
rect 13277 11713 13311 11747
rect 14749 11713 14783 11747
rect 17233 11713 17267 11747
rect 17969 11713 18003 11747
rect 19717 11713 19751 11747
rect 19993 11713 20027 11747
rect 20249 11713 20283 11747
rect 5457 11645 5491 11679
rect 7665 11645 7699 11679
rect 8585 11645 8619 11679
rect 8769 11645 8803 11679
rect 10609 11645 10643 11679
rect 13369 11645 13403 11679
rect 13461 11645 13495 11679
rect 14841 11645 14875 11679
rect 15025 11645 15059 11679
rect 16957 11645 16991 11679
rect 17509 11645 17543 11679
rect 4997 11509 5031 11543
rect 6009 11509 6043 11543
rect 9229 11509 9263 11543
rect 10977 11509 11011 11543
rect 11621 11509 11655 11543
rect 13921 11509 13955 11543
rect 19349 11509 19383 11543
rect 21373 11509 21407 11543
rect 5549 11305 5583 11339
rect 6561 11305 6595 11339
rect 7573 11305 7607 11339
rect 7849 11305 7883 11339
rect 14933 11305 14967 11339
rect 15209 11305 15243 11339
rect 17049 11305 17083 11339
rect 19257 11305 19291 11339
rect 9505 11237 9539 11271
rect 12173 11237 12207 11271
rect 5917 11169 5951 11203
rect 6101 11169 6135 11203
rect 7021 11169 7055 11203
rect 8401 11169 8435 11203
rect 11529 11169 11563 11203
rect 13093 11169 13127 11203
rect 14381 11169 14415 11203
rect 15761 11169 15795 11203
rect 17877 11169 17911 11203
rect 19809 11169 19843 11203
rect 20821 11169 20855 11203
rect 7113 11101 7147 11135
rect 10885 11101 10919 11135
rect 11713 11101 11747 11135
rect 14473 11101 14507 11135
rect 15577 11101 15611 11135
rect 16313 11101 16347 11135
rect 18429 11101 18463 11135
rect 20637 11101 20671 11135
rect 6193 11033 6227 11067
rect 8217 11033 8251 11067
rect 8953 11033 8987 11067
rect 10629 11033 10663 11067
rect 12909 11033 12943 11067
rect 15669 11033 15703 11067
rect 16589 11033 16623 11067
rect 17693 11033 17727 11067
rect 17785 11033 17819 11067
rect 18705 11033 18739 11067
rect 19717 11033 19751 11067
rect 20729 11033 20763 11067
rect 21281 11033 21315 11067
rect 7205 10965 7239 10999
rect 8309 10965 8343 10999
rect 11805 10965 11839 10999
rect 12449 10965 12483 10999
rect 12817 10965 12851 10999
rect 13461 10965 13495 10999
rect 14565 10965 14599 10999
rect 17325 10965 17359 10999
rect 19625 10965 19659 10999
rect 20269 10965 20303 10999
rect 7389 10761 7423 10795
rect 7941 10761 7975 10795
rect 8309 10761 8343 10795
rect 10149 10761 10183 10795
rect 11161 10761 11195 10795
rect 12817 10761 12851 10795
rect 14381 10761 14415 10795
rect 17509 10761 17543 10795
rect 18245 10761 18279 10795
rect 18705 10761 18739 10795
rect 19533 10761 19567 10795
rect 20269 10761 20303 10795
rect 21281 10761 21315 10795
rect 8769 10693 8803 10727
rect 9781 10693 9815 10727
rect 12725 10693 12759 10727
rect 14841 10693 14875 10727
rect 16129 10693 16163 10727
rect 19625 10693 19659 10727
rect 6745 10625 6779 10659
rect 8677 10625 8711 10659
rect 10793 10625 10827 10659
rect 11529 10625 11563 10659
rect 13737 10625 13771 10659
rect 14749 10625 14783 10659
rect 15853 10625 15887 10659
rect 16681 10625 16715 10659
rect 16957 10625 16991 10659
rect 17693 10625 17727 10659
rect 18337 10625 18371 10659
rect 20637 10625 20671 10659
rect 6469 10557 6503 10591
rect 6653 10557 6687 10591
rect 8953 10557 8987 10591
rect 9597 10557 9631 10591
rect 9689 10557 9723 10591
rect 10609 10557 10643 10591
rect 10701 10557 10735 10591
rect 12081 10557 12115 10591
rect 12909 10557 12943 10591
rect 13461 10557 13495 10591
rect 13645 10557 13679 10591
rect 14933 10557 14967 10591
rect 18153 10557 18187 10591
rect 19349 10557 19383 10591
rect 20729 10557 20763 10591
rect 20821 10557 20855 10591
rect 14105 10489 14139 10523
rect 5917 10421 5951 10455
rect 7113 10421 7147 10455
rect 12357 10421 12391 10455
rect 15485 10421 15519 10455
rect 19993 10421 20027 10455
rect 7389 10217 7423 10251
rect 13093 10217 13127 10251
rect 14565 10217 14599 10251
rect 17693 10217 17727 10251
rect 21189 10217 21223 10251
rect 6377 10149 6411 10183
rect 5457 10081 5491 10115
rect 5641 10081 5675 10115
rect 6929 10081 6963 10115
rect 9229 10081 9263 10115
rect 10241 10081 10275 10115
rect 11161 10081 11195 10115
rect 11621 10081 11655 10115
rect 12541 10081 12575 10115
rect 14105 10081 14139 10115
rect 15761 10081 15795 10115
rect 18337 10081 18371 10115
rect 18705 10081 18739 10115
rect 6745 10013 6779 10047
rect 9413 10013 9447 10047
rect 12725 10013 12759 10047
rect 15485 10013 15519 10047
rect 16957 10013 16991 10047
rect 17233 10013 17267 10047
rect 19533 10013 19567 10047
rect 20269 10013 20303 10047
rect 21005 10013 21039 10047
rect 7757 9945 7791 9979
rect 16221 9945 16255 9979
rect 19809 9945 19843 9979
rect 20545 9945 20579 9979
rect 5733 9877 5767 9911
rect 6101 9877 6135 9911
rect 6837 9877 6871 9911
rect 8125 9877 8159 9911
rect 8585 9877 8619 9911
rect 9505 9877 9539 9911
rect 9873 9877 9907 9911
rect 10425 9877 10459 9911
rect 10517 9877 10551 9911
rect 10885 9877 10919 9911
rect 12633 9877 12667 9911
rect 13461 9877 13495 9911
rect 15117 9877 15151 9911
rect 15577 9877 15611 9911
rect 16681 9877 16715 9911
rect 18061 9877 18095 9911
rect 18153 9877 18187 9911
rect 6745 9673 6779 9707
rect 10241 9673 10275 9707
rect 10885 9673 10919 9707
rect 14749 9673 14783 9707
rect 17049 9673 17083 9707
rect 18429 9673 18463 9707
rect 6653 9605 6687 9639
rect 8677 9605 8711 9639
rect 11621 9605 11655 9639
rect 20637 9605 20671 9639
rect 4997 9537 5031 9571
rect 5641 9537 5675 9571
rect 7757 9537 7791 9571
rect 8769 9537 8803 9571
rect 9413 9537 9447 9571
rect 12541 9537 12575 9571
rect 12633 9537 12667 9571
rect 13553 9537 13587 9571
rect 14657 9537 14691 9571
rect 15669 9537 15703 9571
rect 18061 9537 18095 9571
rect 18705 9537 18739 9571
rect 19901 9537 19935 9571
rect 20545 9537 20579 9571
rect 21189 9537 21223 9571
rect 5365 9469 5399 9503
rect 5549 9469 5583 9503
rect 6561 9469 6595 9503
rect 7573 9469 7607 9503
rect 7665 9469 7699 9503
rect 8585 9469 8619 9503
rect 10057 9469 10091 9503
rect 10149 9469 10183 9503
rect 12817 9469 12851 9503
rect 13645 9469 13679 9503
rect 13829 9469 13863 9503
rect 14841 9469 14875 9503
rect 15393 9469 15427 9503
rect 15577 9469 15611 9503
rect 16865 9469 16899 9503
rect 16957 9469 16991 9503
rect 17877 9469 17911 9503
rect 17969 9469 18003 9503
rect 18889 9469 18923 9503
rect 20729 9469 20763 9503
rect 7113 9401 7147 9435
rect 8125 9401 8159 9435
rect 9137 9401 9171 9435
rect 12173 9401 12207 9435
rect 13185 9401 13219 9435
rect 14289 9401 14323 9435
rect 16037 9401 16071 9435
rect 20177 9401 20211 9435
rect 4629 9333 4663 9367
rect 6009 9333 6043 9367
rect 10609 9333 10643 9367
rect 17417 9333 17451 9367
rect 19717 9333 19751 9367
rect 5917 9129 5951 9163
rect 9965 9129 9999 9163
rect 11897 9129 11931 9163
rect 14197 9129 14231 9163
rect 15117 9129 15151 9163
rect 17693 9129 17727 9163
rect 20453 9129 20487 9163
rect 5365 8993 5399 9027
rect 7021 8993 7055 9027
rect 9413 8993 9447 9027
rect 10241 8993 10275 9027
rect 12541 8993 12575 9027
rect 13277 8993 13311 9027
rect 15945 8993 15979 9027
rect 18153 8993 18187 9027
rect 18337 8993 18371 9027
rect 19993 8993 20027 9027
rect 21005 8993 21039 9027
rect 5549 8925 5583 8959
rect 7205 8925 7239 8959
rect 9597 8925 9631 8959
rect 12265 8925 12299 8959
rect 16865 8925 16899 8959
rect 18061 8925 18095 8959
rect 19257 8925 19291 8959
rect 5457 8857 5491 8891
rect 7113 8857 7147 8891
rect 9505 8857 9539 8891
rect 17141 8857 17175 8891
rect 19533 8857 19567 8891
rect 6285 8789 6319 8823
rect 7573 8789 7607 8823
rect 7849 8789 7883 8823
rect 8585 8789 8619 8823
rect 10701 8789 10735 8823
rect 11529 8789 11563 8823
rect 12357 8789 12391 8823
rect 13645 8789 13679 8823
rect 14841 8789 14875 8823
rect 16037 8789 16071 8823
rect 16129 8789 16163 8823
rect 16497 8789 16531 8823
rect 18797 8789 18831 8823
rect 20821 8789 20855 8823
rect 20913 8789 20947 8823
rect 9505 8585 9539 8619
rect 10149 8585 10183 8619
rect 13093 8585 13127 8619
rect 13645 8585 13679 8619
rect 15209 8585 15243 8619
rect 15577 8585 15611 8619
rect 16957 8585 16991 8619
rect 17049 8585 17083 8619
rect 17417 8585 17451 8619
rect 17785 8585 17819 8619
rect 18153 8585 18187 8619
rect 19165 8585 19199 8619
rect 19717 8585 19751 8619
rect 20269 8585 20303 8619
rect 20637 8585 20671 8619
rect 7297 8517 7331 8551
rect 7941 8517 7975 8551
rect 10517 8517 10551 8551
rect 16037 8517 16071 8551
rect 18521 8517 18555 8551
rect 7389 8449 7423 8483
rect 8401 8449 8435 8483
rect 13737 8449 13771 8483
rect 16313 8449 16347 8483
rect 18613 8449 18647 8483
rect 19533 8449 19567 8483
rect 20085 8449 20119 8483
rect 21005 8449 21039 8483
rect 5365 8381 5399 8415
rect 6377 8381 6411 8415
rect 7481 8381 7515 8415
rect 9597 8381 9631 8415
rect 9781 8381 9815 8415
rect 10609 8381 10643 8415
rect 10793 8381 10827 8415
rect 12449 8381 12483 8415
rect 13553 8381 13587 8415
rect 16865 8381 16899 8415
rect 18705 8381 18739 8415
rect 21097 8381 21131 8415
rect 21281 8381 21315 8415
rect 11989 8313 12023 8347
rect 14381 8313 14415 8347
rect 14841 8313 14875 8347
rect 6929 8245 6963 8279
rect 9137 8245 9171 8279
rect 11621 8245 11655 8279
rect 14105 8245 14139 8279
rect 6837 8041 6871 8075
rect 8953 8041 8987 8075
rect 10149 8041 10183 8075
rect 10885 8041 10919 8075
rect 12909 8041 12943 8075
rect 13737 8041 13771 8075
rect 18061 8041 18095 8075
rect 21097 8041 21131 8075
rect 13277 7973 13311 8007
rect 5273 7905 5307 7939
rect 6193 7905 6227 7939
rect 6377 7905 6411 7939
rect 9413 7905 9447 7939
rect 9597 7905 9631 7939
rect 11345 7905 11379 7939
rect 11529 7905 11563 7939
rect 12357 7905 12391 7939
rect 14289 7905 14323 7939
rect 17049 7905 17083 7939
rect 17233 7905 17267 7939
rect 18705 7905 18739 7939
rect 20453 7905 20487 7939
rect 5457 7837 5491 7871
rect 12541 7837 12575 7871
rect 19257 7837 19291 7871
rect 20177 7837 20211 7871
rect 20913 7837 20947 7871
rect 9321 7769 9355 7803
rect 12449 7769 12483 7803
rect 14381 7769 14415 7803
rect 14473 7769 14507 7803
rect 15117 7769 15151 7803
rect 16957 7769 16991 7803
rect 19533 7769 19567 7803
rect 4721 7701 4755 7735
rect 5365 7701 5399 7735
rect 5825 7701 5859 7735
rect 6469 7701 6503 7735
rect 10517 7701 10551 7735
rect 11253 7701 11287 7735
rect 14841 7701 14875 7735
rect 15853 7701 15887 7735
rect 16313 7701 16347 7735
rect 16589 7701 16623 7735
rect 17785 7701 17819 7735
rect 18429 7701 18463 7735
rect 18521 7701 18555 7735
rect 5273 7497 5307 7531
rect 5641 7497 5675 7531
rect 7113 7497 7147 7531
rect 9781 7497 9815 7531
rect 11529 7497 11563 7531
rect 11989 7497 12023 7531
rect 13921 7497 13955 7531
rect 14565 7497 14599 7531
rect 14933 7497 14967 7531
rect 17049 7497 17083 7531
rect 18245 7497 18279 7531
rect 18613 7497 18647 7531
rect 9413 7429 9447 7463
rect 10149 7429 10183 7463
rect 10517 7429 10551 7463
rect 12541 7429 12575 7463
rect 13461 7429 13495 7463
rect 14473 7429 14507 7463
rect 15669 7429 15703 7463
rect 19165 7429 19199 7463
rect 6745 7361 6779 7395
rect 9321 7361 9355 7395
rect 11897 7361 11931 7395
rect 13553 7361 13587 7395
rect 15577 7361 15611 7395
rect 18889 7361 18923 7395
rect 20177 7361 20211 7395
rect 20729 7361 20763 7395
rect 4997 7293 5031 7327
rect 5181 7293 5215 7327
rect 6469 7293 6503 7327
rect 6653 7293 6687 7327
rect 9137 7293 9171 7327
rect 12081 7293 12115 7327
rect 13369 7293 13403 7327
rect 14381 7293 14415 7327
rect 15853 7293 15887 7327
rect 16773 7293 16807 7327
rect 16957 7293 16991 7327
rect 17969 7293 18003 7327
rect 18153 7293 18187 7327
rect 19625 7293 19659 7327
rect 20913 7293 20947 7327
rect 11069 7225 11103 7259
rect 15209 7225 15243 7259
rect 17417 7225 17451 7259
rect 4537 7157 4571 7191
rect 5917 7157 5951 7191
rect 16313 7157 16347 7191
rect 20361 7157 20395 7191
rect 15577 6953 15611 6987
rect 17325 6953 17359 6987
rect 18613 6953 18647 6987
rect 6193 6817 6227 6851
rect 10701 6817 10735 6851
rect 11161 6817 11195 6851
rect 11989 6817 12023 6851
rect 13001 6817 13035 6851
rect 13277 6817 13311 6851
rect 14749 6817 14783 6851
rect 16037 6817 16071 6851
rect 16221 6817 16255 6851
rect 16773 6817 16807 6851
rect 17969 6817 18003 6851
rect 19349 6817 19383 6851
rect 20453 6817 20487 6851
rect 12081 6749 12115 6783
rect 18153 6749 18187 6783
rect 20821 6749 20855 6783
rect 9321 6681 9355 6715
rect 13737 6681 13771 6715
rect 14473 6681 14507 6715
rect 16865 6681 16899 6715
rect 19625 6681 19659 6715
rect 9597 6613 9631 6647
rect 10425 6613 10459 6647
rect 11437 6613 11471 6647
rect 12173 6613 12207 6647
rect 12541 6613 12575 6647
rect 14105 6613 14139 6647
rect 14565 6613 14599 6647
rect 15301 6613 15335 6647
rect 15945 6613 15979 6647
rect 16957 6613 16991 6647
rect 18245 6613 18279 6647
rect 20177 6613 20211 6647
rect 21005 6613 21039 6647
rect 9505 6409 9539 6443
rect 10057 6409 10091 6443
rect 10517 6409 10551 6443
rect 12081 6409 12115 6443
rect 12541 6409 12575 6443
rect 13185 6409 13219 6443
rect 14565 6409 14599 6443
rect 16681 6409 16715 6443
rect 17049 6409 17083 6443
rect 18153 6409 18187 6443
rect 18061 6341 18095 6375
rect 19993 6341 20027 6375
rect 21005 6341 21039 6375
rect 9137 6273 9171 6307
rect 10149 6273 10183 6307
rect 11161 6273 11195 6307
rect 12173 6273 12207 6307
rect 14473 6273 14507 6307
rect 15485 6273 15519 6307
rect 19717 6273 19751 6307
rect 8953 6205 8987 6239
rect 9045 6205 9079 6239
rect 9965 6205 9999 6239
rect 11897 6205 11931 6239
rect 13277 6205 13311 6239
rect 13369 6205 13403 6239
rect 14749 6205 14783 6239
rect 15301 6205 15335 6239
rect 15393 6205 15427 6239
rect 17141 6205 17175 6239
rect 17325 6205 17359 6239
rect 18245 6205 18279 6239
rect 18797 6205 18831 6239
rect 21097 6205 21131 6239
rect 21189 6205 21223 6239
rect 12817 6137 12851 6171
rect 15853 6137 15887 6171
rect 19073 6137 19107 6171
rect 14105 6069 14139 6103
rect 16221 6069 16255 6103
rect 17693 6069 17727 6103
rect 20637 6069 20671 6103
rect 9045 5865 9079 5899
rect 10057 5865 10091 5899
rect 10425 5865 10459 5899
rect 11897 5865 11931 5899
rect 12909 5865 12943 5899
rect 15945 5865 15979 5899
rect 16957 5865 16991 5899
rect 14933 5797 14967 5831
rect 9505 5729 9539 5763
rect 11253 5729 11287 5763
rect 12449 5729 12483 5763
rect 13553 5729 13587 5763
rect 15485 5729 15519 5763
rect 16405 5729 16439 5763
rect 16589 5729 16623 5763
rect 17509 5729 17543 5763
rect 18337 5729 18371 5763
rect 18429 5729 18463 5763
rect 19717 5729 19751 5763
rect 21097 5729 21131 5763
rect 9689 5661 9723 5695
rect 11069 5661 11103 5695
rect 12265 5661 12299 5695
rect 13369 5661 13403 5695
rect 15301 5661 15335 5695
rect 17417 5661 17451 5695
rect 18521 5661 18555 5695
rect 19901 5661 19935 5695
rect 21005 5661 21039 5695
rect 12357 5593 12391 5627
rect 14657 5593 14691 5627
rect 16313 5593 16347 5627
rect 19809 5593 19843 5627
rect 9597 5525 9631 5559
rect 10701 5525 10735 5559
rect 11161 5525 11195 5559
rect 13277 5525 13311 5559
rect 14197 5525 14231 5559
rect 15393 5525 15427 5559
rect 17325 5525 17359 5559
rect 18889 5525 18923 5559
rect 20269 5525 20303 5559
rect 20545 5525 20579 5559
rect 20913 5525 20947 5559
rect 9505 5321 9539 5355
rect 9965 5321 9999 5355
rect 10609 5321 10643 5355
rect 11713 5321 11747 5355
rect 13461 5321 13495 5355
rect 13921 5321 13955 5355
rect 14933 5321 14967 5355
rect 15853 5321 15887 5355
rect 16313 5321 16347 5355
rect 17785 5321 17819 5355
rect 18337 5321 18371 5355
rect 18705 5321 18739 5355
rect 20729 5321 20763 5355
rect 12081 5253 12115 5287
rect 20821 5253 20855 5287
rect 8769 5185 8803 5219
rect 9137 5185 9171 5219
rect 9873 5185 9907 5219
rect 13553 5185 13587 5219
rect 14841 5185 14875 5219
rect 15945 5185 15979 5219
rect 16681 5185 16715 5219
rect 17693 5185 17727 5219
rect 19717 5185 19751 5219
rect 10149 5117 10183 5151
rect 12173 5117 12207 5151
rect 12357 5117 12391 5151
rect 12909 5117 12943 5151
rect 13369 5117 13403 5151
rect 14657 5117 14691 5151
rect 15761 5117 15795 5151
rect 17877 5117 17911 5151
rect 18797 5117 18831 5151
rect 18981 5117 19015 5151
rect 19809 5117 19843 5151
rect 19993 5117 20027 5151
rect 21005 5117 21039 5151
rect 11161 5049 11195 5083
rect 16865 5049 16899 5083
rect 19349 5049 19383 5083
rect 8493 4981 8527 5015
rect 14197 4981 14231 5015
rect 15301 4981 15335 5015
rect 17325 4981 17359 5015
rect 20361 4981 20395 5015
rect 8493 4777 8527 4811
rect 9505 4777 9539 4811
rect 10609 4777 10643 4811
rect 14105 4777 14139 4811
rect 16129 4777 16163 4811
rect 17877 4777 17911 4811
rect 19717 4777 19751 4811
rect 20177 4777 20211 4811
rect 21281 4777 21315 4811
rect 13645 4709 13679 4743
rect 10057 4641 10091 4675
rect 11161 4641 11195 4675
rect 12265 4641 12299 4675
rect 13277 4641 13311 4675
rect 14749 4641 14783 4675
rect 15669 4641 15703 4675
rect 16497 4641 16531 4675
rect 18521 4641 18555 4675
rect 20453 4641 20487 4675
rect 21005 4641 21039 4675
rect 8953 4573 8987 4607
rect 9965 4573 9999 4607
rect 13001 4573 13035 4607
rect 17141 4573 17175 4607
rect 18337 4573 18371 4607
rect 9873 4505 9907 4539
rect 10977 4505 11011 4539
rect 11989 4505 12023 4539
rect 13093 4505 13127 4539
rect 15485 4505 15519 4539
rect 17417 4505 17451 4539
rect 18245 4505 18279 4539
rect 19257 4505 19291 4539
rect 9137 4437 9171 4471
rect 11069 4437 11103 4471
rect 11621 4437 11655 4471
rect 12081 4437 12115 4471
rect 12633 4437 12667 4471
rect 14473 4437 14507 4471
rect 14565 4437 14599 4471
rect 15117 4437 15151 4471
rect 15577 4437 15611 4471
rect 8861 4233 8895 4267
rect 9689 4233 9723 4267
rect 10333 4233 10367 4267
rect 11069 4233 11103 4267
rect 11897 4233 11931 4267
rect 12265 4233 12299 4267
rect 13001 4233 13035 4267
rect 13369 4233 13403 4267
rect 14197 4233 14231 4267
rect 15761 4233 15795 4267
rect 16773 4233 16807 4267
rect 10701 4165 10735 4199
rect 11805 4165 11839 4199
rect 12633 4165 12667 4199
rect 15117 4165 15151 4199
rect 17325 4097 17359 4131
rect 18705 4097 18739 4131
rect 20545 4097 20579 4131
rect 21189 4097 21223 4131
rect 11713 4029 11747 4063
rect 13461 4029 13495 4063
rect 13553 4029 13587 4063
rect 15485 4029 15519 4063
rect 15669 4029 15703 4063
rect 17509 4029 17543 4063
rect 18521 4029 18555 4063
rect 19717 4029 19751 4063
rect 20085 4029 20119 4063
rect 14473 3961 14507 3995
rect 10057 3893 10091 3927
rect 16129 3893 16163 3927
rect 18981 3893 19015 3927
rect 19441 3893 19475 3927
rect 12909 3689 12943 3723
rect 17601 3689 17635 3723
rect 19625 3689 19659 3723
rect 21281 3689 21315 3723
rect 18337 3621 18371 3655
rect 10241 3553 10275 3587
rect 10701 3553 10735 3587
rect 14841 3553 14875 3587
rect 15761 3553 15795 3587
rect 16681 3553 16715 3587
rect 16773 3553 16807 3587
rect 20361 3553 20395 3587
rect 20821 3553 20855 3587
rect 10977 3485 11011 3519
rect 12173 3485 12207 3519
rect 12725 3485 12759 3519
rect 13277 3485 13311 3519
rect 15669 3485 15703 3519
rect 16589 3485 16623 3519
rect 17233 3485 17267 3519
rect 18153 3485 18187 3519
rect 9965 3417 9999 3451
rect 11253 3417 11287 3451
rect 11897 3417 11931 3451
rect 14565 3417 14599 3451
rect 19993 3417 20027 3451
rect 13461 3349 13495 3383
rect 14197 3349 14231 3383
rect 14657 3349 14691 3383
rect 15209 3349 15243 3383
rect 15577 3349 15611 3383
rect 16221 3349 16255 3383
rect 18705 3349 18739 3383
rect 19349 3349 19383 3383
rect 9413 3145 9447 3179
rect 9873 3145 9907 3179
rect 10149 3145 10183 3179
rect 10609 3145 10643 3179
rect 13829 3145 13863 3179
rect 14197 3145 14231 3179
rect 14841 3145 14875 3179
rect 15301 3145 15335 3179
rect 17693 3145 17727 3179
rect 18797 3145 18831 3179
rect 14289 3077 14323 3111
rect 15209 3077 15243 3111
rect 11161 3009 11195 3043
rect 11897 3009 11931 3043
rect 13277 3009 13311 3043
rect 15945 3009 15979 3043
rect 16957 3009 16991 3043
rect 17509 3009 17543 3043
rect 18337 3009 18371 3043
rect 18613 3009 18647 3043
rect 19165 3009 19199 3043
rect 19717 3009 19751 3043
rect 20821 3009 20855 3043
rect 11529 2941 11563 2975
rect 12173 2941 12207 2975
rect 13093 2941 13127 2975
rect 14473 2941 14507 2975
rect 15485 2941 15519 2975
rect 20269 2941 20303 2975
rect 10977 2873 11011 2907
rect 16129 2873 16163 2907
rect 18153 2873 18187 2907
rect 19349 2873 19383 2907
rect 19901 2873 19935 2907
rect 16773 2805 16807 2839
rect 21005 2805 21039 2839
rect 10701 2601 10735 2635
rect 11161 2601 11195 2635
rect 11713 2601 11747 2635
rect 13645 2601 13679 2635
rect 15945 2601 15979 2635
rect 17141 2601 17175 2635
rect 18705 2601 18739 2635
rect 19625 2601 19659 2635
rect 19993 2601 20027 2635
rect 21281 2601 21315 2635
rect 10425 2533 10459 2567
rect 15117 2533 15151 2567
rect 16865 2533 16899 2567
rect 18337 2533 18371 2567
rect 16221 2465 16255 2499
rect 17509 2465 17543 2499
rect 19257 2465 19291 2499
rect 11989 2397 12023 2431
rect 12541 2397 12575 2431
rect 13093 2397 13127 2431
rect 14105 2397 14139 2431
rect 14933 2397 14967 2431
rect 18153 2397 18187 2431
rect 20729 2397 20763 2431
rect 10057 2329 10091 2363
rect 12173 2261 12207 2295
rect 12725 2261 12759 2295
rect 13277 2261 13311 2295
rect 14289 2261 14323 2295
rect 15485 2261 15519 2295
rect 20361 2261 20395 2295
<< metal1 >>
rect 10226 21020 10232 21072
rect 10284 21060 10290 21072
rect 11974 21060 11980 21072
rect 10284 21032 11980 21060
rect 10284 21020 10290 21032
rect 11974 21020 11980 21032
rect 12032 21020 12038 21072
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 7929 20587 7987 20593
rect 7929 20553 7941 20587
rect 7975 20584 7987 20587
rect 8481 20587 8539 20593
rect 7975 20556 8432 20584
rect 7975 20553 7987 20556
rect 7929 20547 7987 20553
rect 6546 20476 6552 20528
rect 6604 20516 6610 20528
rect 6604 20488 8340 20516
rect 6604 20476 6610 20488
rect 6641 20451 6699 20457
rect 6641 20417 6653 20451
rect 6687 20448 6699 20451
rect 6730 20448 6736 20460
rect 6687 20420 6736 20448
rect 6687 20417 6699 20420
rect 6641 20411 6699 20417
rect 6730 20408 6736 20420
rect 6788 20408 6794 20460
rect 7193 20451 7251 20457
rect 7193 20417 7205 20451
rect 7239 20417 7251 20451
rect 7742 20448 7748 20460
rect 7703 20420 7748 20448
rect 7193 20411 7251 20417
rect 7208 20380 7236 20411
rect 7742 20408 7748 20420
rect 7800 20408 7806 20460
rect 8312 20457 8340 20488
rect 8297 20451 8355 20457
rect 8297 20417 8309 20451
rect 8343 20417 8355 20451
rect 8404 20448 8432 20556
rect 8481 20553 8493 20587
rect 8527 20553 8539 20587
rect 8481 20547 8539 20553
rect 9309 20587 9367 20593
rect 9309 20553 9321 20587
rect 9355 20584 9367 20587
rect 11609 20587 11667 20593
rect 11609 20584 11621 20587
rect 9355 20556 11621 20584
rect 9355 20553 9367 20556
rect 9309 20547 9367 20553
rect 11609 20553 11621 20556
rect 11655 20584 11667 20587
rect 11698 20584 11704 20596
rect 11655 20556 11704 20584
rect 11655 20553 11667 20556
rect 11609 20547 11667 20553
rect 8496 20516 8524 20547
rect 11698 20544 11704 20556
rect 11756 20544 11762 20596
rect 14277 20587 14335 20593
rect 14277 20553 14289 20587
rect 14323 20584 14335 20587
rect 18598 20584 18604 20596
rect 14323 20556 18604 20584
rect 14323 20553 14335 20556
rect 14277 20547 14335 20553
rect 18598 20544 18604 20556
rect 18656 20544 18662 20596
rect 18690 20544 18696 20596
rect 18748 20584 18754 20596
rect 19429 20587 19487 20593
rect 18748 20556 18793 20584
rect 18748 20544 18754 20556
rect 19429 20553 19441 20587
rect 19475 20584 19487 20587
rect 21358 20584 21364 20596
rect 19475 20556 21364 20584
rect 19475 20553 19487 20556
rect 19429 20547 19487 20553
rect 21358 20544 21364 20556
rect 21416 20544 21422 20596
rect 12989 20519 13047 20525
rect 8496 20488 12434 20516
rect 10226 20448 10232 20460
rect 8404 20420 10232 20448
rect 8297 20411 8355 20417
rect 10226 20408 10232 20420
rect 10284 20408 10290 20460
rect 10502 20408 10508 20460
rect 10560 20448 10566 20460
rect 12406 20448 12434 20488
rect 12989 20485 13001 20519
rect 13035 20516 13047 20519
rect 13035 20488 16574 20516
rect 13035 20485 13047 20488
rect 12989 20479 13047 20485
rect 12618 20448 12624 20460
rect 10560 20420 10605 20448
rect 12406 20420 12624 20448
rect 10560 20408 10566 20420
rect 12618 20408 12624 20420
rect 12676 20408 12682 20460
rect 14093 20451 14151 20457
rect 14093 20417 14105 20451
rect 14139 20417 14151 20451
rect 14093 20411 14151 20417
rect 5644 20352 7236 20380
rect 5644 20256 5672 20352
rect 7374 20340 7380 20392
rect 7432 20380 7438 20392
rect 7558 20380 7564 20392
rect 7432 20352 7564 20380
rect 7432 20340 7438 20352
rect 7558 20340 7564 20352
rect 7616 20380 7622 20392
rect 9401 20383 9459 20389
rect 9401 20380 9413 20383
rect 7616 20352 9413 20380
rect 7616 20340 7622 20352
rect 9401 20349 9413 20352
rect 9447 20349 9459 20383
rect 9401 20343 9459 20349
rect 9585 20383 9643 20389
rect 9585 20349 9597 20383
rect 9631 20349 9643 20383
rect 9585 20343 9643 20349
rect 10321 20383 10379 20389
rect 10321 20349 10333 20383
rect 10367 20380 10379 20383
rect 14108 20380 14136 20411
rect 14642 20408 14648 20460
rect 14700 20448 14706 20460
rect 15013 20451 15071 20457
rect 15013 20448 15025 20451
rect 14700 20420 15025 20448
rect 14700 20408 14706 20420
rect 15013 20417 15025 20420
rect 15059 20417 15071 20451
rect 15654 20448 15660 20460
rect 15615 20420 15660 20448
rect 15013 20411 15071 20417
rect 15654 20408 15660 20420
rect 15712 20408 15718 20460
rect 15672 20380 15700 20408
rect 10367 20352 10456 20380
rect 10367 20349 10379 20352
rect 10321 20343 10379 20349
rect 9600 20312 9628 20343
rect 9600 20284 10364 20312
rect 10336 20256 10364 20284
rect 5626 20244 5632 20256
rect 5587 20216 5632 20244
rect 5626 20204 5632 20216
rect 5684 20204 5690 20256
rect 5997 20247 6055 20253
rect 5997 20213 6009 20247
rect 6043 20244 6055 20247
rect 6546 20244 6552 20256
rect 6043 20216 6552 20244
rect 6043 20213 6055 20216
rect 5997 20207 6055 20213
rect 6546 20204 6552 20216
rect 6604 20204 6610 20256
rect 6825 20247 6883 20253
rect 6825 20213 6837 20247
rect 6871 20244 6883 20247
rect 7282 20244 7288 20256
rect 6871 20216 7288 20244
rect 6871 20213 6883 20216
rect 6825 20207 6883 20213
rect 7282 20204 7288 20216
rect 7340 20204 7346 20256
rect 7377 20247 7435 20253
rect 7377 20213 7389 20247
rect 7423 20244 7435 20247
rect 8386 20244 8392 20256
rect 7423 20216 8392 20244
rect 7423 20213 7435 20216
rect 7377 20207 7435 20213
rect 8386 20204 8392 20216
rect 8444 20204 8450 20256
rect 8570 20204 8576 20256
rect 8628 20244 8634 20256
rect 8941 20247 8999 20253
rect 8941 20244 8953 20247
rect 8628 20216 8953 20244
rect 8628 20204 8634 20216
rect 8941 20213 8953 20216
rect 8987 20213 8999 20247
rect 8941 20207 8999 20213
rect 10318 20204 10324 20256
rect 10376 20204 10382 20256
rect 10428 20244 10456 20352
rect 10796 20352 14136 20380
rect 14476 20352 15700 20380
rect 16546 20380 16574 20488
rect 17586 20476 17592 20528
rect 17644 20516 17650 20528
rect 20254 20516 20260 20528
rect 17644 20488 18552 20516
rect 17644 20476 17650 20488
rect 16669 20451 16727 20457
rect 16669 20417 16681 20451
rect 16715 20448 16727 20451
rect 17681 20451 17739 20457
rect 16715 20420 16749 20448
rect 16715 20417 16727 20420
rect 16669 20411 16727 20417
rect 17681 20417 17693 20451
rect 17727 20448 17739 20451
rect 18138 20448 18144 20460
rect 17727 20420 18144 20448
rect 17727 20417 17739 20420
rect 17681 20411 17739 20417
rect 16684 20380 16712 20411
rect 18138 20408 18144 20420
rect 18196 20408 18202 20460
rect 18233 20451 18291 20457
rect 18233 20417 18245 20451
rect 18279 20448 18291 20451
rect 18414 20448 18420 20460
rect 18279 20420 18420 20448
rect 18279 20417 18291 20420
rect 18233 20411 18291 20417
rect 18414 20408 18420 20420
rect 18472 20408 18478 20460
rect 18524 20457 18552 20488
rect 18708 20488 20260 20516
rect 18509 20451 18567 20457
rect 18509 20417 18521 20451
rect 18555 20417 18567 20451
rect 18509 20411 18567 20417
rect 16758 20380 16764 20392
rect 16546 20352 16764 20380
rect 10796 20244 10824 20352
rect 13722 20312 13728 20324
rect 13683 20284 13728 20312
rect 13722 20272 13728 20284
rect 13780 20272 13786 20324
rect 10428 20216 10824 20244
rect 10873 20247 10931 20253
rect 10873 20213 10885 20247
rect 10919 20244 10931 20247
rect 10962 20244 10968 20256
rect 10919 20216 10968 20244
rect 10919 20213 10931 20216
rect 10873 20207 10931 20213
rect 10962 20204 10968 20216
rect 11020 20204 11026 20256
rect 12158 20244 12164 20256
rect 12119 20216 12164 20244
rect 12158 20204 12164 20216
rect 12216 20204 12222 20256
rect 12621 20247 12679 20253
rect 12621 20213 12633 20247
rect 12667 20244 12679 20247
rect 12710 20244 12716 20256
rect 12667 20216 12716 20244
rect 12667 20213 12679 20216
rect 12621 20207 12679 20213
rect 12710 20204 12716 20216
rect 12768 20204 12774 20256
rect 13357 20247 13415 20253
rect 13357 20213 13369 20247
rect 13403 20244 13415 20247
rect 14476 20244 14504 20352
rect 16758 20340 16764 20352
rect 16816 20340 16822 20392
rect 18708 20380 18736 20488
rect 20254 20476 20260 20488
rect 20312 20476 20318 20528
rect 18874 20408 18880 20460
rect 18932 20448 18938 20460
rect 19245 20451 19303 20457
rect 19245 20448 19257 20451
rect 18932 20420 19257 20448
rect 18932 20408 18938 20420
rect 19245 20417 19257 20420
rect 19291 20417 19303 20451
rect 20806 20448 20812 20460
rect 19245 20411 19303 20417
rect 19444 20420 20812 20448
rect 16868 20352 18736 20380
rect 15841 20315 15899 20321
rect 15841 20281 15853 20315
rect 15887 20312 15899 20315
rect 16298 20312 16304 20324
rect 15887 20284 16304 20312
rect 15887 20281 15899 20284
rect 15841 20275 15899 20281
rect 16298 20272 16304 20284
rect 16356 20272 16362 20324
rect 16868 20321 16896 20352
rect 16853 20315 16911 20321
rect 16853 20281 16865 20315
rect 16899 20281 16911 20315
rect 16853 20275 16911 20281
rect 18049 20315 18107 20321
rect 18049 20281 18061 20315
rect 18095 20312 18107 20315
rect 19444 20312 19472 20420
rect 20806 20408 20812 20420
rect 20864 20408 20870 20460
rect 21082 20448 21088 20460
rect 21140 20457 21146 20460
rect 21052 20420 21088 20448
rect 21082 20408 21088 20420
rect 21140 20411 21152 20457
rect 21140 20408 21146 20411
rect 21358 20380 21364 20392
rect 21319 20352 21364 20380
rect 21358 20340 21364 20352
rect 21416 20340 21422 20392
rect 20162 20312 20168 20324
rect 18095 20284 19472 20312
rect 19505 20284 20168 20312
rect 18095 20281 18107 20284
rect 18049 20275 18107 20281
rect 14642 20244 14648 20256
rect 13403 20216 14504 20244
rect 14603 20216 14648 20244
rect 13403 20213 13415 20216
rect 13357 20207 13415 20213
rect 14642 20204 14648 20216
rect 14700 20204 14706 20256
rect 15197 20247 15255 20253
rect 15197 20213 15209 20247
rect 15243 20244 15255 20247
rect 15930 20244 15936 20256
rect 15243 20216 15936 20244
rect 15243 20213 15255 20216
rect 15197 20207 15255 20213
rect 15930 20204 15936 20216
rect 15988 20204 15994 20256
rect 16206 20244 16212 20256
rect 16167 20216 16212 20244
rect 16206 20204 16212 20216
rect 16264 20204 16270 20256
rect 17497 20247 17555 20253
rect 17497 20213 17509 20247
rect 17543 20244 17555 20247
rect 17954 20244 17960 20256
rect 17543 20216 17960 20244
rect 17543 20213 17555 20216
rect 17497 20207 17555 20213
rect 17954 20204 17960 20216
rect 18012 20204 18018 20256
rect 18138 20204 18144 20256
rect 18196 20244 18202 20256
rect 19505 20244 19533 20284
rect 20162 20272 20168 20284
rect 20220 20272 20226 20324
rect 19978 20244 19984 20256
rect 18196 20216 19533 20244
rect 19939 20216 19984 20244
rect 18196 20204 18202 20216
rect 19978 20204 19984 20216
rect 20036 20204 20042 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 7929 20043 7987 20049
rect 7929 20009 7941 20043
rect 7975 20040 7987 20043
rect 13078 20040 13084 20052
rect 7975 20012 13084 20040
rect 7975 20009 7987 20012
rect 7929 20003 7987 20009
rect 13078 20000 13084 20012
rect 13136 20000 13142 20052
rect 16132 20012 18000 20040
rect 5718 19932 5724 19984
rect 5776 19972 5782 19984
rect 5776 19944 8340 19972
rect 5776 19932 5782 19944
rect 6730 19904 6736 19916
rect 6691 19876 6736 19904
rect 6730 19864 6736 19876
rect 6788 19864 6794 19916
rect 4433 19839 4491 19845
rect 4433 19805 4445 19839
rect 4479 19836 4491 19839
rect 6273 19839 6331 19845
rect 4479 19808 5120 19836
rect 4479 19805 4491 19808
rect 4433 19799 4491 19805
rect 4614 19700 4620 19712
rect 4575 19672 4620 19700
rect 4614 19660 4620 19672
rect 4672 19660 4678 19712
rect 5092 19709 5120 19808
rect 6273 19805 6285 19839
rect 6319 19805 6331 19839
rect 7006 19836 7012 19848
rect 6967 19808 7012 19836
rect 6273 19799 6331 19805
rect 6288 19768 6316 19799
rect 7006 19796 7012 19808
rect 7064 19796 7070 19848
rect 7190 19796 7196 19848
rect 7248 19836 7254 19848
rect 8312 19845 8340 19944
rect 11974 19864 11980 19916
rect 12032 19904 12038 19916
rect 12032 19876 13400 19904
rect 12032 19864 12038 19876
rect 7745 19839 7803 19845
rect 7745 19836 7757 19839
rect 7248 19808 7757 19836
rect 7248 19796 7254 19808
rect 7745 19805 7757 19808
rect 7791 19805 7803 19839
rect 7745 19799 7803 19805
rect 8297 19839 8355 19845
rect 8297 19805 8309 19839
rect 8343 19805 8355 19839
rect 8297 19799 8355 19805
rect 10597 19839 10655 19845
rect 10597 19805 10609 19839
rect 10643 19836 10655 19839
rect 10873 19839 10931 19845
rect 10873 19836 10885 19839
rect 10643 19808 10885 19836
rect 10643 19805 10655 19808
rect 10597 19799 10655 19805
rect 10873 19805 10885 19808
rect 10919 19836 10931 19839
rect 10962 19836 10968 19848
rect 10919 19808 10968 19836
rect 10919 19805 10931 19808
rect 10873 19799 10931 19805
rect 10962 19796 10968 19808
rect 11020 19796 11026 19848
rect 12897 19839 12955 19845
rect 12897 19836 12909 19839
rect 11072 19808 12909 19836
rect 7098 19768 7104 19780
rect 6288 19740 7104 19768
rect 7098 19728 7104 19740
rect 7156 19728 7162 19780
rect 8496 19740 10272 19768
rect 5077 19703 5135 19709
rect 5077 19669 5089 19703
rect 5123 19700 5135 19703
rect 5166 19700 5172 19712
rect 5123 19672 5172 19700
rect 5123 19669 5135 19672
rect 5077 19663 5135 19669
rect 5166 19660 5172 19672
rect 5224 19660 5230 19712
rect 5718 19700 5724 19712
rect 5679 19672 5724 19700
rect 5718 19660 5724 19672
rect 5776 19660 5782 19712
rect 6089 19703 6147 19709
rect 6089 19669 6101 19703
rect 6135 19700 6147 19703
rect 6914 19700 6920 19712
rect 6135 19672 6920 19700
rect 6135 19669 6147 19672
rect 6089 19663 6147 19669
rect 6914 19660 6920 19672
rect 6972 19660 6978 19712
rect 7374 19700 7380 19712
rect 7335 19672 7380 19700
rect 7374 19660 7380 19672
rect 7432 19660 7438 19712
rect 8496 19709 8524 19740
rect 8481 19703 8539 19709
rect 8481 19669 8493 19703
rect 8527 19669 8539 19703
rect 8481 19663 8539 19669
rect 9217 19703 9275 19709
rect 9217 19669 9229 19703
rect 9263 19700 9275 19703
rect 9306 19700 9312 19712
rect 9263 19672 9312 19700
rect 9263 19669 9275 19672
rect 9217 19663 9275 19669
rect 9306 19660 9312 19672
rect 9364 19660 9370 19712
rect 10244 19700 10272 19740
rect 10318 19728 10324 19780
rect 10376 19777 10382 19780
rect 10376 19768 10388 19777
rect 10376 19740 10421 19768
rect 10376 19731 10388 19740
rect 10376 19728 10382 19731
rect 10686 19728 10692 19780
rect 10744 19768 10750 19780
rect 11072 19768 11100 19808
rect 12897 19805 12909 19808
rect 12943 19836 12955 19839
rect 13265 19839 13323 19845
rect 13265 19836 13277 19839
rect 12943 19808 13277 19836
rect 12943 19805 12955 19808
rect 12897 19799 12955 19805
rect 13265 19805 13277 19808
rect 13311 19805 13323 19839
rect 13372 19836 13400 19876
rect 15470 19836 15476 19848
rect 13372 19808 15332 19836
rect 15431 19808 15476 19836
rect 13265 19799 13323 19805
rect 10744 19740 11100 19768
rect 11140 19771 11198 19777
rect 10744 19728 10750 19740
rect 11140 19737 11152 19771
rect 11186 19768 11198 19771
rect 11186 19740 11376 19768
rect 11186 19737 11198 19740
rect 11140 19731 11198 19737
rect 11054 19700 11060 19712
rect 10244 19672 11060 19700
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 11348 19700 11376 19740
rect 11514 19728 11520 19780
rect 11572 19768 11578 19780
rect 13630 19768 13636 19780
rect 11572 19740 13636 19768
rect 11572 19728 11578 19740
rect 13630 19728 13636 19740
rect 13688 19728 13694 19780
rect 13740 19740 14596 19768
rect 11422 19700 11428 19712
rect 11348 19672 11428 19700
rect 11422 19660 11428 19672
rect 11480 19660 11486 19712
rect 12250 19700 12256 19712
rect 12211 19672 12256 19700
rect 12250 19660 12256 19672
rect 12308 19660 12314 19712
rect 12526 19700 12532 19712
rect 12487 19672 12532 19700
rect 12526 19660 12532 19672
rect 12584 19660 12590 19712
rect 13449 19703 13507 19709
rect 13449 19669 13461 19703
rect 13495 19700 13507 19703
rect 13740 19700 13768 19740
rect 13495 19672 13768 19700
rect 13495 19669 13507 19672
rect 13449 19663 13507 19669
rect 13814 19660 13820 19712
rect 13872 19700 13878 19712
rect 14093 19703 14151 19709
rect 14093 19700 14105 19703
rect 13872 19672 14105 19700
rect 13872 19660 13878 19672
rect 14093 19669 14105 19672
rect 14139 19669 14151 19703
rect 14568 19700 14596 19740
rect 14642 19728 14648 19780
rect 14700 19768 14706 19780
rect 15206 19771 15264 19777
rect 15206 19768 15218 19771
rect 14700 19740 15218 19768
rect 14700 19728 14706 19740
rect 15206 19737 15218 19740
rect 15252 19737 15264 19771
rect 15304 19768 15332 19808
rect 15470 19796 15476 19808
rect 15528 19796 15534 19848
rect 15562 19796 15568 19848
rect 15620 19836 15626 19848
rect 15933 19839 15991 19845
rect 15933 19836 15945 19839
rect 15620 19808 15945 19836
rect 15620 19796 15626 19808
rect 15933 19805 15945 19808
rect 15979 19805 15991 19839
rect 15933 19799 15991 19805
rect 16132 19768 16160 20012
rect 17586 19972 17592 19984
rect 16546 19944 17592 19972
rect 16209 19907 16267 19913
rect 16209 19873 16221 19907
rect 16255 19904 16267 19907
rect 16546 19904 16574 19944
rect 17586 19932 17592 19944
rect 17644 19932 17650 19984
rect 16255 19876 16574 19904
rect 16945 19907 17003 19913
rect 16255 19873 16267 19876
rect 16209 19867 16267 19873
rect 16945 19873 16957 19907
rect 16991 19904 17003 19907
rect 17972 19904 18000 20012
rect 18046 20000 18052 20052
rect 18104 20040 18110 20052
rect 18601 20043 18659 20049
rect 18601 20040 18613 20043
rect 18104 20012 18613 20040
rect 18104 20000 18110 20012
rect 18601 20009 18613 20012
rect 18647 20009 18659 20043
rect 18601 20003 18659 20009
rect 18690 20000 18696 20052
rect 18748 20040 18754 20052
rect 21082 20040 21088 20052
rect 18748 20012 21088 20040
rect 18748 20000 18754 20012
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 16991 19876 17448 19904
rect 17972 19876 18368 19904
rect 16991 19873 17003 19876
rect 16945 19867 17003 19873
rect 17034 19836 17040 19848
rect 15304 19740 16160 19768
rect 16224 19808 17040 19836
rect 15206 19731 15264 19737
rect 16224 19700 16252 19808
rect 17034 19796 17040 19808
rect 17092 19796 17098 19848
rect 17129 19839 17187 19845
rect 17129 19805 17141 19839
rect 17175 19836 17187 19839
rect 17310 19836 17316 19848
rect 17175 19808 17316 19836
rect 17175 19805 17187 19808
rect 17129 19799 17187 19805
rect 17310 19796 17316 19808
rect 17368 19796 17374 19848
rect 17420 19845 17448 19876
rect 17405 19839 17463 19845
rect 17405 19805 17417 19839
rect 17451 19805 17463 19839
rect 18230 19836 18236 19848
rect 18191 19808 18236 19836
rect 17405 19799 17463 19805
rect 18230 19796 18236 19808
rect 18288 19796 18294 19848
rect 16942 19728 16948 19780
rect 17000 19768 17006 19780
rect 17000 19740 18092 19768
rect 17000 19728 17006 19740
rect 14568 19672 16252 19700
rect 14093 19663 14151 19669
rect 16390 19660 16396 19712
rect 16448 19700 16454 19712
rect 18064 19709 18092 19740
rect 17589 19703 17647 19709
rect 17589 19700 17601 19703
rect 16448 19672 17601 19700
rect 16448 19660 16454 19672
rect 17589 19669 17601 19672
rect 17635 19669 17647 19703
rect 17589 19663 17647 19669
rect 18049 19703 18107 19709
rect 18049 19669 18061 19703
rect 18095 19669 18107 19703
rect 18340 19700 18368 19876
rect 18414 19864 18420 19916
rect 18472 19904 18478 19916
rect 19429 19907 19487 19913
rect 19429 19904 19441 19907
rect 18472 19876 19441 19904
rect 18472 19864 18478 19876
rect 19429 19873 19441 19876
rect 19475 19873 19487 19907
rect 21358 19904 21364 19916
rect 21319 19876 21364 19904
rect 19429 19867 19487 19873
rect 21358 19864 21364 19876
rect 21416 19864 21422 19916
rect 18782 19836 18788 19848
rect 18743 19808 18788 19836
rect 18782 19796 18788 19808
rect 18840 19796 18846 19848
rect 19245 19839 19303 19845
rect 19245 19805 19257 19839
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 18414 19728 18420 19780
rect 18472 19768 18478 19780
rect 19260 19768 19288 19799
rect 18472 19740 19288 19768
rect 18472 19728 18478 19740
rect 19702 19728 19708 19780
rect 19760 19768 19766 19780
rect 21094 19771 21152 19777
rect 21094 19768 21106 19771
rect 19760 19740 21106 19768
rect 19760 19728 19766 19740
rect 21094 19737 21106 19740
rect 21140 19737 21152 19771
rect 21094 19731 21152 19737
rect 19981 19703 20039 19709
rect 19981 19700 19993 19703
rect 18340 19672 19993 19700
rect 18049 19663 18107 19669
rect 19981 19669 19993 19672
rect 20027 19669 20039 19703
rect 19981 19663 20039 19669
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 5350 19456 5356 19508
rect 5408 19496 5414 19508
rect 6365 19499 6423 19505
rect 6365 19496 6377 19499
rect 5408 19468 6377 19496
rect 5408 19456 5414 19468
rect 6365 19465 6377 19468
rect 6411 19465 6423 19499
rect 6365 19459 6423 19465
rect 6733 19499 6791 19505
rect 6733 19465 6745 19499
rect 6779 19496 6791 19499
rect 6822 19496 6828 19508
rect 6779 19468 6828 19496
rect 6779 19465 6791 19468
rect 6733 19459 6791 19465
rect 6822 19456 6828 19468
rect 6880 19456 6886 19508
rect 8113 19499 8171 19505
rect 7484 19468 8064 19496
rect 4982 19388 4988 19440
rect 5040 19428 5046 19440
rect 7484 19428 7512 19468
rect 5040 19400 7512 19428
rect 7561 19431 7619 19437
rect 5040 19388 5046 19400
rect 7561 19397 7573 19431
rect 7607 19428 7619 19431
rect 7742 19428 7748 19440
rect 7607 19400 7748 19428
rect 7607 19397 7619 19400
rect 7561 19391 7619 19397
rect 7742 19388 7748 19400
rect 7800 19388 7806 19440
rect 5626 19360 5632 19372
rect 5587 19332 5632 19360
rect 5626 19320 5632 19332
rect 5684 19320 5690 19372
rect 5721 19363 5779 19369
rect 5721 19329 5733 19363
rect 5767 19329 5779 19363
rect 7834 19360 7840 19372
rect 7795 19332 7840 19360
rect 5721 19323 5779 19329
rect 4798 19252 4804 19304
rect 4856 19292 4862 19304
rect 4893 19295 4951 19301
rect 4893 19292 4905 19295
rect 4856 19264 4905 19292
rect 4856 19252 4862 19264
rect 4893 19261 4905 19264
rect 4939 19292 4951 19295
rect 5736 19292 5764 19323
rect 7834 19320 7840 19332
rect 7892 19320 7898 19372
rect 8036 19360 8064 19468
rect 8113 19465 8125 19499
rect 8159 19465 8171 19499
rect 8113 19459 8171 19465
rect 11149 19499 11207 19505
rect 11149 19465 11161 19499
rect 11195 19496 11207 19499
rect 12066 19496 12072 19508
rect 11195 19468 12072 19496
rect 11195 19465 11207 19468
rect 11149 19459 11207 19465
rect 8128 19428 8156 19459
rect 12066 19456 12072 19468
rect 12124 19456 12130 19508
rect 12989 19499 13047 19505
rect 12989 19496 13001 19499
rect 12176 19468 13001 19496
rect 8202 19428 8208 19440
rect 8128 19400 8208 19428
rect 8202 19388 8208 19400
rect 8260 19428 8266 19440
rect 10014 19431 10072 19437
rect 10014 19428 10026 19431
rect 8260 19400 10026 19428
rect 8260 19388 8266 19400
rect 10014 19397 10026 19400
rect 10060 19397 10072 19431
rect 10014 19391 10072 19397
rect 10318 19388 10324 19440
rect 10376 19428 10382 19440
rect 12176 19428 12204 19468
rect 12989 19465 13001 19468
rect 13035 19465 13047 19499
rect 14642 19496 14648 19508
rect 14603 19468 14648 19496
rect 12989 19459 13047 19465
rect 14642 19456 14648 19468
rect 14700 19456 14706 19508
rect 16942 19456 16948 19508
rect 17000 19496 17006 19508
rect 18693 19499 18751 19505
rect 18693 19496 18705 19499
rect 17000 19468 18705 19496
rect 17000 19456 17006 19468
rect 18693 19465 18705 19468
rect 18739 19465 18751 19499
rect 18693 19459 18751 19465
rect 18966 19456 18972 19508
rect 19024 19496 19030 19508
rect 20530 19496 20536 19508
rect 19024 19468 20536 19496
rect 19024 19456 19030 19468
rect 20530 19456 20536 19468
rect 20588 19456 20594 19508
rect 10376 19400 12204 19428
rect 12345 19431 12403 19437
rect 10376 19388 10382 19400
rect 12345 19397 12357 19431
rect 12391 19428 12403 19431
rect 12526 19428 12532 19440
rect 12391 19400 12532 19428
rect 12391 19397 12403 19400
rect 12345 19391 12403 19397
rect 12526 19388 12532 19400
rect 12584 19428 12590 19440
rect 12713 19431 12771 19437
rect 12713 19428 12725 19431
rect 12584 19400 12725 19428
rect 12584 19388 12590 19400
rect 12713 19397 12725 19400
rect 12759 19428 12771 19431
rect 13722 19428 13728 19440
rect 12759 19400 13728 19428
rect 12759 19397 12771 19400
rect 12713 19391 12771 19397
rect 13722 19388 13728 19400
rect 13780 19428 13786 19440
rect 13780 19400 14412 19428
rect 13780 19388 13786 19400
rect 9226 19363 9284 19369
rect 9226 19360 9238 19363
rect 8036 19332 9238 19360
rect 9226 19329 9238 19332
rect 9272 19360 9284 19363
rect 9272 19332 10824 19360
rect 9272 19329 9284 19332
rect 9226 19323 9284 19329
rect 4939 19264 5764 19292
rect 5905 19295 5963 19301
rect 4939 19261 4951 19264
rect 4893 19255 4951 19261
rect 5905 19261 5917 19295
rect 5951 19261 5963 19295
rect 5905 19255 5963 19261
rect 5920 19224 5948 19255
rect 5994 19252 6000 19304
rect 6052 19292 6058 19304
rect 6825 19295 6883 19301
rect 6825 19292 6837 19295
rect 6052 19264 6837 19292
rect 6052 19252 6058 19264
rect 6825 19261 6837 19264
rect 6871 19261 6883 19295
rect 6825 19255 6883 19261
rect 7009 19295 7067 19301
rect 7009 19261 7021 19295
rect 7055 19292 7067 19295
rect 8202 19292 8208 19304
rect 7055 19264 8208 19292
rect 7055 19261 7067 19264
rect 7009 19255 7067 19261
rect 8202 19252 8208 19264
rect 8260 19252 8266 19304
rect 9493 19295 9551 19301
rect 9493 19261 9505 19295
rect 9539 19292 9551 19295
rect 9674 19292 9680 19304
rect 9539 19264 9680 19292
rect 9539 19261 9551 19264
rect 9493 19255 9551 19261
rect 9674 19252 9680 19264
rect 9732 19292 9738 19304
rect 9769 19295 9827 19301
rect 9769 19292 9781 19295
rect 9732 19264 9781 19292
rect 9732 19252 9738 19264
rect 9769 19261 9781 19264
rect 9815 19261 9827 19295
rect 10796 19292 10824 19332
rect 11238 19320 11244 19372
rect 11296 19360 11302 19372
rect 14384 19369 14412 19400
rect 15378 19388 15384 19440
rect 15436 19428 15442 19440
rect 15758 19431 15816 19437
rect 15758 19428 15770 19431
rect 15436 19400 15770 19428
rect 15436 19388 15442 19400
rect 15758 19397 15770 19400
rect 15804 19397 15816 19431
rect 15758 19391 15816 19397
rect 17304 19431 17362 19437
rect 17304 19397 17316 19431
rect 17350 19428 17362 19431
rect 20622 19428 20628 19440
rect 17350 19400 20024 19428
rect 17350 19397 17362 19400
rect 17304 19391 17362 19397
rect 14102 19363 14160 19369
rect 14102 19360 14114 19363
rect 11296 19332 14114 19360
rect 11296 19320 11302 19332
rect 14102 19329 14114 19332
rect 14148 19329 14160 19363
rect 14102 19323 14160 19329
rect 14369 19363 14427 19369
rect 14369 19329 14381 19363
rect 14415 19360 14427 19363
rect 15470 19360 15476 19372
rect 14415 19332 15476 19360
rect 14415 19329 14427 19332
rect 14369 19323 14427 19329
rect 15470 19320 15476 19332
rect 15528 19360 15534 19372
rect 15528 19332 16068 19360
rect 15528 19320 15534 19332
rect 16040 19304 16068 19332
rect 18322 19320 18328 19372
rect 18380 19360 18386 19372
rect 18690 19360 18696 19372
rect 18380 19332 18696 19360
rect 18380 19320 18386 19332
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 19794 19320 19800 19372
rect 19852 19369 19858 19372
rect 19852 19360 19864 19369
rect 19852 19332 19897 19360
rect 19852 19323 19864 19332
rect 19852 19320 19858 19323
rect 11698 19292 11704 19304
rect 10796 19264 11704 19292
rect 9769 19255 9827 19261
rect 11698 19252 11704 19264
rect 11756 19252 11762 19304
rect 16022 19252 16028 19304
rect 16080 19292 16086 19304
rect 17037 19295 17095 19301
rect 17037 19292 17049 19295
rect 16080 19264 17049 19292
rect 16080 19252 16086 19264
rect 8018 19224 8024 19236
rect 5920 19196 8024 19224
rect 8018 19184 8024 19196
rect 8076 19184 8082 19236
rect 10962 19184 10968 19236
rect 11020 19224 11026 19236
rect 11517 19227 11575 19233
rect 11517 19224 11529 19227
rect 11020 19196 11529 19224
rect 11020 19184 11026 19196
rect 11517 19193 11529 19196
rect 11563 19193 11575 19227
rect 12434 19224 12440 19236
rect 11517 19187 11575 19193
rect 11624 19196 12440 19224
rect 5258 19156 5264 19168
rect 5219 19128 5264 19156
rect 5258 19116 5264 19128
rect 5316 19116 5322 19168
rect 7282 19116 7288 19168
rect 7340 19156 7346 19168
rect 11624 19156 11652 19196
rect 12434 19184 12440 19196
rect 12492 19184 12498 19236
rect 11882 19156 11888 19168
rect 7340 19128 11652 19156
rect 11843 19128 11888 19156
rect 7340 19116 7346 19128
rect 11882 19116 11888 19128
rect 11940 19116 11946 19168
rect 12618 19116 12624 19168
rect 12676 19156 12682 19168
rect 15838 19156 15844 19168
rect 12676 19128 15844 19156
rect 12676 19116 12682 19128
rect 15838 19116 15844 19128
rect 15896 19116 15902 19168
rect 16546 19156 16574 19264
rect 17037 19261 17049 19264
rect 17083 19261 17095 19295
rect 19996 19292 20024 19400
rect 20088 19400 20628 19428
rect 20088 19369 20116 19400
rect 20622 19388 20628 19400
rect 20680 19428 20686 19440
rect 21177 19431 21235 19437
rect 21177 19428 21189 19431
rect 20680 19400 21189 19428
rect 20680 19388 20686 19400
rect 21177 19397 21189 19400
rect 21223 19428 21235 19431
rect 21358 19428 21364 19440
rect 21223 19400 21364 19428
rect 21223 19397 21235 19400
rect 21177 19391 21235 19397
rect 21358 19388 21364 19400
rect 21416 19388 21422 19440
rect 20073 19363 20131 19369
rect 20073 19329 20085 19363
rect 20119 19329 20131 19363
rect 20530 19360 20536 19372
rect 20491 19332 20536 19360
rect 20073 19323 20131 19329
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 20254 19292 20260 19304
rect 19996 19264 20260 19292
rect 17037 19255 17095 19261
rect 20254 19252 20260 19264
rect 20312 19252 20318 19304
rect 19058 19224 19064 19236
rect 17972 19196 19064 19224
rect 16669 19159 16727 19165
rect 16669 19156 16681 19159
rect 16546 19128 16681 19156
rect 16669 19125 16681 19128
rect 16715 19125 16727 19159
rect 16669 19119 16727 19125
rect 17034 19116 17040 19168
rect 17092 19156 17098 19168
rect 17972 19156 18000 19196
rect 19058 19184 19064 19196
rect 19116 19184 19122 19236
rect 17092 19128 18000 19156
rect 18417 19159 18475 19165
rect 17092 19116 17098 19128
rect 18417 19125 18429 19159
rect 18463 19156 18475 19159
rect 20346 19156 20352 19168
rect 18463 19128 20352 19156
rect 18463 19125 18475 19128
rect 18417 19119 18475 19125
rect 20346 19116 20352 19128
rect 20404 19116 20410 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 8386 18912 8392 18964
rect 8444 18952 8450 18964
rect 14734 18952 14740 18964
rect 8444 18924 14740 18952
rect 8444 18912 8450 18924
rect 14734 18912 14740 18924
rect 14792 18912 14798 18964
rect 15930 18912 15936 18964
rect 15988 18952 15994 18964
rect 18690 18952 18696 18964
rect 15988 18924 18276 18952
rect 18651 18924 18696 18952
rect 15988 18912 15994 18924
rect 1486 18844 1492 18896
rect 1544 18884 1550 18896
rect 3326 18884 3332 18896
rect 1544 18856 3332 18884
rect 1544 18844 1550 18856
rect 3326 18844 3332 18856
rect 3384 18844 3390 18896
rect 8588 18856 9260 18884
rect 6733 18819 6791 18825
rect 6733 18785 6745 18819
rect 6779 18816 6791 18819
rect 7190 18816 7196 18828
rect 6779 18788 7196 18816
rect 6779 18785 6791 18788
rect 6733 18779 6791 18785
rect 7190 18776 7196 18788
rect 7248 18776 7254 18828
rect 934 18708 940 18760
rect 992 18748 998 18760
rect 4430 18748 4436 18760
rect 992 18720 4436 18748
rect 992 18708 998 18720
rect 4430 18708 4436 18720
rect 4488 18708 4494 18760
rect 6822 18708 6828 18760
rect 6880 18748 6886 18760
rect 8588 18757 8616 18856
rect 6917 18751 6975 18757
rect 6917 18748 6929 18751
rect 6880 18720 6929 18748
rect 6880 18708 6886 18720
rect 6917 18717 6929 18720
rect 6963 18717 6975 18751
rect 6917 18711 6975 18717
rect 8573 18751 8631 18757
rect 8573 18717 8585 18751
rect 8619 18717 8631 18751
rect 9232 18748 9260 18856
rect 10594 18844 10600 18896
rect 10652 18884 10658 18896
rect 11425 18887 11483 18893
rect 11425 18884 11437 18887
rect 10652 18856 11437 18884
rect 10652 18844 10658 18856
rect 11425 18853 11437 18856
rect 11471 18853 11483 18887
rect 11425 18847 11483 18853
rect 16485 18887 16543 18893
rect 16485 18853 16497 18887
rect 16531 18853 16543 18887
rect 18248 18884 18276 18924
rect 18690 18912 18696 18924
rect 18748 18912 18754 18964
rect 22462 18952 22468 18964
rect 19628 18924 22468 18952
rect 19518 18884 19524 18896
rect 18248 18856 19524 18884
rect 16485 18847 16543 18853
rect 9674 18748 9680 18760
rect 9232 18720 9680 18748
rect 8573 18711 8631 18717
rect 9674 18708 9680 18720
rect 9732 18748 9738 18760
rect 10318 18748 10324 18760
rect 9732 18720 10324 18748
rect 9732 18708 9738 18720
rect 10318 18708 10324 18720
rect 10376 18748 10382 18760
rect 12805 18751 12863 18757
rect 12805 18748 12817 18751
rect 10376 18720 12817 18748
rect 10376 18708 10382 18720
rect 8110 18640 8116 18692
rect 8168 18680 8174 18692
rect 8328 18683 8386 18689
rect 8328 18680 8340 18683
rect 8168 18652 8340 18680
rect 8168 18640 8174 18652
rect 8328 18649 8340 18652
rect 8374 18680 8386 18683
rect 8374 18652 8984 18680
rect 8374 18649 8386 18652
rect 8328 18643 8386 18649
rect 5626 18572 5632 18624
rect 5684 18612 5690 18624
rect 5721 18615 5779 18621
rect 5721 18612 5733 18615
rect 5684 18584 5733 18612
rect 5684 18572 5690 18584
rect 5721 18581 5733 18584
rect 5767 18581 5779 18615
rect 5721 18575 5779 18581
rect 5994 18572 6000 18624
rect 6052 18612 6058 18624
rect 6089 18615 6147 18621
rect 6089 18612 6101 18615
rect 6052 18584 6101 18612
rect 6052 18572 6058 18584
rect 6089 18581 6101 18584
rect 6135 18581 6147 18615
rect 6089 18575 6147 18581
rect 7193 18615 7251 18621
rect 7193 18581 7205 18615
rect 7239 18612 7251 18615
rect 7374 18612 7380 18624
rect 7239 18584 7380 18612
rect 7239 18581 7251 18584
rect 7193 18575 7251 18581
rect 7374 18572 7380 18584
rect 7432 18572 7438 18624
rect 8956 18621 8984 18652
rect 9858 18640 9864 18692
rect 9916 18680 9922 18692
rect 10054 18683 10112 18689
rect 10054 18680 10066 18683
rect 9916 18652 10066 18680
rect 9916 18640 9922 18652
rect 10054 18649 10066 18652
rect 10100 18680 10112 18683
rect 10594 18680 10600 18692
rect 10100 18652 10600 18680
rect 10100 18649 10112 18652
rect 10054 18643 10112 18649
rect 10594 18640 10600 18652
rect 10652 18640 10658 18692
rect 10704 18624 10732 18720
rect 12805 18717 12817 18720
rect 12851 18748 12863 18751
rect 13173 18751 13231 18757
rect 13173 18748 13185 18751
rect 12851 18720 13185 18748
rect 12851 18717 12863 18720
rect 12805 18711 12863 18717
rect 13173 18717 13185 18720
rect 13219 18748 13231 18751
rect 13725 18751 13783 18757
rect 13725 18748 13737 18751
rect 13219 18720 13737 18748
rect 13219 18717 13231 18720
rect 13173 18711 13231 18717
rect 13725 18717 13737 18720
rect 13771 18748 13783 18751
rect 14182 18748 14188 18760
rect 13771 18720 14188 18748
rect 13771 18717 13783 18720
rect 13725 18711 13783 18717
rect 14182 18708 14188 18720
rect 14240 18748 14246 18760
rect 14461 18751 14519 18757
rect 14461 18748 14473 18751
rect 14240 18720 14473 18748
rect 14240 18708 14246 18720
rect 14461 18717 14473 18720
rect 14507 18748 14519 18751
rect 16022 18748 16028 18760
rect 14507 18720 16028 18748
rect 14507 18717 14519 18720
rect 14461 18711 14519 18717
rect 16022 18708 16028 18720
rect 16080 18708 16086 18760
rect 16298 18748 16304 18760
rect 16259 18720 16304 18748
rect 16298 18708 16304 18720
rect 16356 18708 16362 18760
rect 16500 18748 16528 18847
rect 19518 18844 19524 18856
rect 19576 18844 19582 18896
rect 19628 18816 19656 18924
rect 22462 18912 22468 18924
rect 22520 18912 22526 18964
rect 20622 18816 20628 18828
rect 18156 18788 19656 18816
rect 20583 18788 20628 18816
rect 18156 18748 18184 18788
rect 20622 18776 20628 18788
rect 20680 18776 20686 18828
rect 16500 18720 18184 18748
rect 18233 18751 18291 18757
rect 18233 18717 18245 18751
rect 18279 18748 18291 18751
rect 18690 18748 18696 18760
rect 18279 18720 18696 18748
rect 18279 18717 18291 18720
rect 18233 18711 18291 18717
rect 18690 18708 18696 18720
rect 18748 18708 18754 18760
rect 18874 18748 18880 18760
rect 18835 18720 18880 18748
rect 18874 18708 18880 18720
rect 18932 18708 18938 18760
rect 20346 18708 20352 18760
rect 20404 18757 20410 18760
rect 20404 18748 20416 18757
rect 20404 18720 20449 18748
rect 20404 18711 20416 18720
rect 20404 18708 20410 18711
rect 20714 18708 20720 18760
rect 20772 18748 20778 18760
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 20772 18720 20913 18748
rect 20772 18708 20778 18720
rect 20901 18717 20913 18720
rect 20947 18717 20959 18751
rect 20901 18711 20959 18717
rect 12066 18640 12072 18692
rect 12124 18680 12130 18692
rect 12560 18683 12618 18689
rect 12560 18680 12572 18683
rect 12124 18652 12572 18680
rect 12124 18640 12130 18652
rect 12560 18649 12572 18652
rect 12606 18680 12618 18683
rect 12606 18652 12848 18680
rect 12606 18649 12618 18652
rect 12560 18643 12618 18649
rect 12820 18624 12848 18652
rect 13262 18640 13268 18692
rect 13320 18680 13326 18692
rect 14706 18683 14764 18689
rect 14706 18680 14718 18683
rect 13320 18652 14718 18680
rect 13320 18640 13326 18652
rect 14706 18649 14718 18652
rect 14752 18649 14764 18683
rect 16482 18680 16488 18692
rect 14706 18643 14764 18649
rect 14844 18652 16488 18680
rect 8941 18615 8999 18621
rect 8941 18581 8953 18615
rect 8987 18581 8999 18615
rect 8941 18575 8999 18581
rect 9030 18572 9036 18624
rect 9088 18612 9094 18624
rect 10502 18612 10508 18624
rect 9088 18584 10508 18612
rect 9088 18572 9094 18584
rect 10502 18572 10508 18584
rect 10560 18572 10566 18624
rect 10686 18612 10692 18624
rect 10647 18584 10692 18612
rect 10686 18572 10692 18584
rect 10744 18612 10750 18624
rect 10962 18612 10968 18624
rect 10744 18584 10968 18612
rect 10744 18572 10750 18584
rect 10962 18572 10968 18584
rect 11020 18572 11026 18624
rect 11054 18572 11060 18624
rect 11112 18612 11118 18624
rect 12710 18612 12716 18624
rect 11112 18584 12716 18612
rect 11112 18572 11118 18584
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 12802 18572 12808 18624
rect 12860 18572 12866 18624
rect 14458 18572 14464 18624
rect 14516 18612 14522 18624
rect 14844 18612 14872 18652
rect 16482 18640 16488 18652
rect 16540 18640 16546 18692
rect 16666 18640 16672 18692
rect 16724 18680 16730 18692
rect 17988 18683 18046 18689
rect 17988 18680 18000 18683
rect 16724 18652 18000 18680
rect 16724 18640 16730 18652
rect 17988 18649 18000 18652
rect 18034 18680 18046 18683
rect 19978 18680 19984 18692
rect 18034 18652 19984 18680
rect 18034 18649 18046 18652
rect 17988 18643 18046 18649
rect 19978 18640 19984 18652
rect 20036 18640 20042 18692
rect 21174 18680 21180 18692
rect 21135 18652 21180 18680
rect 21174 18640 21180 18652
rect 21232 18640 21238 18692
rect 15838 18612 15844 18624
rect 14516 18584 14872 18612
rect 15799 18584 15844 18612
rect 14516 18572 14522 18584
rect 15838 18572 15844 18584
rect 15896 18572 15902 18624
rect 16853 18615 16911 18621
rect 16853 18581 16865 18615
rect 16899 18612 16911 18615
rect 17126 18612 17132 18624
rect 16899 18584 17132 18612
rect 16899 18581 16911 18584
rect 16853 18575 16911 18581
rect 17126 18572 17132 18584
rect 17184 18612 17190 18624
rect 17678 18612 17684 18624
rect 17184 18584 17684 18612
rect 17184 18572 17190 18584
rect 17678 18572 17684 18584
rect 17736 18572 17742 18624
rect 19245 18615 19303 18621
rect 19245 18581 19257 18615
rect 19291 18612 19303 18615
rect 19794 18612 19800 18624
rect 19291 18584 19800 18612
rect 19291 18581 19303 18584
rect 19245 18575 19303 18581
rect 19794 18572 19800 18584
rect 19852 18612 19858 18624
rect 20070 18612 20076 18624
rect 19852 18584 20076 18612
rect 19852 18572 19858 18584
rect 20070 18572 20076 18584
rect 20128 18572 20134 18624
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 6730 18408 6736 18420
rect 6691 18380 6736 18408
rect 6730 18368 6736 18380
rect 6788 18368 6794 18420
rect 7837 18411 7895 18417
rect 7837 18377 7849 18411
rect 7883 18408 7895 18411
rect 8573 18411 8631 18417
rect 8573 18408 8585 18411
rect 7883 18380 8585 18408
rect 7883 18377 7895 18380
rect 7837 18371 7895 18377
rect 8573 18377 8585 18380
rect 8619 18408 8631 18411
rect 9214 18408 9220 18420
rect 8619 18380 9220 18408
rect 8619 18377 8631 18380
rect 8573 18371 8631 18377
rect 9214 18368 9220 18380
rect 9272 18368 9278 18420
rect 14274 18408 14280 18420
rect 9324 18380 14280 18408
rect 6914 18300 6920 18352
rect 6972 18340 6978 18352
rect 9324 18340 9352 18380
rect 14274 18368 14280 18380
rect 14332 18368 14338 18420
rect 16022 18408 16028 18420
rect 15983 18380 16028 18408
rect 16022 18368 16028 18380
rect 16080 18368 16086 18420
rect 18782 18408 18788 18420
rect 16546 18380 18788 18408
rect 11146 18340 11152 18352
rect 6972 18312 9352 18340
rect 9407 18312 11152 18340
rect 6972 18300 6978 18312
rect 6638 18232 6644 18284
rect 6696 18272 6702 18284
rect 7101 18275 7159 18281
rect 7101 18272 7113 18275
rect 6696 18244 7113 18272
rect 6696 18232 6702 18244
rect 7101 18241 7113 18244
rect 7147 18272 7159 18275
rect 7929 18275 7987 18281
rect 7929 18272 7941 18275
rect 7147 18244 7941 18272
rect 7147 18241 7159 18244
rect 7101 18235 7159 18241
rect 7929 18241 7941 18244
rect 7975 18241 7987 18275
rect 7929 18235 7987 18241
rect 2590 18096 2596 18148
rect 2648 18136 2654 18148
rect 4890 18136 4896 18148
rect 2648 18108 4896 18136
rect 2648 18096 2654 18108
rect 4890 18096 4896 18108
rect 4948 18096 4954 18148
rect 3142 18028 3148 18080
rect 3200 18068 3206 18080
rect 5442 18068 5448 18080
rect 3200 18040 5448 18068
rect 3200 18028 3206 18040
rect 5442 18028 5448 18040
rect 5500 18028 5506 18080
rect 7466 18068 7472 18080
rect 7427 18040 7472 18068
rect 7466 18028 7472 18040
rect 7524 18028 7530 18080
rect 7944 18068 7972 18235
rect 8110 18204 8116 18216
rect 8071 18176 8116 18204
rect 8110 18164 8116 18176
rect 8168 18164 8174 18216
rect 8018 18096 8024 18148
rect 8076 18136 8082 18148
rect 9033 18139 9091 18145
rect 9033 18136 9045 18139
rect 8076 18108 9045 18136
rect 8076 18096 8082 18108
rect 9033 18105 9045 18108
rect 9079 18136 9091 18139
rect 9407 18136 9435 18312
rect 11146 18300 11152 18312
rect 11204 18300 11210 18352
rect 12250 18300 12256 18352
rect 12308 18340 12314 18352
rect 13642 18343 13700 18349
rect 13642 18340 13654 18343
rect 12308 18312 13654 18340
rect 12308 18300 12314 18312
rect 13642 18309 13654 18312
rect 13688 18309 13700 18343
rect 13642 18303 13700 18309
rect 13814 18300 13820 18352
rect 13872 18340 13878 18352
rect 14522 18343 14580 18349
rect 14522 18340 14534 18343
rect 13872 18312 14534 18340
rect 13872 18300 13878 18312
rect 14522 18309 14534 18312
rect 14568 18309 14580 18343
rect 16546 18340 16574 18380
rect 18782 18368 18788 18380
rect 18840 18368 18846 18420
rect 19702 18408 19708 18420
rect 19663 18380 19708 18408
rect 19702 18368 19708 18380
rect 19760 18368 19766 18420
rect 18690 18340 18696 18352
rect 14522 18303 14580 18309
rect 15764 18312 16574 18340
rect 18340 18312 18696 18340
rect 9674 18232 9680 18284
rect 9732 18272 9738 18284
rect 9858 18272 9864 18284
rect 9732 18244 9864 18272
rect 9732 18232 9738 18244
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 10134 18232 10140 18284
rect 10192 18281 10198 18284
rect 10192 18272 10204 18281
rect 10192 18244 10237 18272
rect 10192 18235 10204 18244
rect 10192 18232 10198 18235
rect 10318 18232 10324 18284
rect 10376 18272 10382 18284
rect 10413 18275 10471 18281
rect 10413 18272 10425 18275
rect 10376 18244 10425 18272
rect 10376 18232 10382 18244
rect 10413 18241 10425 18244
rect 10459 18241 10471 18275
rect 10413 18235 10471 18241
rect 11330 18232 11336 18284
rect 11388 18272 11394 18284
rect 11882 18272 11888 18284
rect 11388 18244 11888 18272
rect 11388 18232 11394 18244
rect 11882 18232 11888 18244
rect 11940 18272 11946 18284
rect 13909 18275 13967 18281
rect 11940 18244 13860 18272
rect 11940 18232 11946 18244
rect 12618 18204 12624 18216
rect 9079 18108 9435 18136
rect 10520 18176 12624 18204
rect 9079 18105 9091 18108
rect 9033 18099 9091 18105
rect 10520 18068 10548 18176
rect 12618 18164 12624 18176
rect 12676 18164 12682 18216
rect 13832 18204 13860 18244
rect 13909 18241 13921 18275
rect 13955 18272 13967 18275
rect 14182 18272 14188 18284
rect 13955 18244 14188 18272
rect 13955 18241 13967 18244
rect 13909 18235 13967 18241
rect 14182 18232 14188 18244
rect 14240 18272 14246 18284
rect 14277 18275 14335 18281
rect 14277 18272 14289 18275
rect 14240 18244 14289 18272
rect 14240 18232 14246 18244
rect 14277 18241 14289 18244
rect 14323 18241 14335 18275
rect 15764 18272 15792 18312
rect 14277 18235 14335 18241
rect 14384 18244 15792 18272
rect 14384 18204 14412 18244
rect 15838 18232 15844 18284
rect 15896 18272 15902 18284
rect 18340 18281 18368 18312
rect 18690 18300 18696 18312
rect 18748 18340 18754 18352
rect 20622 18340 20628 18352
rect 18748 18312 20628 18340
rect 18748 18300 18754 18312
rect 19996 18281 20024 18312
rect 20622 18300 20628 18312
rect 20680 18300 20686 18352
rect 16925 18275 16983 18281
rect 16925 18272 16937 18275
rect 15896 18244 16937 18272
rect 15896 18232 15902 18244
rect 16925 18241 16937 18244
rect 16971 18241 16983 18275
rect 16925 18235 16983 18241
rect 18325 18275 18383 18281
rect 18325 18241 18337 18275
rect 18371 18241 18383 18275
rect 18581 18275 18639 18281
rect 18581 18272 18593 18275
rect 18325 18235 18383 18241
rect 18432 18244 18593 18272
rect 13832 18176 14412 18204
rect 16022 18164 16028 18216
rect 16080 18204 16086 18216
rect 16482 18204 16488 18216
rect 16080 18176 16488 18204
rect 16080 18164 16086 18176
rect 16482 18164 16488 18176
rect 16540 18204 16546 18216
rect 16669 18207 16727 18213
rect 16669 18204 16681 18207
rect 16540 18176 16681 18204
rect 16540 18164 16546 18176
rect 16669 18173 16681 18176
rect 16715 18173 16727 18207
rect 16669 18167 16727 18173
rect 18138 18164 18144 18216
rect 18196 18204 18202 18216
rect 18432 18204 18460 18244
rect 18581 18241 18593 18244
rect 18627 18241 18639 18275
rect 18581 18235 18639 18241
rect 19981 18275 20039 18281
rect 19981 18241 19993 18275
rect 20027 18241 20039 18275
rect 20237 18275 20295 18281
rect 20237 18272 20249 18275
rect 19981 18235 20039 18241
rect 20088 18244 20249 18272
rect 20088 18204 20116 18244
rect 20237 18241 20249 18244
rect 20283 18241 20295 18275
rect 20237 18235 20295 18241
rect 18196 18176 18460 18204
rect 19352 18176 20116 18204
rect 18196 18164 18202 18176
rect 11698 18096 11704 18148
rect 11756 18136 11762 18148
rect 12529 18139 12587 18145
rect 12529 18136 12541 18139
rect 11756 18108 12541 18136
rect 11756 18096 11762 18108
rect 12529 18105 12541 18108
rect 12575 18105 12587 18139
rect 16298 18136 16304 18148
rect 12529 18099 12587 18105
rect 15580 18108 16304 18136
rect 10686 18068 10692 18080
rect 7944 18040 10548 18068
rect 10647 18040 10692 18068
rect 10686 18028 10692 18040
rect 10744 18068 10750 18080
rect 11057 18071 11115 18077
rect 11057 18068 11069 18071
rect 10744 18040 11069 18068
rect 10744 18028 10750 18040
rect 11057 18037 11069 18040
rect 11103 18068 11115 18071
rect 11793 18071 11851 18077
rect 11793 18068 11805 18071
rect 11103 18040 11805 18068
rect 11103 18037 11115 18040
rect 11057 18031 11115 18037
rect 11793 18037 11805 18040
rect 11839 18068 11851 18071
rect 12161 18071 12219 18077
rect 12161 18068 12173 18071
rect 11839 18040 12173 18068
rect 11839 18037 11851 18040
rect 11793 18031 11851 18037
rect 12161 18037 12173 18040
rect 12207 18037 12219 18071
rect 12161 18031 12219 18037
rect 13538 18028 13544 18080
rect 13596 18068 13602 18080
rect 15580 18068 15608 18108
rect 16298 18096 16304 18108
rect 16356 18096 16362 18148
rect 17678 18096 17684 18148
rect 17736 18136 17742 18148
rect 17736 18108 18184 18136
rect 17736 18096 17742 18108
rect 13596 18040 15608 18068
rect 15657 18071 15715 18077
rect 13596 18028 13602 18040
rect 15657 18037 15669 18071
rect 15703 18068 15715 18071
rect 17034 18068 17040 18080
rect 15703 18040 17040 18068
rect 15703 18037 15715 18040
rect 15657 18031 15715 18037
rect 17034 18028 17040 18040
rect 17092 18028 17098 18080
rect 18046 18068 18052 18080
rect 18007 18040 18052 18068
rect 18046 18028 18052 18040
rect 18104 18028 18110 18080
rect 18156 18068 18184 18108
rect 19352 18068 19380 18176
rect 18156 18040 19380 18068
rect 21361 18071 21419 18077
rect 21361 18037 21373 18071
rect 21407 18068 21419 18071
rect 21450 18068 21456 18080
rect 21407 18040 21456 18068
rect 21407 18037 21419 18040
rect 21361 18031 21419 18037
rect 21450 18028 21456 18040
rect 21508 18028 21514 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 9766 17824 9772 17876
rect 9824 17864 9830 17876
rect 13173 17867 13231 17873
rect 13173 17864 13185 17867
rect 9824 17836 13185 17864
rect 9824 17824 9830 17836
rect 13173 17833 13185 17836
rect 13219 17833 13231 17867
rect 13173 17827 13231 17833
rect 7098 17688 7104 17740
rect 7156 17728 7162 17740
rect 7193 17731 7251 17737
rect 7193 17728 7205 17731
rect 7156 17700 7205 17728
rect 7156 17688 7162 17700
rect 7193 17697 7205 17700
rect 7239 17697 7251 17731
rect 7193 17691 7251 17697
rect 7374 17688 7380 17740
rect 7432 17728 7438 17740
rect 11698 17728 11704 17740
rect 7432 17700 9904 17728
rect 7432 17688 7438 17700
rect 7469 17663 7527 17669
rect 7469 17629 7481 17663
rect 7515 17660 7527 17663
rect 7650 17660 7656 17672
rect 7515 17632 7656 17660
rect 7515 17629 7527 17632
rect 7469 17623 7527 17629
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 9033 17663 9091 17669
rect 9033 17629 9045 17663
rect 9079 17660 9091 17663
rect 9122 17660 9128 17672
rect 9079 17632 9128 17660
rect 9079 17629 9091 17632
rect 9033 17623 9091 17629
rect 9122 17620 9128 17632
rect 9180 17660 9186 17672
rect 9769 17663 9827 17669
rect 9769 17660 9781 17663
rect 9180 17632 9781 17660
rect 9180 17620 9186 17632
rect 9769 17629 9781 17632
rect 9815 17629 9827 17663
rect 9876 17660 9904 17700
rect 11348 17700 11704 17728
rect 10025 17663 10083 17669
rect 10025 17660 10037 17663
rect 9876 17632 10037 17660
rect 9769 17623 9827 17629
rect 10025 17629 10037 17632
rect 10071 17629 10083 17663
rect 11348 17660 11376 17700
rect 11698 17688 11704 17700
rect 11756 17688 11762 17740
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 10025 17623 10083 17629
rect 10704 17632 11376 17660
rect 11440 17632 11805 17660
rect 4062 17552 4068 17604
rect 4120 17592 4126 17604
rect 10704 17592 10732 17632
rect 4120 17564 10732 17592
rect 4120 17552 4126 17564
rect 6730 17484 6736 17536
rect 6788 17524 6794 17536
rect 10962 17524 10968 17536
rect 6788 17496 10968 17524
rect 6788 17484 6794 17496
rect 10962 17484 10968 17496
rect 11020 17484 11026 17536
rect 11146 17524 11152 17536
rect 11107 17496 11152 17524
rect 11146 17484 11152 17496
rect 11204 17484 11210 17536
rect 11238 17484 11244 17536
rect 11296 17524 11302 17536
rect 11440 17533 11468 17632
rect 11793 17629 11805 17632
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 11882 17552 11888 17604
rect 11940 17592 11946 17604
rect 12038 17595 12096 17601
rect 12038 17592 12050 17595
rect 11940 17564 12050 17592
rect 11940 17552 11946 17564
rect 12038 17561 12050 17564
rect 12084 17561 12096 17595
rect 13188 17592 13216 17827
rect 16022 17824 16028 17876
rect 16080 17864 16086 17876
rect 17129 17867 17187 17873
rect 17129 17864 17141 17867
rect 16080 17836 17141 17864
rect 16080 17824 16086 17836
rect 17129 17833 17141 17836
rect 17175 17833 17187 17867
rect 17129 17827 17187 17833
rect 18138 17824 18144 17876
rect 18196 17864 18202 17876
rect 19981 17867 20039 17873
rect 19981 17864 19993 17867
rect 18196 17836 19993 17864
rect 18196 17824 18202 17836
rect 19981 17833 19993 17836
rect 20027 17833 20039 17867
rect 19981 17827 20039 17833
rect 19610 17796 19616 17808
rect 19571 17768 19616 17796
rect 19610 17756 19616 17768
rect 19668 17756 19674 17808
rect 13541 17663 13599 17669
rect 13541 17629 13553 17663
rect 13587 17660 13599 17663
rect 14185 17663 14243 17669
rect 14185 17660 14197 17663
rect 13587 17632 14197 17660
rect 13587 17629 13599 17632
rect 13541 17623 13599 17629
rect 14185 17629 14197 17632
rect 14231 17660 14243 17663
rect 14829 17663 14887 17669
rect 14829 17660 14841 17663
rect 14231 17632 14841 17660
rect 14231 17629 14243 17632
rect 14185 17623 14243 17629
rect 14829 17629 14841 17632
rect 14875 17660 14887 17663
rect 15105 17663 15163 17669
rect 15105 17660 15117 17663
rect 14875 17632 15117 17660
rect 14875 17629 14887 17632
rect 14829 17623 14887 17629
rect 15105 17629 15117 17632
rect 15151 17660 15163 17663
rect 16482 17660 16488 17672
rect 15151 17632 16488 17660
rect 15151 17629 15163 17632
rect 15105 17623 15163 17629
rect 16482 17620 16488 17632
rect 16540 17660 16546 17672
rect 16853 17663 16911 17669
rect 16853 17660 16865 17663
rect 16540 17632 16865 17660
rect 16540 17620 16546 17632
rect 16853 17629 16865 17632
rect 16899 17660 16911 17663
rect 18509 17663 18567 17669
rect 18509 17660 18521 17663
rect 16899 17632 18521 17660
rect 16899 17629 16911 17632
rect 16853 17623 16911 17629
rect 18509 17629 18521 17632
rect 18555 17629 18567 17663
rect 18509 17623 18567 17629
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17660 19487 17663
rect 19518 17660 19524 17672
rect 19475 17632 19524 17660
rect 19475 17629 19487 17632
rect 19429 17623 19487 17629
rect 19518 17620 19524 17632
rect 19576 17620 19582 17672
rect 20622 17620 20628 17672
rect 20680 17660 20686 17672
rect 21361 17663 21419 17669
rect 21361 17660 21373 17663
rect 20680 17632 21373 17660
rect 20680 17620 20686 17632
rect 21361 17629 21373 17632
rect 21407 17629 21419 17663
rect 21361 17623 21419 17629
rect 15350 17595 15408 17601
rect 15350 17592 15362 17595
rect 13188 17564 15362 17592
rect 12038 17555 12096 17561
rect 15350 17561 15362 17564
rect 15396 17561 15408 17595
rect 15350 17555 15408 17561
rect 18046 17552 18052 17604
rect 18104 17592 18110 17604
rect 18242 17595 18300 17601
rect 18242 17592 18254 17595
rect 18104 17564 18254 17592
rect 18104 17552 18110 17564
rect 18242 17561 18254 17564
rect 18288 17561 18300 17595
rect 18242 17555 18300 17561
rect 18598 17552 18604 17604
rect 18656 17592 18662 17604
rect 21116 17595 21174 17601
rect 18656 17564 18920 17592
rect 18656 17552 18662 17564
rect 11425 17527 11483 17533
rect 11425 17524 11437 17527
rect 11296 17496 11437 17524
rect 11296 17484 11302 17496
rect 11425 17493 11437 17496
rect 11471 17493 11483 17527
rect 11425 17487 11483 17493
rect 15102 17484 15108 17536
rect 15160 17524 15166 17536
rect 16485 17527 16543 17533
rect 16485 17524 16497 17527
rect 15160 17496 16497 17524
rect 15160 17484 15166 17496
rect 16485 17493 16497 17496
rect 16531 17493 16543 17527
rect 18782 17524 18788 17536
rect 18743 17496 18788 17524
rect 16485 17487 16543 17493
rect 18782 17484 18788 17496
rect 18840 17484 18846 17536
rect 18892 17524 18920 17564
rect 21116 17561 21128 17595
rect 21162 17592 21174 17595
rect 21450 17592 21456 17604
rect 21162 17564 21456 17592
rect 21162 17561 21174 17564
rect 21116 17555 21174 17561
rect 21450 17552 21456 17564
rect 21508 17552 21514 17604
rect 21542 17524 21548 17536
rect 18892 17496 21548 17524
rect 21542 17484 21548 17496
rect 21600 17484 21606 17536
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 4246 17280 4252 17332
rect 4304 17320 4310 17332
rect 4525 17323 4583 17329
rect 4525 17320 4537 17323
rect 4304 17292 4537 17320
rect 4304 17280 4310 17292
rect 4525 17289 4537 17292
rect 4571 17289 4583 17323
rect 4890 17320 4896 17332
rect 4851 17292 4896 17320
rect 4525 17283 4583 17289
rect 4540 17252 4568 17283
rect 4890 17280 4896 17292
rect 4948 17320 4954 17332
rect 5537 17323 5595 17329
rect 5537 17320 5549 17323
rect 4948 17292 5549 17320
rect 4948 17280 4954 17292
rect 5537 17289 5549 17292
rect 5583 17289 5595 17323
rect 7650 17320 7656 17332
rect 7611 17292 7656 17320
rect 5537 17283 5595 17289
rect 7650 17280 7656 17292
rect 7708 17280 7714 17332
rect 8021 17323 8079 17329
rect 8021 17289 8033 17323
rect 8067 17320 8079 17323
rect 8202 17320 8208 17332
rect 8067 17292 8208 17320
rect 8067 17289 8079 17292
rect 8021 17283 8079 17289
rect 8202 17280 8208 17292
rect 8260 17280 8266 17332
rect 10042 17280 10048 17332
rect 10100 17320 10106 17332
rect 10870 17320 10876 17332
rect 10100 17292 10876 17320
rect 10100 17280 10106 17292
rect 10870 17280 10876 17292
rect 10928 17280 10934 17332
rect 11977 17323 12035 17329
rect 11977 17289 11989 17323
rect 12023 17320 12035 17323
rect 18966 17320 18972 17332
rect 12023 17292 18972 17320
rect 12023 17289 12035 17292
rect 11977 17283 12035 17289
rect 18966 17280 18972 17292
rect 19024 17280 19030 17332
rect 19076 17292 20668 17320
rect 5629 17255 5687 17261
rect 5629 17252 5641 17255
rect 4540 17224 5641 17252
rect 5629 17221 5641 17224
rect 5675 17252 5687 17255
rect 5994 17252 6000 17264
rect 5675 17224 6000 17252
rect 5675 17221 5687 17224
rect 5629 17215 5687 17221
rect 5994 17212 6000 17224
rect 6052 17212 6058 17264
rect 8220 17224 10824 17252
rect 5445 17119 5503 17125
rect 5445 17085 5457 17119
rect 5491 17116 5503 17119
rect 5534 17116 5540 17128
rect 5491 17088 5540 17116
rect 5491 17085 5503 17088
rect 5445 17079 5503 17085
rect 5534 17076 5540 17088
rect 5592 17076 5598 17128
rect 8220 17125 8248 17224
rect 9858 17144 9864 17196
rect 9916 17184 9922 17196
rect 10146 17187 10204 17193
rect 10146 17184 10158 17187
rect 9916 17156 10158 17184
rect 9916 17144 9922 17156
rect 10146 17153 10158 17156
rect 10192 17153 10204 17187
rect 10146 17147 10204 17153
rect 8113 17119 8171 17125
rect 8113 17085 8125 17119
rect 8159 17085 8171 17119
rect 8113 17079 8171 17085
rect 8205 17119 8263 17125
rect 8205 17085 8217 17119
rect 8251 17085 8263 17119
rect 8205 17079 8263 17085
rect 10413 17119 10471 17125
rect 10413 17085 10425 17119
rect 10459 17116 10471 17119
rect 10796 17116 10824 17224
rect 12342 17212 12348 17264
rect 12400 17252 12406 17264
rect 12621 17255 12679 17261
rect 12621 17252 12633 17255
rect 12400 17224 12633 17252
rect 12400 17212 12406 17224
rect 12621 17221 12633 17224
rect 12667 17252 12679 17255
rect 12989 17255 13047 17261
rect 12989 17252 13001 17255
rect 12667 17224 13001 17252
rect 12667 17221 12679 17224
rect 12621 17215 12679 17221
rect 12989 17221 13001 17224
rect 13035 17221 13047 17255
rect 19076 17252 19104 17292
rect 12989 17215 13047 17221
rect 13096 17224 19104 17252
rect 12894 17144 12900 17196
rect 12952 17184 12958 17196
rect 13096 17184 13124 17224
rect 19702 17212 19708 17264
rect 19760 17252 19766 17264
rect 19760 17224 20300 17252
rect 19760 17212 19766 17224
rect 12952 17156 13124 17184
rect 12952 17144 12958 17156
rect 14826 17144 14832 17196
rect 14884 17193 14890 17196
rect 14884 17184 14896 17193
rect 18049 17187 18107 17193
rect 14884 17156 14929 17184
rect 14884 17147 14896 17156
rect 18049 17153 18061 17187
rect 18095 17153 18107 17187
rect 18049 17147 18107 17153
rect 18325 17187 18383 17193
rect 18325 17153 18337 17187
rect 18371 17184 18383 17187
rect 18782 17184 18788 17196
rect 18371 17156 18788 17184
rect 18371 17153 18383 17156
rect 18325 17147 18383 17153
rect 14884 17144 14890 17147
rect 15105 17119 15163 17125
rect 10459 17088 10732 17116
rect 10796 17088 14136 17116
rect 10459 17085 10471 17088
rect 10413 17079 10471 17085
rect 8128 17048 8156 17079
rect 8662 17048 8668 17060
rect 8128 17020 8668 17048
rect 8662 17008 8668 17020
rect 8720 17008 8726 17060
rect 8757 17051 8815 17057
rect 8757 17017 8769 17051
rect 8803 17048 8815 17051
rect 9122 17048 9128 17060
rect 8803 17020 9128 17048
rect 8803 17017 8815 17020
rect 8757 17011 8815 17017
rect 9122 17008 9128 17020
rect 9180 17008 9186 17060
rect 10704 16992 10732 17088
rect 12710 17008 12716 17060
rect 12768 17048 12774 17060
rect 13725 17051 13783 17057
rect 13725 17048 13737 17051
rect 12768 17020 13737 17048
rect 12768 17008 12774 17020
rect 13725 17017 13737 17020
rect 13771 17017 13783 17051
rect 13725 17011 13783 17017
rect 5997 16983 6055 16989
rect 5997 16949 6009 16983
rect 6043 16980 6055 16983
rect 6638 16980 6644 16992
rect 6043 16952 6644 16980
rect 6043 16949 6055 16952
rect 5997 16943 6055 16949
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 9033 16983 9091 16989
rect 9033 16949 9045 16983
rect 9079 16980 9091 16983
rect 10502 16980 10508 16992
rect 9079 16952 10508 16980
rect 9079 16949 9091 16952
rect 9033 16943 9091 16949
rect 10502 16940 10508 16952
rect 10560 16940 10566 16992
rect 10686 16980 10692 16992
rect 10647 16952 10692 16980
rect 10686 16940 10692 16952
rect 10744 16980 10750 16992
rect 11057 16983 11115 16989
rect 11057 16980 11069 16983
rect 10744 16952 11069 16980
rect 10744 16940 10750 16952
rect 11057 16949 11069 16952
rect 11103 16980 11115 16983
rect 11238 16980 11244 16992
rect 11103 16952 11244 16980
rect 11103 16949 11115 16952
rect 11057 16943 11115 16949
rect 11238 16940 11244 16952
rect 11296 16980 11302 16992
rect 11517 16983 11575 16989
rect 11517 16980 11529 16983
rect 11296 16952 11529 16980
rect 11296 16940 11302 16952
rect 11517 16949 11529 16952
rect 11563 16980 11575 16983
rect 12253 16983 12311 16989
rect 12253 16980 12265 16983
rect 11563 16952 12265 16980
rect 11563 16949 11575 16952
rect 11517 16943 11575 16949
rect 12253 16949 12265 16952
rect 12299 16980 12311 16983
rect 12342 16980 12348 16992
rect 12299 16952 12348 16980
rect 12299 16949 12311 16952
rect 12253 16943 12311 16949
rect 12342 16940 12348 16952
rect 12400 16940 12406 16992
rect 13446 16980 13452 16992
rect 13407 16952 13452 16980
rect 13446 16940 13452 16952
rect 13504 16940 13510 16992
rect 14108 16980 14136 17088
rect 15105 17085 15117 17119
rect 15151 17116 15163 17119
rect 15565 17119 15623 17125
rect 15565 17116 15577 17119
rect 15151 17088 15577 17116
rect 15151 17085 15163 17088
rect 15105 17079 15163 17085
rect 15565 17085 15577 17088
rect 15611 17116 15623 17119
rect 15746 17116 15752 17128
rect 15611 17088 15752 17116
rect 15611 17085 15623 17088
rect 15565 17079 15623 17085
rect 15746 17076 15752 17088
rect 15804 17116 15810 17128
rect 15933 17119 15991 17125
rect 15933 17116 15945 17119
rect 15804 17088 15945 17116
rect 15804 17076 15810 17088
rect 15933 17085 15945 17088
rect 15979 17116 15991 17119
rect 18064 17116 18092 17147
rect 18782 17144 18788 17156
rect 18840 17144 18846 17196
rect 19978 17184 19984 17196
rect 20036 17193 20042 17196
rect 19948 17156 19984 17184
rect 19978 17144 19984 17156
rect 20036 17147 20048 17193
rect 20036 17144 20042 17147
rect 20162 17144 20168 17196
rect 20220 17144 20226 17196
rect 20272 17193 20300 17224
rect 20257 17187 20315 17193
rect 20257 17153 20269 17187
rect 20303 17184 20315 17187
rect 20530 17184 20536 17196
rect 20303 17156 20536 17184
rect 20303 17153 20315 17156
rect 20257 17147 20315 17153
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 20640 17193 20668 17292
rect 20625 17187 20683 17193
rect 20625 17153 20637 17187
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 20180 17116 20208 17144
rect 20809 17119 20867 17125
rect 20809 17116 20821 17119
rect 15979 17088 16574 17116
rect 18064 17088 19104 17116
rect 20180 17088 20821 17116
rect 15979 17085 15991 17088
rect 15933 17079 15991 17085
rect 16022 16980 16028 16992
rect 14108 16952 16028 16980
rect 16022 16940 16028 16952
rect 16080 16940 16086 16992
rect 16546 16980 16574 17088
rect 18509 17051 18567 17057
rect 18509 17017 18521 17051
rect 18555 17048 18567 17051
rect 18598 17048 18604 17060
rect 18555 17020 18604 17048
rect 18555 17017 18567 17020
rect 18509 17011 18567 17017
rect 18598 17008 18604 17020
rect 18656 17008 18662 17060
rect 16761 16983 16819 16989
rect 16761 16980 16773 16983
rect 16546 16952 16773 16980
rect 16761 16949 16773 16952
rect 16807 16980 16819 16983
rect 17221 16983 17279 16989
rect 17221 16980 17233 16983
rect 16807 16952 17233 16980
rect 16807 16949 16819 16952
rect 16761 16943 16819 16949
rect 17221 16949 17233 16952
rect 17267 16949 17279 16983
rect 17221 16943 17279 16949
rect 17865 16983 17923 16989
rect 17865 16949 17877 16983
rect 17911 16980 17923 16983
rect 18690 16980 18696 16992
rect 17911 16952 18696 16980
rect 17911 16949 17923 16952
rect 17865 16943 17923 16949
rect 18690 16940 18696 16952
rect 18748 16940 18754 16992
rect 18877 16983 18935 16989
rect 18877 16949 18889 16983
rect 18923 16980 18935 16983
rect 18966 16980 18972 16992
rect 18923 16952 18972 16980
rect 18923 16949 18935 16952
rect 18877 16943 18935 16949
rect 18966 16940 18972 16952
rect 19024 16940 19030 16992
rect 19076 16980 19104 17088
rect 20809 17085 20821 17088
rect 20855 17085 20867 17119
rect 20809 17079 20867 17085
rect 21174 16980 21180 16992
rect 19076 16952 21180 16980
rect 21174 16940 21180 16952
rect 21232 16940 21238 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 8662 16736 8668 16788
rect 8720 16776 8726 16788
rect 11698 16776 11704 16788
rect 8720 16748 11704 16776
rect 8720 16736 8726 16748
rect 11698 16736 11704 16748
rect 11756 16736 11762 16788
rect 12986 16736 12992 16788
rect 13044 16776 13050 16788
rect 13446 16776 13452 16788
rect 13044 16748 13452 16776
rect 13044 16736 13050 16748
rect 13446 16736 13452 16748
rect 13504 16776 13510 16788
rect 19518 16776 19524 16788
rect 13504 16748 19524 16776
rect 13504 16736 13510 16748
rect 19518 16736 19524 16748
rect 19576 16736 19582 16788
rect 17497 16711 17555 16717
rect 17497 16677 17509 16711
rect 17543 16677 17555 16711
rect 17497 16671 17555 16677
rect 12250 16640 12256 16652
rect 11992 16612 12256 16640
rect 8573 16575 8631 16581
rect 8573 16541 8585 16575
rect 8619 16572 8631 16575
rect 9033 16575 9091 16581
rect 9033 16572 9045 16575
rect 8619 16544 9045 16572
rect 8619 16541 8631 16544
rect 8573 16535 8631 16541
rect 9033 16541 9045 16544
rect 9079 16572 9091 16575
rect 9122 16572 9128 16584
rect 9079 16544 9128 16572
rect 9079 16541 9091 16544
rect 9033 16535 9091 16541
rect 9122 16532 9128 16544
rect 9180 16532 9186 16584
rect 10686 16572 10692 16584
rect 10647 16544 10692 16572
rect 10686 16532 10692 16544
rect 10744 16532 10750 16584
rect 11992 16572 12020 16612
rect 12250 16600 12256 16612
rect 12308 16600 12314 16652
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 13372 16612 14105 16640
rect 10897 16544 12020 16572
rect 5534 16464 5540 16516
rect 5592 16504 5598 16516
rect 5592 16476 7236 16504
rect 5592 16464 5598 16476
rect 4154 16396 4160 16448
rect 4212 16436 4218 16448
rect 4525 16439 4583 16445
rect 4525 16436 4537 16439
rect 4212 16408 4537 16436
rect 4212 16396 4218 16408
rect 4525 16405 4537 16408
rect 4571 16405 4583 16439
rect 4525 16399 4583 16405
rect 5902 16396 5908 16448
rect 5960 16436 5966 16448
rect 7208 16445 7236 16476
rect 7558 16464 7564 16516
rect 7616 16504 7622 16516
rect 8306 16507 8364 16513
rect 8306 16504 8318 16507
rect 7616 16476 8318 16504
rect 7616 16464 7622 16476
rect 8306 16473 8318 16476
rect 8352 16473 8364 16507
rect 9278 16507 9336 16513
rect 9278 16504 9290 16507
rect 8306 16467 8364 16473
rect 8404 16476 9290 16504
rect 6457 16439 6515 16445
rect 6457 16436 6469 16439
rect 5960 16408 6469 16436
rect 5960 16396 5966 16408
rect 6457 16405 6469 16408
rect 6503 16405 6515 16439
rect 6457 16399 6515 16405
rect 7193 16439 7251 16445
rect 7193 16405 7205 16439
rect 7239 16436 7251 16439
rect 8404 16436 8432 16476
rect 9278 16473 9290 16476
rect 9324 16473 9336 16507
rect 9278 16467 9336 16473
rect 9950 16464 9956 16516
rect 10008 16504 10014 16516
rect 10897 16504 10925 16544
rect 12066 16532 12072 16584
rect 12124 16572 12130 16584
rect 13262 16572 13268 16584
rect 12124 16544 13268 16572
rect 12124 16532 12130 16544
rect 13262 16532 13268 16544
rect 13320 16532 13326 16584
rect 10008 16476 10925 16504
rect 10956 16507 11014 16513
rect 10008 16464 10014 16476
rect 10956 16473 10968 16507
rect 11002 16504 11014 16507
rect 12710 16504 12716 16516
rect 11002 16476 12716 16504
rect 11002 16473 11014 16476
rect 10956 16467 11014 16473
rect 12710 16464 12716 16476
rect 12768 16464 12774 16516
rect 7239 16408 8432 16436
rect 7239 16405 7251 16408
rect 7193 16399 7251 16405
rect 9582 16396 9588 16448
rect 9640 16436 9646 16448
rect 10413 16439 10471 16445
rect 10413 16436 10425 16439
rect 9640 16408 10425 16436
rect 9640 16396 9646 16408
rect 10413 16405 10425 16408
rect 10459 16405 10471 16439
rect 10413 16399 10471 16405
rect 10594 16396 10600 16448
rect 10652 16436 10658 16448
rect 11238 16436 11244 16448
rect 10652 16408 11244 16436
rect 10652 16396 10658 16408
rect 11238 16396 11244 16408
rect 11296 16396 11302 16448
rect 12066 16436 12072 16448
rect 12027 16408 12072 16436
rect 12066 16396 12072 16408
rect 12124 16396 12130 16448
rect 12437 16439 12495 16445
rect 12437 16405 12449 16439
rect 12483 16436 12495 16439
rect 12989 16439 13047 16445
rect 12989 16436 13001 16439
rect 12483 16408 13001 16436
rect 12483 16405 12495 16408
rect 12437 16399 12495 16405
rect 12989 16405 13001 16408
rect 13035 16436 13047 16439
rect 13262 16436 13268 16448
rect 13035 16408 13268 16436
rect 13035 16405 13047 16408
rect 12989 16399 13047 16405
rect 13262 16396 13268 16408
rect 13320 16436 13326 16448
rect 13372 16445 13400 16612
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 15746 16572 15752 16584
rect 15707 16544 15752 16572
rect 15746 16532 15752 16544
rect 15804 16532 15810 16584
rect 16022 16581 16028 16584
rect 16016 16535 16028 16581
rect 16080 16572 16086 16584
rect 17512 16572 17540 16671
rect 18322 16572 18328 16584
rect 16080 16544 16116 16572
rect 16546 16544 18328 16572
rect 16022 16532 16028 16535
rect 16080 16532 16086 16544
rect 13446 16464 13452 16516
rect 13504 16504 13510 16516
rect 14338 16507 14396 16513
rect 14338 16504 14350 16507
rect 13504 16476 14350 16504
rect 13504 16464 13510 16476
rect 14338 16473 14350 16476
rect 14384 16473 14396 16507
rect 14338 16467 14396 16473
rect 15930 16464 15936 16516
rect 15988 16504 15994 16516
rect 16546 16504 16574 16544
rect 18322 16532 18328 16544
rect 18380 16532 18386 16584
rect 18877 16575 18935 16581
rect 18877 16541 18889 16575
rect 18923 16572 18935 16575
rect 19245 16575 19303 16581
rect 19245 16572 19257 16575
rect 18923 16544 19257 16572
rect 18923 16541 18935 16544
rect 18877 16535 18935 16541
rect 19245 16541 19257 16544
rect 19291 16572 19303 16575
rect 19291 16544 19748 16572
rect 19291 16541 19303 16544
rect 19245 16535 19303 16541
rect 19720 16516 19748 16544
rect 20806 16532 20812 16584
rect 20864 16572 20870 16584
rect 20901 16575 20959 16581
rect 20901 16572 20913 16575
rect 20864 16544 20913 16572
rect 20864 16532 20870 16544
rect 20901 16541 20913 16544
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 15988 16476 16574 16504
rect 15988 16464 15994 16476
rect 18230 16464 18236 16516
rect 18288 16504 18294 16516
rect 18610 16507 18668 16513
rect 18610 16504 18622 16507
rect 18288 16476 18622 16504
rect 18288 16464 18294 16476
rect 18610 16473 18622 16476
rect 18656 16504 18668 16507
rect 18966 16504 18972 16516
rect 18656 16476 18972 16504
rect 18656 16473 18668 16476
rect 18610 16467 18668 16473
rect 18966 16464 18972 16476
rect 19024 16464 19030 16516
rect 19490 16507 19548 16513
rect 19490 16504 19502 16507
rect 19076 16476 19502 16504
rect 13357 16439 13415 16445
rect 13357 16436 13369 16439
rect 13320 16408 13369 16436
rect 13320 16396 13326 16408
rect 13357 16405 13369 16408
rect 13403 16405 13415 16439
rect 13357 16399 13415 16405
rect 14734 16396 14740 16448
rect 14792 16436 14798 16448
rect 15473 16439 15531 16445
rect 15473 16436 15485 16439
rect 14792 16408 15485 16436
rect 14792 16396 14798 16408
rect 15473 16405 15485 16408
rect 15519 16405 15531 16439
rect 15473 16399 15531 16405
rect 17129 16439 17187 16445
rect 17129 16405 17141 16439
rect 17175 16436 17187 16439
rect 18690 16436 18696 16448
rect 17175 16408 18696 16436
rect 17175 16405 17187 16408
rect 17129 16399 17187 16405
rect 18690 16396 18696 16408
rect 18748 16436 18754 16448
rect 19076 16436 19104 16476
rect 19490 16473 19502 16476
rect 19536 16473 19548 16507
rect 19490 16467 19548 16473
rect 19702 16464 19708 16516
rect 19760 16464 19766 16516
rect 19978 16464 19984 16516
rect 20036 16504 20042 16516
rect 20036 16476 20208 16504
rect 20036 16464 20042 16476
rect 20180 16448 20208 16476
rect 18748 16408 19104 16436
rect 18748 16396 18754 16408
rect 19150 16396 19156 16448
rect 19208 16436 19214 16448
rect 20070 16436 20076 16448
rect 19208 16408 20076 16436
rect 19208 16396 19214 16408
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 20162 16396 20168 16448
rect 20220 16436 20226 16448
rect 20625 16439 20683 16445
rect 20625 16436 20637 16439
rect 20220 16408 20637 16436
rect 20220 16396 20226 16408
rect 20625 16405 20637 16408
rect 20671 16405 20683 16439
rect 21082 16436 21088 16448
rect 21043 16408 21088 16436
rect 20625 16399 20683 16405
rect 21082 16396 21088 16408
rect 21140 16396 21146 16448
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 4154 16232 4160 16244
rect 4115 16204 4160 16232
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 5261 16235 5319 16241
rect 5261 16201 5273 16235
rect 5307 16232 5319 16235
rect 5350 16232 5356 16244
rect 5307 16204 5356 16232
rect 5307 16201 5319 16204
rect 5261 16195 5319 16201
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 6641 16235 6699 16241
rect 6641 16201 6653 16235
rect 6687 16232 6699 16235
rect 7466 16232 7472 16244
rect 6687 16204 7472 16232
rect 6687 16201 6699 16204
rect 6641 16195 6699 16201
rect 7466 16192 7472 16204
rect 7524 16192 7530 16244
rect 11885 16235 11943 16241
rect 11885 16232 11897 16235
rect 8689 16204 11897 16232
rect 4080 16136 5488 16164
rect 4080 16096 4108 16136
rect 3988 16068 4108 16096
rect 5169 16099 5227 16105
rect 3988 16037 4016 16068
rect 5169 16065 5181 16099
rect 5215 16096 5227 16099
rect 5215 16068 5396 16096
rect 5215 16065 5227 16068
rect 5169 16059 5227 16065
rect 3973 16031 4031 16037
rect 3973 15997 3985 16031
rect 4019 15997 4031 16031
rect 3973 15991 4031 15997
rect 4065 16031 4123 16037
rect 4065 15997 4077 16031
rect 4111 16028 4123 16031
rect 4614 16028 4620 16040
rect 4111 16000 4620 16028
rect 4111 15997 4123 16000
rect 4065 15991 4123 15997
rect 4614 15988 4620 16000
rect 4672 15988 4678 16040
rect 4522 15892 4528 15904
rect 4483 15864 4528 15892
rect 4522 15852 4528 15864
rect 4580 15852 4586 15904
rect 4798 15892 4804 15904
rect 4759 15864 4804 15892
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 5368 15892 5396 16068
rect 5460 16037 5488 16136
rect 6733 16099 6791 16105
rect 6733 16065 6745 16099
rect 6779 16096 6791 16099
rect 7650 16096 7656 16108
rect 6779 16068 7656 16096
rect 6779 16065 6791 16068
rect 6733 16059 6791 16065
rect 7650 16056 7656 16068
rect 7708 16056 7714 16108
rect 7742 16056 7748 16108
rect 7800 16096 7806 16108
rect 8689 16105 8717 16204
rect 11885 16201 11897 16204
rect 11931 16201 11943 16235
rect 12802 16232 12808 16244
rect 11885 16195 11943 16201
rect 12406 16204 12808 16232
rect 12406 16164 12434 16204
rect 12802 16192 12808 16204
rect 12860 16192 12866 16244
rect 18049 16235 18107 16241
rect 18049 16201 18061 16235
rect 18095 16201 18107 16235
rect 18049 16195 18107 16201
rect 20349 16235 20407 16241
rect 20349 16201 20361 16235
rect 20395 16232 20407 16235
rect 20438 16232 20444 16244
rect 20395 16204 20444 16232
rect 20395 16201 20407 16204
rect 20349 16195 20407 16201
rect 9600 16136 12434 16164
rect 16936 16167 16994 16173
rect 8674 16099 8732 16105
rect 8674 16096 8686 16099
rect 7800 16068 8686 16096
rect 7800 16056 7806 16068
rect 8674 16065 8686 16068
rect 8720 16065 8732 16099
rect 8674 16059 8732 16065
rect 5445 16031 5503 16037
rect 5445 15997 5457 16031
rect 5491 15997 5503 16031
rect 5445 15991 5503 15997
rect 6549 16031 6607 16037
rect 6549 15997 6561 16031
rect 6595 16028 6607 16031
rect 6914 16028 6920 16040
rect 6595 16000 6920 16028
rect 6595 15997 6607 16000
rect 6549 15991 6607 15997
rect 5460 15960 5488 15991
rect 6914 15988 6920 16000
rect 6972 16028 6978 16040
rect 7374 16028 7380 16040
rect 6972 16000 7380 16028
rect 6972 15988 6978 16000
rect 7374 15988 7380 16000
rect 7432 15988 7438 16040
rect 8941 16031 8999 16037
rect 8941 15997 8953 16031
rect 8987 16028 8999 16031
rect 9122 16028 9128 16040
rect 8987 16000 9128 16028
rect 8987 15997 8999 16000
rect 8941 15991 8999 15997
rect 9122 15988 9128 16000
rect 9180 15988 9186 16040
rect 9600 15960 9628 16136
rect 16936 16133 16948 16167
rect 16982 16164 16994 16167
rect 17034 16164 17040 16176
rect 16982 16136 17040 16164
rect 16982 16133 16994 16136
rect 16936 16127 16994 16133
rect 17034 16124 17040 16136
rect 17092 16124 17098 16176
rect 17126 16124 17132 16176
rect 17184 16164 17190 16176
rect 18064 16164 18092 16195
rect 20438 16192 20444 16204
rect 20496 16192 20502 16244
rect 20898 16232 20904 16244
rect 20859 16204 20904 16232
rect 20898 16192 20904 16204
rect 20956 16192 20962 16244
rect 18754 16167 18812 16173
rect 18754 16164 18766 16167
rect 17184 16136 18766 16164
rect 17184 16124 17190 16136
rect 18754 16133 18766 16136
rect 18800 16133 18812 16167
rect 18754 16127 18812 16133
rect 10341 16099 10399 16105
rect 10341 16065 10353 16099
rect 10387 16096 10399 16099
rect 10502 16096 10508 16108
rect 10387 16068 10508 16096
rect 10387 16065 10399 16068
rect 10341 16059 10399 16065
rect 10502 16056 10508 16068
rect 10560 16056 10566 16108
rect 12250 16056 12256 16108
rect 12308 16096 12314 16108
rect 12998 16099 13056 16105
rect 12998 16096 13010 16099
rect 12308 16068 13010 16096
rect 12308 16056 12314 16068
rect 12998 16065 13010 16068
rect 13044 16065 13056 16099
rect 12998 16059 13056 16065
rect 13808 16099 13866 16105
rect 13808 16065 13820 16099
rect 13854 16096 13866 16099
rect 14274 16096 14280 16108
rect 13854 16068 14280 16096
rect 13854 16065 13866 16068
rect 13808 16059 13866 16065
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 20165 16099 20223 16105
rect 20165 16065 20177 16099
rect 20211 16096 20223 16099
rect 20714 16096 20720 16108
rect 20211 16068 20576 16096
rect 20675 16068 20720 16096
rect 20211 16065 20223 16068
rect 20165 16059 20223 16065
rect 10597 16031 10655 16037
rect 10597 15997 10609 16031
rect 10643 16028 10655 16031
rect 10686 16028 10692 16040
rect 10643 16000 10692 16028
rect 10643 15997 10655 16000
rect 10597 15991 10655 15997
rect 10686 15988 10692 16000
rect 10744 16028 10750 16040
rect 13262 16028 13268 16040
rect 10744 16000 11008 16028
rect 13223 16000 13268 16028
rect 10744 15988 10750 16000
rect 5460 15932 7696 15960
rect 5810 15892 5816 15904
rect 5368 15864 5816 15892
rect 5810 15852 5816 15864
rect 5868 15852 5874 15904
rect 7098 15892 7104 15904
rect 7059 15864 7104 15892
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 7466 15852 7472 15904
rect 7524 15892 7530 15904
rect 7561 15895 7619 15901
rect 7561 15892 7573 15895
rect 7524 15864 7573 15892
rect 7524 15852 7530 15864
rect 7561 15861 7573 15864
rect 7607 15861 7619 15895
rect 7668 15892 7696 15932
rect 8956 15932 9628 15960
rect 8956 15892 8984 15932
rect 7668 15864 8984 15892
rect 9217 15895 9275 15901
rect 7561 15855 7619 15861
rect 9217 15861 9229 15895
rect 9263 15892 9275 15895
rect 9398 15892 9404 15904
rect 9263 15864 9404 15892
rect 9263 15861 9275 15864
rect 9217 15855 9275 15861
rect 9398 15852 9404 15864
rect 9456 15852 9462 15904
rect 10980 15901 11008 16000
rect 13262 15988 13268 16000
rect 13320 16028 13326 16040
rect 13541 16031 13599 16037
rect 13541 16028 13553 16031
rect 13320 16000 13553 16028
rect 13320 15988 13326 16000
rect 13541 15997 13553 16000
rect 13587 15997 13599 16031
rect 16669 16031 16727 16037
rect 16669 16028 16681 16031
rect 13541 15991 13599 15997
rect 16546 16000 16681 16028
rect 14921 15963 14979 15969
rect 14921 15929 14933 15963
rect 14967 15960 14979 15963
rect 15470 15960 15476 15972
rect 14967 15932 15476 15960
rect 14967 15929 14979 15932
rect 14921 15923 14979 15929
rect 15470 15920 15476 15932
rect 15528 15920 15534 15972
rect 10965 15895 11023 15901
rect 10965 15861 10977 15895
rect 11011 15892 11023 15895
rect 11054 15892 11060 15904
rect 11011 15864 11060 15892
rect 11011 15861 11023 15864
rect 10965 15855 11023 15861
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 12158 15852 12164 15904
rect 12216 15892 12222 15904
rect 14642 15892 14648 15904
rect 12216 15864 14648 15892
rect 12216 15852 12222 15864
rect 14642 15852 14648 15864
rect 14700 15852 14706 15904
rect 15194 15892 15200 15904
rect 15155 15864 15200 15892
rect 15194 15852 15200 15864
rect 15252 15892 15258 15904
rect 15657 15895 15715 15901
rect 15657 15892 15669 15895
rect 15252 15864 15669 15892
rect 15252 15852 15258 15864
rect 15657 15861 15669 15864
rect 15703 15892 15715 15895
rect 15746 15892 15752 15904
rect 15703 15864 15752 15892
rect 15703 15861 15715 15864
rect 15657 15855 15715 15861
rect 15746 15852 15752 15864
rect 15804 15892 15810 15904
rect 16209 15895 16267 15901
rect 16209 15892 16221 15895
rect 15804 15864 16221 15892
rect 15804 15852 15810 15864
rect 16209 15861 16221 15864
rect 16255 15892 16267 15895
rect 16546 15892 16574 16000
rect 16669 15997 16681 16000
rect 16715 15997 16727 16031
rect 18506 16028 18512 16040
rect 18467 16000 18512 16028
rect 16669 15991 16727 15997
rect 18506 15988 18512 16000
rect 18564 15988 18570 16040
rect 20548 16028 20576 16068
rect 20714 16056 20720 16068
rect 20772 16056 20778 16108
rect 20990 16028 20996 16040
rect 20548 16000 20996 16028
rect 20990 15988 20996 16000
rect 21048 15988 21054 16040
rect 16255 15864 16574 15892
rect 19889 15895 19947 15901
rect 16255 15861 16267 15864
rect 16209 15855 16267 15861
rect 19889 15861 19901 15895
rect 19935 15892 19947 15895
rect 20070 15892 20076 15904
rect 19935 15864 20076 15892
rect 19935 15861 19947 15864
rect 19889 15855 19947 15861
rect 20070 15852 20076 15864
rect 20128 15852 20134 15904
rect 21266 15892 21272 15904
rect 21227 15864 21272 15892
rect 21266 15852 21272 15864
rect 21324 15852 21330 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 11146 15688 11152 15700
rect 7852 15660 11152 15688
rect 6914 15620 6920 15632
rect 5736 15592 6920 15620
rect 5736 15561 5764 15592
rect 6914 15580 6920 15592
rect 6972 15580 6978 15632
rect 5721 15555 5779 15561
rect 5721 15521 5733 15555
rect 5767 15521 5779 15555
rect 5721 15515 5779 15521
rect 6733 15555 6791 15561
rect 6733 15521 6745 15555
rect 6779 15521 6791 15555
rect 6733 15515 6791 15521
rect 6825 15555 6883 15561
rect 6825 15521 6837 15555
rect 6871 15552 6883 15555
rect 7098 15552 7104 15564
rect 6871 15524 7104 15552
rect 6871 15521 6883 15524
rect 6825 15515 6883 15521
rect 5902 15484 5908 15496
rect 5863 15456 5908 15484
rect 5902 15444 5908 15456
rect 5960 15444 5966 15496
rect 6748 15484 6776 15515
rect 7098 15512 7104 15524
rect 7156 15512 7162 15564
rect 7852 15484 7880 15660
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 11698 15648 11704 15700
rect 11756 15688 11762 15700
rect 14366 15688 14372 15700
rect 11756 15660 14372 15688
rect 11756 15648 11762 15660
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 7926 15580 7932 15632
rect 7984 15620 7990 15632
rect 9769 15623 9827 15629
rect 9769 15620 9781 15623
rect 7984 15592 9781 15620
rect 7984 15580 7990 15592
rect 9769 15589 9781 15592
rect 9815 15620 9827 15623
rect 10134 15620 10140 15632
rect 9815 15592 10140 15620
rect 9815 15589 9827 15592
rect 9769 15583 9827 15589
rect 10134 15580 10140 15592
rect 10192 15580 10198 15632
rect 11164 15592 11376 15620
rect 11164 15552 11192 15592
rect 11072 15524 11192 15552
rect 6748 15456 7880 15484
rect 10318 15444 10324 15496
rect 10376 15484 10382 15496
rect 11072 15484 11100 15524
rect 10376 15456 11100 15484
rect 11149 15487 11207 15493
rect 10376 15444 10382 15456
rect 11149 15453 11161 15487
rect 11195 15453 11207 15487
rect 11348 15484 11376 15592
rect 13090 15487 13148 15493
rect 13090 15484 13102 15487
rect 11348 15456 13102 15484
rect 11149 15447 11207 15453
rect 13090 15453 13102 15456
rect 13136 15453 13148 15487
rect 13090 15447 13148 15453
rect 5813 15419 5871 15425
rect 5813 15385 5825 15419
rect 5859 15416 5871 15419
rect 6086 15416 6092 15428
rect 5859 15388 6092 15416
rect 5859 15385 5871 15388
rect 5813 15379 5871 15385
rect 6086 15376 6092 15388
rect 6144 15376 6150 15428
rect 6917 15419 6975 15425
rect 6917 15416 6929 15419
rect 6288 15388 6929 15416
rect 4614 15348 4620 15360
rect 4575 15320 4620 15348
rect 4614 15308 4620 15320
rect 4672 15308 4678 15360
rect 6288 15357 6316 15388
rect 6917 15385 6929 15388
rect 6963 15385 6975 15419
rect 6917 15379 6975 15385
rect 7558 15376 7564 15428
rect 7616 15416 7622 15428
rect 7929 15419 7987 15425
rect 7929 15416 7941 15419
rect 7616 15388 7941 15416
rect 7616 15376 7622 15388
rect 7929 15385 7941 15388
rect 7975 15385 7987 15419
rect 7929 15379 7987 15385
rect 9582 15376 9588 15428
rect 9640 15416 9646 15428
rect 10882 15419 10940 15425
rect 10882 15416 10894 15419
rect 9640 15388 10894 15416
rect 9640 15376 9646 15388
rect 10882 15385 10894 15388
rect 10928 15385 10940 15419
rect 10882 15379 10940 15385
rect 6273 15351 6331 15357
rect 6273 15317 6285 15351
rect 6319 15317 6331 15351
rect 7282 15348 7288 15360
rect 7243 15320 7288 15348
rect 6273 15311 6331 15317
rect 7282 15308 7288 15320
rect 7340 15308 7346 15360
rect 7650 15348 7656 15360
rect 7611 15320 7656 15348
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 9122 15348 9128 15360
rect 9083 15320 9128 15348
rect 9122 15308 9128 15320
rect 9180 15308 9186 15360
rect 11054 15308 11060 15360
rect 11112 15348 11118 15360
rect 11164 15348 11192 15447
rect 13262 15444 13268 15496
rect 13320 15484 13326 15496
rect 13357 15487 13415 15493
rect 13357 15484 13369 15487
rect 13320 15456 13369 15484
rect 13320 15444 13326 15456
rect 13357 15453 13369 15456
rect 13403 15484 13415 15487
rect 15565 15487 15623 15493
rect 15565 15484 15577 15487
rect 13403 15456 13768 15484
rect 13403 15453 13415 15456
rect 13357 15447 13415 15453
rect 13740 15360 13768 15456
rect 15212 15456 15577 15484
rect 15212 15428 15240 15456
rect 15565 15453 15577 15456
rect 15611 15484 15623 15487
rect 15841 15487 15899 15493
rect 15841 15484 15853 15487
rect 15611 15456 15853 15484
rect 15611 15453 15623 15456
rect 15565 15447 15623 15453
rect 15841 15453 15853 15456
rect 15887 15484 15899 15487
rect 16390 15484 16396 15496
rect 15887 15456 16396 15484
rect 15887 15453 15899 15456
rect 15841 15447 15899 15453
rect 16390 15444 16396 15456
rect 16448 15484 16454 15496
rect 17497 15487 17555 15493
rect 17497 15484 17509 15487
rect 16448 15456 17509 15484
rect 16448 15444 16454 15456
rect 17497 15453 17509 15456
rect 17543 15484 17555 15487
rect 18141 15487 18199 15493
rect 18141 15484 18153 15487
rect 17543 15456 18153 15484
rect 17543 15453 17555 15456
rect 17497 15447 17555 15453
rect 18141 15453 18153 15456
rect 18187 15484 18199 15487
rect 18506 15484 18512 15496
rect 18187 15456 18512 15484
rect 18187 15453 18199 15456
rect 18141 15447 18199 15453
rect 18506 15444 18512 15456
rect 18564 15484 18570 15496
rect 18785 15487 18843 15493
rect 18785 15484 18797 15487
rect 18564 15456 18797 15484
rect 18564 15444 18570 15456
rect 18785 15453 18797 15456
rect 18831 15484 18843 15487
rect 19245 15487 19303 15493
rect 19245 15484 19257 15487
rect 18831 15456 19257 15484
rect 18831 15453 18843 15456
rect 18785 15447 18843 15453
rect 19245 15453 19257 15456
rect 19291 15453 19303 15487
rect 19245 15447 19303 15453
rect 21266 15444 21272 15496
rect 21324 15484 21330 15496
rect 21361 15487 21419 15493
rect 21361 15484 21373 15487
rect 21324 15456 21373 15484
rect 21324 15444 21330 15456
rect 21361 15453 21373 15456
rect 21407 15453 21419 15487
rect 21361 15447 21419 15453
rect 15194 15376 15200 15428
rect 15252 15376 15258 15428
rect 15286 15376 15292 15428
rect 15344 15425 15350 15428
rect 15344 15416 15356 15425
rect 15344 15388 15389 15416
rect 15344 15379 15356 15388
rect 15344 15376 15350 15379
rect 15470 15376 15476 15428
rect 15528 15416 15534 15428
rect 16086 15419 16144 15425
rect 16086 15416 16098 15419
rect 15528 15388 16098 15416
rect 15528 15376 15534 15388
rect 16086 15385 16098 15388
rect 16132 15385 16144 15419
rect 16086 15379 16144 15385
rect 21082 15376 21088 15428
rect 21140 15425 21146 15428
rect 21140 15416 21152 15425
rect 21140 15388 21185 15416
rect 21140 15379 21152 15388
rect 21140 15376 21146 15379
rect 11425 15351 11483 15357
rect 11425 15348 11437 15351
rect 11112 15320 11437 15348
rect 11112 15308 11118 15320
rect 11425 15317 11437 15320
rect 11471 15317 11483 15351
rect 11425 15311 11483 15317
rect 11698 15308 11704 15360
rect 11756 15348 11762 15360
rect 11977 15351 12035 15357
rect 11977 15348 11989 15351
rect 11756 15320 11989 15348
rect 11756 15308 11762 15320
rect 11977 15317 11989 15320
rect 12023 15317 12035 15351
rect 13722 15348 13728 15360
rect 13683 15320 13728 15348
rect 11977 15311 12035 15317
rect 13722 15308 13728 15320
rect 13780 15308 13786 15360
rect 14185 15351 14243 15357
rect 14185 15317 14197 15351
rect 14231 15348 14243 15351
rect 14274 15348 14280 15360
rect 14231 15320 14280 15348
rect 14231 15317 14243 15320
rect 14185 15311 14243 15317
rect 14274 15308 14280 15320
rect 14332 15348 14338 15360
rect 15102 15348 15108 15360
rect 14332 15320 15108 15348
rect 14332 15308 14338 15320
rect 15102 15308 15108 15320
rect 15160 15308 15166 15360
rect 17221 15351 17279 15357
rect 17221 15317 17233 15351
rect 17267 15348 17279 15351
rect 18046 15348 18052 15360
rect 17267 15320 18052 15348
rect 17267 15317 17279 15320
rect 17221 15311 17279 15317
rect 18046 15308 18052 15320
rect 18104 15308 18110 15360
rect 18506 15308 18512 15360
rect 18564 15348 18570 15360
rect 18690 15348 18696 15360
rect 18564 15320 18696 15348
rect 18564 15308 18570 15320
rect 18690 15308 18696 15320
rect 18748 15308 18754 15360
rect 19702 15348 19708 15360
rect 19663 15320 19708 15348
rect 19702 15308 19708 15320
rect 19760 15308 19766 15360
rect 19886 15308 19892 15360
rect 19944 15348 19950 15360
rect 19981 15351 20039 15357
rect 19981 15348 19993 15351
rect 19944 15320 19993 15348
rect 19944 15308 19950 15320
rect 19981 15317 19993 15320
rect 20027 15348 20039 15351
rect 20254 15348 20260 15360
rect 20027 15320 20260 15348
rect 20027 15317 20039 15320
rect 19981 15311 20039 15317
rect 20254 15308 20260 15320
rect 20312 15308 20318 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 4522 15104 4528 15156
rect 4580 15144 4586 15156
rect 4617 15147 4675 15153
rect 4617 15144 4629 15147
rect 4580 15116 4629 15144
rect 4580 15104 4586 15116
rect 4617 15113 4629 15116
rect 4663 15113 4675 15147
rect 6822 15144 6828 15156
rect 6783 15116 6828 15144
rect 4617 15107 4675 15113
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 8018 15104 8024 15156
rect 8076 15144 8082 15156
rect 12066 15144 12072 15156
rect 8076 15116 12072 15144
rect 8076 15104 8082 15116
rect 12066 15104 12072 15116
rect 12124 15104 12130 15156
rect 12342 15104 12348 15156
rect 12400 15144 12406 15156
rect 14921 15147 14979 15153
rect 14921 15144 14933 15147
rect 12400 15116 14933 15144
rect 12400 15104 12406 15116
rect 14921 15113 14933 15116
rect 14967 15144 14979 15147
rect 15286 15144 15292 15156
rect 14967 15116 15292 15144
rect 14967 15113 14979 15116
rect 14921 15107 14979 15113
rect 15286 15104 15292 15116
rect 15344 15104 15350 15156
rect 5721 15079 5779 15085
rect 5721 15045 5733 15079
rect 5767 15076 5779 15079
rect 6178 15076 6184 15088
rect 5767 15048 6184 15076
rect 5767 15045 5779 15048
rect 5721 15039 5779 15045
rect 6178 15036 6184 15048
rect 6236 15076 6242 15088
rect 6730 15076 6736 15088
rect 6236 15048 6736 15076
rect 6236 15036 6242 15048
rect 6730 15036 6736 15048
rect 6788 15036 6794 15088
rect 7285 15079 7343 15085
rect 7285 15045 7297 15079
rect 7331 15076 7343 15079
rect 7331 15048 8717 15076
rect 7331 15045 7343 15048
rect 7285 15039 7343 15045
rect 4525 15011 4583 15017
rect 4525 14977 4537 15011
rect 4571 15008 4583 15011
rect 4798 15008 4804 15020
rect 4571 14980 4804 15008
rect 4571 14977 4583 14980
rect 4525 14971 4583 14977
rect 4798 14968 4804 14980
rect 4856 14968 4862 15020
rect 5629 15011 5687 15017
rect 5629 14977 5641 15011
rect 5675 15008 5687 15011
rect 6365 15011 6423 15017
rect 6365 15008 6377 15011
rect 5675 14980 6377 15008
rect 5675 14977 5687 14980
rect 5629 14971 5687 14977
rect 6365 14977 6377 14980
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 7193 15011 7251 15017
rect 7193 14977 7205 15011
rect 7239 15008 7251 15011
rect 7558 15008 7564 15020
rect 7239 14980 7564 15008
rect 7239 14977 7251 14980
rect 7193 14971 7251 14977
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 8689 15008 8717 15048
rect 8864 15048 12434 15076
rect 8864 15008 8892 15048
rect 8689 14980 8892 15008
rect 9398 14968 9404 15020
rect 9456 15008 9462 15020
rect 10025 15011 10083 15017
rect 10025 15008 10037 15011
rect 9456 14980 10037 15008
rect 9456 14968 9462 14980
rect 10025 14977 10037 14980
rect 10071 14977 10083 15011
rect 12406 15008 12434 15048
rect 20070 15036 20076 15088
rect 20128 15036 20134 15088
rect 12894 15008 12900 15020
rect 12406 14980 12900 15008
rect 10025 14971 10083 14977
rect 12894 14968 12900 14980
rect 12952 14968 12958 15020
rect 13630 14968 13636 15020
rect 13688 15008 13694 15020
rect 16034 15011 16092 15017
rect 16034 15008 16046 15011
rect 13688 14980 16046 15008
rect 13688 14968 13694 14980
rect 16034 14977 16046 14980
rect 16080 14977 16092 15011
rect 16034 14971 16092 14977
rect 16301 15011 16359 15017
rect 16301 14977 16313 15011
rect 16347 15008 16359 15011
rect 16390 15008 16396 15020
rect 16347 14980 16396 15008
rect 16347 14977 16359 14980
rect 16301 14971 16359 14977
rect 16390 14968 16396 14980
rect 16448 14968 16454 15020
rect 17310 14968 17316 15020
rect 17368 15008 17374 15020
rect 19961 15011 20019 15017
rect 19961 15008 19973 15011
rect 17368 14980 19973 15008
rect 17368 14968 17374 14980
rect 19961 14977 19973 14980
rect 20007 15008 20019 15011
rect 20088 15008 20116 15036
rect 20007 14980 20116 15008
rect 20007 14977 20019 14980
rect 19961 14971 20019 14977
rect 4433 14943 4491 14949
rect 4433 14909 4445 14943
rect 4479 14909 4491 14943
rect 4433 14903 4491 14909
rect 5905 14943 5963 14949
rect 5905 14909 5917 14943
rect 5951 14940 5963 14943
rect 6730 14940 6736 14952
rect 5951 14912 6736 14940
rect 5951 14909 5963 14912
rect 5905 14903 5963 14909
rect 4448 14872 4476 14903
rect 6730 14900 6736 14912
rect 6788 14900 6794 14952
rect 7469 14943 7527 14949
rect 7469 14909 7481 14943
rect 7515 14940 7527 14943
rect 8018 14940 8024 14952
rect 7515 14912 8024 14940
rect 7515 14909 7527 14912
rect 7469 14903 7527 14909
rect 8018 14900 8024 14912
rect 8076 14900 8082 14952
rect 9122 14900 9128 14952
rect 9180 14940 9186 14952
rect 9769 14943 9827 14949
rect 9769 14940 9781 14943
rect 9180 14912 9781 14940
rect 9180 14900 9186 14912
rect 9769 14909 9781 14912
rect 9815 14909 9827 14943
rect 16408 14940 16436 14968
rect 16761 14943 16819 14949
rect 16761 14940 16773 14943
rect 16408 14912 16773 14940
rect 9769 14903 9827 14909
rect 16761 14909 16773 14912
rect 16807 14940 16819 14943
rect 17129 14943 17187 14949
rect 17129 14940 17141 14943
rect 16807 14912 17141 14940
rect 16807 14909 16819 14912
rect 16761 14903 16819 14909
rect 17129 14909 17141 14912
rect 17175 14940 17187 14943
rect 17681 14943 17739 14949
rect 17681 14940 17693 14943
rect 17175 14912 17693 14940
rect 17175 14909 17187 14912
rect 17129 14903 17187 14909
rect 17681 14909 17693 14912
rect 17727 14940 17739 14943
rect 18049 14943 18107 14949
rect 18049 14940 18061 14943
rect 17727 14912 18061 14940
rect 17727 14909 17739 14912
rect 17681 14903 17739 14909
rect 18049 14909 18061 14912
rect 18095 14940 18107 14943
rect 18693 14943 18751 14949
rect 18693 14940 18705 14943
rect 18095 14912 18705 14940
rect 18095 14909 18107 14912
rect 18049 14903 18107 14909
rect 18693 14909 18705 14912
rect 18739 14940 18751 14943
rect 19429 14943 19487 14949
rect 19429 14940 19441 14943
rect 18739 14912 19441 14940
rect 18739 14909 18751 14912
rect 18693 14903 18751 14909
rect 19429 14909 19441 14912
rect 19475 14940 19487 14943
rect 19702 14940 19708 14952
rect 19475 14912 19708 14940
rect 19475 14909 19487 14912
rect 19429 14903 19487 14909
rect 9674 14872 9680 14884
rect 4448 14844 9680 14872
rect 9674 14832 9680 14844
rect 9732 14832 9738 14884
rect 4985 14807 5043 14813
rect 4985 14773 4997 14807
rect 5031 14804 5043 14807
rect 5074 14804 5080 14816
rect 5031 14776 5080 14804
rect 5031 14773 5043 14776
rect 4985 14767 5043 14773
rect 5074 14764 5080 14776
rect 5132 14764 5138 14816
rect 5261 14807 5319 14813
rect 5261 14773 5273 14807
rect 5307 14804 5319 14807
rect 5350 14804 5356 14816
rect 5307 14776 5356 14804
rect 5307 14773 5319 14776
rect 5261 14767 5319 14773
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 9784 14804 9812 14903
rect 19702 14900 19708 14912
rect 19760 14900 19766 14952
rect 11054 14832 11060 14884
rect 11112 14872 11118 14884
rect 11517 14875 11575 14881
rect 11517 14872 11529 14875
rect 11112 14844 11529 14872
rect 11112 14832 11118 14844
rect 11517 14841 11529 14844
rect 11563 14841 11575 14875
rect 21542 14872 21548 14884
rect 11517 14835 11575 14841
rect 20640 14844 21548 14872
rect 11072 14804 11100 14832
rect 9784 14776 11100 14804
rect 11146 14764 11152 14816
rect 11204 14804 11210 14816
rect 12250 14804 12256 14816
rect 11204 14776 12256 14804
rect 11204 14764 11210 14776
rect 12250 14764 12256 14776
rect 12308 14764 12314 14816
rect 13722 14764 13728 14816
rect 13780 14804 13786 14816
rect 14185 14807 14243 14813
rect 14185 14804 14197 14807
rect 13780 14776 14197 14804
rect 13780 14764 13786 14776
rect 14185 14773 14197 14776
rect 14231 14804 14243 14807
rect 14553 14807 14611 14813
rect 14553 14804 14565 14807
rect 14231 14776 14565 14804
rect 14231 14773 14243 14776
rect 14185 14767 14243 14773
rect 14553 14773 14565 14776
rect 14599 14804 14611 14807
rect 15194 14804 15200 14816
rect 14599 14776 15200 14804
rect 14599 14773 14611 14776
rect 14553 14767 14611 14773
rect 15194 14764 15200 14776
rect 15252 14764 15258 14816
rect 18046 14764 18052 14816
rect 18104 14804 18110 14816
rect 19061 14807 19119 14813
rect 19061 14804 19073 14807
rect 18104 14776 19073 14804
rect 18104 14764 18110 14776
rect 19061 14773 19073 14776
rect 19107 14804 19119 14807
rect 20640 14804 20668 14844
rect 21542 14832 21548 14844
rect 21600 14832 21606 14884
rect 21082 14804 21088 14816
rect 19107 14776 20668 14804
rect 20995 14776 21088 14804
rect 19107 14773 19119 14776
rect 19061 14767 19119 14773
rect 21082 14764 21088 14776
rect 21140 14804 21146 14816
rect 22186 14804 22192 14816
rect 21140 14776 22192 14804
rect 21140 14764 21146 14776
rect 22186 14764 22192 14776
rect 22244 14764 22250 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 3326 14600 3332 14612
rect 3287 14572 3332 14600
rect 3326 14560 3332 14572
rect 3384 14600 3390 14612
rect 3384 14572 4292 14600
rect 3384 14560 3390 14572
rect 4264 14473 4292 14572
rect 4522 14560 4528 14612
rect 4580 14600 4586 14612
rect 6178 14600 6184 14612
rect 4580 14572 6184 14600
rect 4580 14560 4586 14572
rect 6178 14560 6184 14572
rect 6236 14560 6242 14612
rect 7653 14603 7711 14609
rect 7653 14569 7665 14603
rect 7699 14600 7711 14603
rect 7834 14600 7840 14612
rect 7699 14572 7840 14600
rect 7699 14569 7711 14572
rect 7653 14563 7711 14569
rect 7834 14560 7840 14572
rect 7892 14560 7898 14612
rect 9858 14600 9864 14612
rect 9600 14572 9864 14600
rect 9600 14532 9628 14572
rect 9858 14560 9864 14572
rect 9916 14600 9922 14612
rect 11698 14600 11704 14612
rect 9916 14572 11704 14600
rect 9916 14560 9922 14572
rect 11698 14560 11704 14572
rect 11756 14560 11762 14612
rect 13262 14560 13268 14612
rect 13320 14600 13326 14612
rect 16209 14603 16267 14609
rect 16209 14600 16221 14603
rect 13320 14572 16221 14600
rect 13320 14560 13326 14572
rect 16209 14569 16221 14572
rect 16255 14569 16267 14603
rect 16209 14563 16267 14569
rect 5092 14504 9628 14532
rect 4157 14467 4215 14473
rect 4157 14433 4169 14467
rect 4203 14433 4215 14467
rect 4157 14427 4215 14433
rect 4249 14467 4307 14473
rect 4249 14433 4261 14467
rect 4295 14433 4307 14467
rect 4249 14427 4307 14433
rect 4172 14396 4200 14427
rect 4798 14424 4804 14476
rect 4856 14464 4862 14476
rect 5092 14473 5120 14504
rect 5077 14467 5135 14473
rect 5077 14464 5089 14467
rect 4856 14436 5089 14464
rect 4856 14424 4862 14436
rect 5077 14433 5089 14436
rect 5123 14433 5135 14467
rect 5077 14427 5135 14433
rect 7101 14467 7159 14473
rect 7101 14433 7113 14467
rect 7147 14433 7159 14467
rect 14550 14464 14556 14476
rect 7101 14427 7159 14433
rect 10520 14436 14556 14464
rect 4172 14368 4292 14396
rect 4264 14328 4292 14368
rect 4430 14356 4436 14408
rect 4488 14396 4494 14408
rect 5261 14399 5319 14405
rect 5261 14396 5273 14399
rect 4488 14368 5273 14396
rect 4488 14356 4494 14368
rect 5261 14365 5273 14368
rect 5307 14365 5319 14399
rect 5261 14359 5319 14365
rect 5353 14399 5411 14405
rect 5353 14365 5365 14399
rect 5399 14396 5411 14399
rect 5442 14396 5448 14408
rect 5399 14368 5448 14396
rect 5399 14365 5411 14368
rect 5353 14359 5411 14365
rect 5442 14356 5448 14368
rect 5500 14356 5506 14408
rect 7116 14396 7144 14427
rect 9766 14396 9772 14408
rect 7116 14368 9772 14396
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 7098 14328 7104 14340
rect 4264 14300 7104 14328
rect 7098 14288 7104 14300
rect 7156 14288 7162 14340
rect 10318 14288 10324 14340
rect 10376 14337 10382 14340
rect 10376 14328 10388 14337
rect 10520 14328 10548 14436
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 10597 14399 10655 14405
rect 10597 14365 10609 14399
rect 10643 14396 10655 14399
rect 11054 14396 11060 14408
rect 10643 14368 11060 14396
rect 10643 14365 10655 14368
rect 10597 14359 10655 14365
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 14829 14399 14887 14405
rect 14829 14396 14841 14399
rect 14476 14368 14841 14396
rect 10376 14300 10548 14328
rect 10888 14300 12434 14328
rect 10376 14291 10388 14300
rect 10376 14288 10382 14291
rect 3878 14220 3884 14272
rect 3936 14260 3942 14272
rect 4341 14263 4399 14269
rect 4341 14260 4353 14263
rect 3936 14232 4353 14260
rect 3936 14220 3942 14232
rect 4341 14229 4353 14232
rect 4387 14229 4399 14263
rect 4706 14260 4712 14272
rect 4667 14232 4712 14260
rect 4341 14223 4399 14229
rect 4706 14220 4712 14232
rect 4764 14220 4770 14272
rect 5721 14263 5779 14269
rect 5721 14229 5733 14263
rect 5767 14260 5779 14263
rect 5810 14260 5816 14272
rect 5767 14232 5816 14260
rect 5767 14229 5779 14232
rect 5721 14223 5779 14229
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 6914 14220 6920 14272
rect 6972 14260 6978 14272
rect 7193 14263 7251 14269
rect 7193 14260 7205 14263
rect 6972 14232 7205 14260
rect 6972 14220 6978 14232
rect 7193 14229 7205 14232
rect 7239 14229 7251 14263
rect 7193 14223 7251 14229
rect 7282 14220 7288 14272
rect 7340 14260 7346 14272
rect 9214 14260 9220 14272
rect 7340 14232 7385 14260
rect 9175 14232 9220 14260
rect 7340 14220 7346 14232
rect 9214 14220 9220 14232
rect 9272 14260 9278 14272
rect 10888 14260 10916 14300
rect 9272 14232 10916 14260
rect 10965 14263 11023 14269
rect 9272 14220 9278 14232
rect 10965 14229 10977 14263
rect 11011 14260 11023 14263
rect 11054 14260 11060 14272
rect 11011 14232 11060 14260
rect 11011 14229 11023 14232
rect 10965 14223 11023 14229
rect 11054 14220 11060 14232
rect 11112 14220 11118 14272
rect 12406 14260 12434 14300
rect 13446 14260 13452 14272
rect 12406 14232 13452 14260
rect 13446 14220 13452 14232
rect 13504 14220 13510 14272
rect 13722 14220 13728 14272
rect 13780 14260 13786 14272
rect 14476 14269 14504 14368
rect 14829 14365 14841 14368
rect 14875 14365 14887 14399
rect 14829 14359 14887 14365
rect 14918 14288 14924 14340
rect 14976 14328 14982 14340
rect 15074 14331 15132 14337
rect 15074 14328 15086 14331
rect 14976 14300 15086 14328
rect 14976 14288 14982 14300
rect 15074 14297 15086 14300
rect 15120 14297 15132 14331
rect 16224 14328 16252 14563
rect 19518 14424 19524 14476
rect 19576 14464 19582 14476
rect 20070 14464 20076 14476
rect 19576 14436 20076 14464
rect 19576 14424 19582 14436
rect 20070 14424 20076 14436
rect 20128 14424 20134 14476
rect 16390 14356 16396 14408
rect 16448 14396 16454 14408
rect 16485 14399 16543 14405
rect 16485 14396 16497 14399
rect 16448 14368 16497 14396
rect 16448 14356 16454 14368
rect 16485 14365 16497 14368
rect 16531 14396 16543 14399
rect 18141 14399 18199 14405
rect 18141 14396 18153 14399
rect 16531 14368 18153 14396
rect 16531 14365 16543 14368
rect 16485 14359 16543 14365
rect 18141 14365 18153 14368
rect 18187 14396 18199 14399
rect 18509 14399 18567 14405
rect 18509 14396 18521 14399
rect 18187 14368 18521 14396
rect 18187 14365 18199 14368
rect 18141 14359 18199 14365
rect 18509 14365 18521 14368
rect 18555 14365 18567 14399
rect 19702 14396 19708 14408
rect 19615 14368 19708 14396
rect 18509 14359 18567 14365
rect 19702 14356 19708 14368
rect 19760 14396 19766 14408
rect 21266 14396 21272 14408
rect 19760 14368 21272 14396
rect 19760 14356 19766 14368
rect 21266 14356 21272 14368
rect 21324 14396 21330 14408
rect 21361 14399 21419 14405
rect 21361 14396 21373 14399
rect 21324 14368 21373 14396
rect 21324 14356 21330 14368
rect 21361 14365 21373 14368
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 16730 14331 16788 14337
rect 16730 14328 16742 14331
rect 16224 14300 16742 14328
rect 15074 14291 15132 14297
rect 16730 14297 16742 14300
rect 16776 14297 16788 14331
rect 20162 14328 20168 14340
rect 16730 14291 16788 14297
rect 19352 14300 20168 14328
rect 19352 14272 19380 14300
rect 20162 14288 20168 14300
rect 20220 14288 20226 14340
rect 21082 14288 21088 14340
rect 21140 14337 21146 14340
rect 21140 14328 21152 14337
rect 21140 14300 21185 14328
rect 21140 14291 21152 14300
rect 21140 14288 21146 14291
rect 14093 14263 14151 14269
rect 14093 14260 14105 14263
rect 13780 14232 14105 14260
rect 13780 14220 13786 14232
rect 14093 14229 14105 14232
rect 14139 14260 14151 14263
rect 14461 14263 14519 14269
rect 14461 14260 14473 14263
rect 14139 14232 14473 14260
rect 14139 14229 14151 14232
rect 14093 14223 14151 14229
rect 14461 14229 14473 14232
rect 14507 14229 14519 14263
rect 14461 14223 14519 14229
rect 17586 14220 17592 14272
rect 17644 14260 17650 14272
rect 17865 14263 17923 14269
rect 17865 14260 17877 14263
rect 17644 14232 17877 14260
rect 17644 14220 17650 14232
rect 17865 14229 17877 14232
rect 17911 14229 17923 14263
rect 19334 14260 19340 14272
rect 19295 14232 19340 14260
rect 17865 14223 17923 14229
rect 19334 14220 19340 14232
rect 19392 14220 19398 14272
rect 19886 14220 19892 14272
rect 19944 14260 19950 14272
rect 19981 14263 20039 14269
rect 19981 14260 19993 14263
rect 19944 14232 19993 14260
rect 19944 14220 19950 14232
rect 19981 14229 19993 14232
rect 20027 14229 20039 14263
rect 19981 14223 20039 14229
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 3697 14059 3755 14065
rect 3697 14025 3709 14059
rect 3743 14056 3755 14059
rect 3878 14056 3884 14068
rect 3743 14028 3884 14056
rect 3743 14025 3755 14028
rect 3697 14019 3755 14025
rect 3878 14016 3884 14028
rect 3936 14016 3942 14068
rect 4430 14016 4436 14068
rect 4488 14056 4494 14068
rect 4801 14059 4859 14065
rect 4801 14056 4813 14059
rect 4488 14028 4813 14056
rect 4488 14016 4494 14028
rect 4801 14025 4813 14028
rect 4847 14025 4859 14059
rect 4801 14019 4859 14025
rect 5261 14059 5319 14065
rect 5261 14025 5273 14059
rect 5307 14056 5319 14059
rect 5442 14056 5448 14068
rect 5307 14028 5448 14056
rect 5307 14025 5319 14028
rect 5261 14019 5319 14025
rect 5442 14016 5448 14028
rect 5500 14016 5506 14068
rect 9674 14016 9680 14068
rect 9732 14056 9738 14068
rect 9732 14028 12572 14056
rect 9732 14016 9738 14028
rect 7098 13948 7104 14000
rect 7156 13988 7162 14000
rect 10134 13988 10140 14000
rect 7156 13960 10140 13988
rect 7156 13948 7162 13960
rect 10134 13948 10140 13960
rect 10192 13948 10198 14000
rect 10318 13948 10324 14000
rect 10376 13997 10382 14000
rect 10376 13988 10388 13997
rect 12544 13988 12572 14028
rect 13170 14016 13176 14068
rect 13228 14056 13234 14068
rect 13630 14056 13636 14068
rect 13228 14028 13636 14056
rect 13228 14016 13234 14028
rect 13630 14016 13636 14028
rect 13688 14056 13694 14068
rect 14277 14059 14335 14065
rect 14277 14056 14289 14059
rect 13688 14028 14289 14056
rect 13688 14016 13694 14028
rect 14277 14025 14289 14028
rect 14323 14025 14335 14059
rect 19334 14056 19340 14068
rect 14277 14019 14335 14025
rect 14384 14028 19340 14056
rect 14384 13988 14412 14028
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 21634 14056 21640 14068
rect 19536 14028 21640 14056
rect 10376 13960 10421 13988
rect 12544 13960 14412 13988
rect 10376 13951 10388 13960
rect 10376 13948 10382 13951
rect 15286 13948 15292 14000
rect 15344 13988 15350 14000
rect 15390 13991 15448 13997
rect 15390 13988 15402 13991
rect 15344 13960 15402 13988
rect 15344 13948 15350 13960
rect 15390 13957 15402 13960
rect 15436 13957 15448 13991
rect 15390 13951 15448 13957
rect 16936 13991 16994 13997
rect 16936 13957 16948 13991
rect 16982 13988 16994 13991
rect 17586 13988 17592 14000
rect 16982 13960 17592 13988
rect 16982 13957 16994 13960
rect 16936 13951 16994 13957
rect 17586 13948 17592 13960
rect 17644 13948 17650 14000
rect 19058 13988 19064 14000
rect 18156 13960 19064 13988
rect 6086 13880 6092 13932
rect 6144 13920 6150 13932
rect 6730 13920 6736 13932
rect 6144 13892 6736 13920
rect 6144 13880 6150 13892
rect 6730 13880 6736 13892
rect 6788 13920 6794 13932
rect 9950 13920 9956 13932
rect 6788 13892 9956 13920
rect 6788 13880 6794 13892
rect 9950 13880 9956 13892
rect 10008 13880 10014 13932
rect 12526 13880 12532 13932
rect 12584 13920 12590 13932
rect 12877 13923 12935 13929
rect 12877 13920 12889 13923
rect 12584 13892 12889 13920
rect 12584 13880 12590 13892
rect 12877 13889 12889 13892
rect 12923 13889 12935 13923
rect 12877 13883 12935 13889
rect 10597 13855 10655 13861
rect 10597 13821 10609 13855
rect 10643 13852 10655 13855
rect 10873 13855 10931 13861
rect 10873 13852 10885 13855
rect 10643 13824 10885 13852
rect 10643 13821 10655 13824
rect 10597 13815 10655 13821
rect 10873 13821 10885 13824
rect 10919 13852 10931 13855
rect 11054 13852 11060 13864
rect 10919 13824 11060 13852
rect 10919 13821 10931 13824
rect 10873 13815 10931 13821
rect 8849 13787 8907 13793
rect 8849 13784 8861 13787
rect 8312 13756 8861 13784
rect 8312 13728 8340 13756
rect 8849 13753 8861 13756
rect 8895 13784 8907 13787
rect 8895 13756 9720 13784
rect 8895 13753 8907 13756
rect 8849 13747 8907 13753
rect 7837 13719 7895 13725
rect 7837 13685 7849 13719
rect 7883 13716 7895 13719
rect 8205 13719 8263 13725
rect 8205 13716 8217 13719
rect 7883 13688 8217 13716
rect 7883 13685 7895 13688
rect 7837 13679 7895 13685
rect 8205 13685 8217 13688
rect 8251 13716 8263 13719
rect 8294 13716 8300 13728
rect 8251 13688 8300 13716
rect 8251 13685 8263 13688
rect 8205 13679 8263 13685
rect 8294 13676 8300 13688
rect 8352 13676 8358 13728
rect 8386 13676 8392 13728
rect 8444 13716 8450 13728
rect 8481 13719 8539 13725
rect 8481 13716 8493 13719
rect 8444 13688 8493 13716
rect 8444 13676 8450 13688
rect 8481 13685 8493 13688
rect 8527 13685 8539 13719
rect 8481 13679 8539 13685
rect 8662 13676 8668 13728
rect 8720 13716 8726 13728
rect 9217 13719 9275 13725
rect 9217 13716 9229 13719
rect 8720 13688 9229 13716
rect 8720 13676 8726 13688
rect 9217 13685 9229 13688
rect 9263 13685 9275 13719
rect 9692 13716 9720 13756
rect 10612 13716 10640 13815
rect 11054 13812 11060 13824
rect 11112 13852 11118 13864
rect 12621 13855 12679 13861
rect 12621 13852 12633 13855
rect 11112 13824 12633 13852
rect 11112 13812 11118 13824
rect 12621 13821 12633 13824
rect 12667 13821 12679 13855
rect 15654 13852 15660 13864
rect 15615 13824 15660 13852
rect 12621 13815 12679 13821
rect 15654 13812 15660 13824
rect 15712 13852 15718 13864
rect 15933 13855 15991 13861
rect 15933 13852 15945 13855
rect 15712 13824 15945 13852
rect 15712 13812 15718 13824
rect 15933 13821 15945 13824
rect 15979 13852 15991 13855
rect 16669 13855 16727 13861
rect 16669 13852 16681 13855
rect 15979 13824 16681 13852
rect 15979 13821 15991 13824
rect 15933 13815 15991 13821
rect 16669 13821 16681 13824
rect 16715 13821 16727 13855
rect 18156 13852 18184 13960
rect 19058 13948 19064 13960
rect 19116 13948 19122 14000
rect 19536 13988 19564 14028
rect 21634 14016 21640 14028
rect 21692 14016 21698 14068
rect 19352 13960 19564 13988
rect 19720 13960 21312 13988
rect 19352 13920 19380 13960
rect 18708 13892 19380 13920
rect 18708 13852 18736 13892
rect 19426 13880 19432 13932
rect 19484 13929 19490 13932
rect 19720 13929 19748 13960
rect 21284 13932 21312 13960
rect 19484 13920 19496 13929
rect 19705 13923 19763 13929
rect 19484 13892 19529 13920
rect 19484 13883 19496 13892
rect 19705 13889 19717 13923
rect 19751 13889 19763 13923
rect 19705 13883 19763 13889
rect 19484 13880 19490 13883
rect 20162 13880 20168 13932
rect 20220 13920 20226 13932
rect 21094 13923 21152 13929
rect 21094 13920 21106 13923
rect 20220 13892 21106 13920
rect 20220 13880 20226 13892
rect 21094 13889 21106 13892
rect 21140 13889 21152 13923
rect 21094 13883 21152 13889
rect 21266 13880 21272 13932
rect 21324 13920 21330 13932
rect 21361 13923 21419 13929
rect 21361 13920 21373 13923
rect 21324 13892 21373 13920
rect 21324 13880 21330 13892
rect 21361 13889 21373 13892
rect 21407 13889 21419 13923
rect 21361 13883 21419 13889
rect 16669 13815 16727 13821
rect 18064 13824 18184 13852
rect 18340 13824 18736 13852
rect 18064 13793 18092 13824
rect 18340 13793 18368 13824
rect 18049 13787 18107 13793
rect 18049 13753 18061 13787
rect 18095 13753 18107 13787
rect 18049 13747 18107 13753
rect 18325 13787 18383 13793
rect 18325 13753 18337 13787
rect 18371 13753 18383 13787
rect 18325 13747 18383 13753
rect 9692 13688 10640 13716
rect 9217 13679 9275 13685
rect 13538 13676 13544 13728
rect 13596 13716 13602 13728
rect 14001 13719 14059 13725
rect 14001 13716 14013 13719
rect 13596 13688 14013 13716
rect 13596 13676 13602 13688
rect 14001 13685 14013 13688
rect 14047 13685 14059 13719
rect 14001 13679 14059 13685
rect 15010 13676 15016 13728
rect 15068 13716 15074 13728
rect 16850 13716 16856 13728
rect 15068 13688 16856 13716
rect 15068 13676 15074 13688
rect 16850 13676 16856 13688
rect 16908 13676 16914 13728
rect 17034 13676 17040 13728
rect 17092 13716 17098 13728
rect 17770 13716 17776 13728
rect 17092 13688 17776 13716
rect 17092 13676 17098 13688
rect 17770 13676 17776 13688
rect 17828 13716 17834 13728
rect 19981 13719 20039 13725
rect 19981 13716 19993 13719
rect 17828 13688 19993 13716
rect 17828 13676 17834 13688
rect 19981 13685 19993 13688
rect 20027 13685 20039 13719
rect 19981 13679 20039 13685
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 6730 13472 6736 13524
rect 6788 13512 6794 13524
rect 8662 13512 8668 13524
rect 6788 13484 8668 13512
rect 6788 13472 6794 13484
rect 8662 13472 8668 13484
rect 8720 13472 8726 13524
rect 10226 13512 10232 13524
rect 9048 13484 10232 13512
rect 6086 13444 6092 13456
rect 5092 13416 6092 13444
rect 5092 13385 5120 13416
rect 6086 13404 6092 13416
rect 6144 13404 6150 13456
rect 8573 13447 8631 13453
rect 8573 13413 8585 13447
rect 8619 13444 8631 13447
rect 9048 13444 9076 13484
rect 10226 13472 10232 13484
rect 10284 13472 10290 13524
rect 10689 13515 10747 13521
rect 10689 13481 10701 13515
rect 10735 13512 10747 13515
rect 11698 13512 11704 13524
rect 10735 13484 11704 13512
rect 10735 13481 10747 13484
rect 10689 13475 10747 13481
rect 11698 13472 11704 13484
rect 11756 13512 11762 13524
rect 11882 13512 11888 13524
rect 11756 13484 11888 13512
rect 11756 13472 11762 13484
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 12250 13472 12256 13524
rect 12308 13512 12314 13524
rect 12345 13515 12403 13521
rect 12345 13512 12357 13515
rect 12308 13484 12357 13512
rect 12308 13472 12314 13484
rect 12345 13481 12357 13484
rect 12391 13481 12403 13515
rect 12345 13475 12403 13481
rect 13538 13472 13544 13524
rect 13596 13512 13602 13524
rect 13596 13484 13952 13512
rect 13596 13472 13602 13484
rect 8619 13416 9076 13444
rect 8619 13413 8631 13416
rect 8573 13407 8631 13413
rect 5077 13379 5135 13385
rect 5077 13345 5089 13379
rect 5123 13345 5135 13379
rect 5258 13376 5264 13388
rect 5219 13348 5264 13376
rect 5077 13339 5135 13345
rect 5258 13336 5264 13348
rect 5316 13336 5322 13388
rect 8294 13336 8300 13388
rect 8352 13376 8358 13388
rect 9033 13379 9091 13385
rect 9033 13376 9045 13379
rect 8352 13348 9045 13376
rect 8352 13336 8358 13348
rect 9033 13345 9045 13348
rect 9079 13345 9091 13379
rect 9033 13339 9091 13345
rect 5442 13268 5448 13320
rect 5500 13308 5506 13320
rect 6454 13308 6460 13320
rect 5500 13280 6460 13308
rect 5500 13268 5506 13280
rect 6454 13268 6460 13280
rect 6512 13268 6518 13320
rect 6546 13268 6552 13320
rect 6604 13308 6610 13320
rect 7193 13311 7251 13317
rect 7193 13308 7205 13311
rect 6604 13280 7205 13308
rect 6604 13268 6610 13280
rect 7193 13277 7205 13280
rect 7239 13277 7251 13311
rect 7193 13271 7251 13277
rect 7460 13311 7518 13317
rect 7460 13277 7472 13311
rect 7506 13308 7518 13311
rect 9122 13308 9128 13320
rect 7506 13280 9128 13308
rect 7506 13277 7518 13280
rect 7460 13271 7518 13277
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 12066 13308 12072 13320
rect 12027 13280 12072 13308
rect 12066 13268 12072 13280
rect 12124 13308 12130 13320
rect 13722 13308 13728 13320
rect 12124 13280 13728 13308
rect 12124 13268 12130 13280
rect 13722 13268 13728 13280
rect 13780 13268 13786 13320
rect 13924 13308 13952 13484
rect 17862 13472 17868 13524
rect 17920 13512 17926 13524
rect 19245 13515 19303 13521
rect 19245 13512 19257 13515
rect 17920 13484 19257 13512
rect 17920 13472 17926 13484
rect 19245 13481 19257 13484
rect 19291 13481 19303 13515
rect 19245 13475 19303 13481
rect 20622 13472 20628 13524
rect 20680 13512 20686 13524
rect 21085 13515 21143 13521
rect 21085 13512 21097 13515
rect 20680 13484 21097 13512
rect 20680 13472 20686 13484
rect 21085 13481 21097 13484
rect 21131 13481 21143 13515
rect 21085 13475 21143 13481
rect 18230 13444 18236 13456
rect 18191 13416 18236 13444
rect 18230 13404 18236 13416
rect 18288 13404 18294 13456
rect 18782 13444 18788 13456
rect 18743 13416 18788 13444
rect 18782 13404 18788 13416
rect 18840 13404 18846 13456
rect 17494 13336 17500 13388
rect 17552 13376 17558 13388
rect 20625 13379 20683 13385
rect 17552 13348 18644 13376
rect 17552 13336 17558 13348
rect 15206 13311 15264 13317
rect 15206 13308 15218 13311
rect 13924 13280 15218 13308
rect 15206 13277 15218 13280
rect 15252 13277 15264 13311
rect 15470 13308 15476 13320
rect 15431 13280 15476 13308
rect 15206 13271 15264 13277
rect 15470 13268 15476 13280
rect 15528 13308 15534 13320
rect 15654 13308 15660 13320
rect 15528 13280 15660 13308
rect 15528 13268 15534 13280
rect 15654 13268 15660 13280
rect 15712 13308 15718 13320
rect 15749 13311 15807 13317
rect 15749 13308 15761 13311
rect 15712 13280 15761 13308
rect 15712 13268 15718 13280
rect 15749 13277 15761 13280
rect 15795 13308 15807 13311
rect 16209 13311 16267 13317
rect 16209 13308 16221 13311
rect 15795 13280 16221 13308
rect 15795 13277 15807 13280
rect 15749 13271 15807 13277
rect 16209 13277 16221 13280
rect 16255 13277 16267 13311
rect 16209 13271 16267 13277
rect 16298 13268 16304 13320
rect 16356 13308 16362 13320
rect 18616 13317 18644 13348
rect 20625 13345 20637 13379
rect 20671 13376 20683 13379
rect 21266 13376 21272 13388
rect 20671 13348 21272 13376
rect 20671 13345 20683 13348
rect 20625 13339 20683 13345
rect 21266 13336 21272 13348
rect 21324 13336 21330 13388
rect 18049 13311 18107 13317
rect 18049 13308 18061 13311
rect 16356 13280 18061 13308
rect 16356 13268 16362 13280
rect 18049 13277 18061 13280
rect 18095 13277 18107 13311
rect 18049 13271 18107 13277
rect 18601 13311 18659 13317
rect 18601 13277 18613 13311
rect 18647 13277 18659 13311
rect 20898 13308 20904 13320
rect 20859 13280 20904 13308
rect 18601 13271 18659 13277
rect 20898 13268 20904 13280
rect 20956 13268 20962 13320
rect 5353 13243 5411 13249
rect 5353 13209 5365 13243
rect 5399 13240 5411 13243
rect 5399 13212 6132 13240
rect 5399 13209 5411 13212
rect 5353 13203 5411 13209
rect 5718 13172 5724 13184
rect 5679 13144 5724 13172
rect 5718 13132 5724 13144
rect 5776 13132 5782 13184
rect 6104 13181 6132 13212
rect 8386 13200 8392 13252
rect 8444 13240 8450 13252
rect 9278 13243 9336 13249
rect 9278 13240 9290 13243
rect 8444 13212 9290 13240
rect 8444 13200 8450 13212
rect 9278 13209 9290 13212
rect 9324 13209 9336 13243
rect 11824 13243 11882 13249
rect 11824 13240 11836 13243
rect 9278 13203 9336 13209
rect 10428 13212 11836 13240
rect 10428 13184 10456 13212
rect 11824 13209 11836 13212
rect 11870 13240 11882 13243
rect 13078 13240 13084 13252
rect 11870 13212 13084 13240
rect 11870 13209 11882 13212
rect 11824 13203 11882 13209
rect 13078 13200 13084 13212
rect 13136 13200 13142 13252
rect 13480 13243 13538 13249
rect 13480 13209 13492 13243
rect 13526 13240 13538 13243
rect 15010 13240 15016 13252
rect 13526 13212 15016 13240
rect 13526 13209 13538 13212
rect 13480 13203 13538 13209
rect 15010 13200 15016 13212
rect 15068 13200 15074 13252
rect 16022 13240 16028 13252
rect 15120 13212 16028 13240
rect 6089 13175 6147 13181
rect 6089 13141 6101 13175
rect 6135 13172 6147 13175
rect 6822 13172 6828 13184
rect 6135 13144 6828 13172
rect 6135 13141 6147 13144
rect 6089 13135 6147 13141
rect 6822 13132 6828 13144
rect 6880 13132 6886 13184
rect 7834 13132 7840 13184
rect 7892 13172 7898 13184
rect 9674 13172 9680 13184
rect 7892 13144 9680 13172
rect 7892 13132 7898 13144
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 10410 13172 10416 13184
rect 10323 13144 10416 13172
rect 10410 13132 10416 13144
rect 10468 13132 10474 13184
rect 13998 13132 14004 13184
rect 14056 13172 14062 13184
rect 14093 13175 14151 13181
rect 14093 13172 14105 13175
rect 14056 13144 14105 13172
rect 14056 13132 14062 13144
rect 14093 13141 14105 13144
rect 14139 13141 14151 13175
rect 14093 13135 14151 13141
rect 14274 13132 14280 13184
rect 14332 13172 14338 13184
rect 15120 13172 15148 13212
rect 16022 13200 16028 13212
rect 16080 13200 16086 13252
rect 16476 13243 16534 13249
rect 16476 13209 16488 13243
rect 16522 13240 16534 13243
rect 17034 13240 17040 13252
rect 16522 13212 17040 13240
rect 16522 13209 16534 13212
rect 16476 13203 16534 13209
rect 17034 13200 17040 13212
rect 17092 13200 17098 13252
rect 20358 13243 20416 13249
rect 20358 13240 20370 13243
rect 17604 13212 20370 13240
rect 14332 13144 15148 13172
rect 14332 13132 14338 13144
rect 15838 13132 15844 13184
rect 15896 13172 15902 13184
rect 17604 13181 17632 13212
rect 20358 13209 20370 13212
rect 20404 13209 20416 13243
rect 20358 13203 20416 13209
rect 17589 13175 17647 13181
rect 17589 13172 17601 13175
rect 15896 13144 17601 13172
rect 15896 13132 15902 13144
rect 17589 13141 17601 13144
rect 17635 13141 17647 13175
rect 17589 13135 17647 13141
rect 22002 13132 22008 13184
rect 22060 13172 22066 13184
rect 22554 13172 22560 13184
rect 22060 13144 22560 13172
rect 22060 13132 22066 13144
rect 22554 13132 22560 13144
rect 22612 13132 22618 13184
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 5261 12971 5319 12977
rect 5261 12937 5273 12971
rect 5307 12968 5319 12971
rect 5718 12968 5724 12980
rect 5307 12940 5724 12968
rect 5307 12937 5319 12940
rect 5261 12931 5319 12937
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 7834 12968 7840 12980
rect 7795 12940 7840 12968
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 8478 12928 8484 12980
rect 8536 12968 8542 12980
rect 17218 12968 17224 12980
rect 8536 12940 17224 12968
rect 8536 12928 8542 12940
rect 17218 12928 17224 12940
rect 17276 12928 17282 12980
rect 5350 12900 5356 12912
rect 5311 12872 5356 12900
rect 5350 12860 5356 12872
rect 5408 12860 5414 12912
rect 8294 12900 8300 12912
rect 6564 12872 8300 12900
rect 6564 12844 6592 12872
rect 8128 12844 8156 12872
rect 8294 12860 8300 12872
rect 8352 12900 8358 12912
rect 11054 12900 11060 12912
rect 8352 12872 11060 12900
rect 8352 12860 8358 12872
rect 5718 12792 5724 12844
rect 5776 12832 5782 12844
rect 5902 12832 5908 12844
rect 5776 12804 5908 12832
rect 5776 12792 5782 12804
rect 5902 12792 5908 12804
rect 5960 12792 5966 12844
rect 6457 12835 6515 12841
rect 6457 12801 6469 12835
rect 6503 12832 6515 12835
rect 6546 12832 6552 12844
rect 6503 12804 6552 12832
rect 6503 12801 6515 12804
rect 6457 12795 6515 12801
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 6730 12841 6736 12844
rect 6724 12832 6736 12841
rect 6691 12804 6736 12832
rect 6724 12795 6736 12804
rect 6730 12792 6736 12795
rect 6788 12792 6794 12844
rect 8110 12832 8116 12844
rect 8023 12804 8116 12832
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 8380 12835 8438 12841
rect 8380 12801 8392 12835
rect 8426 12832 8438 12835
rect 9306 12832 9312 12844
rect 8426 12804 9312 12832
rect 8426 12801 8438 12804
rect 8380 12795 8438 12801
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 9784 12841 9812 12872
rect 11054 12860 11060 12872
rect 11112 12900 11118 12912
rect 11517 12903 11575 12909
rect 11517 12900 11529 12903
rect 11112 12872 11529 12900
rect 11112 12860 11118 12872
rect 11517 12869 11529 12872
rect 11563 12900 11575 12903
rect 12066 12900 12072 12912
rect 11563 12872 12072 12900
rect 11563 12869 11575 12872
rect 11517 12863 11575 12869
rect 12066 12860 12072 12872
rect 12124 12900 12130 12912
rect 12161 12903 12219 12909
rect 12161 12900 12173 12903
rect 12124 12872 12173 12900
rect 12124 12860 12130 12872
rect 12161 12869 12173 12872
rect 12207 12900 12219 12903
rect 12529 12903 12587 12909
rect 12529 12900 12541 12903
rect 12207 12872 12541 12900
rect 12207 12869 12219 12872
rect 12161 12863 12219 12869
rect 12529 12869 12541 12872
rect 12575 12900 12587 12903
rect 12710 12900 12716 12912
rect 12575 12872 12716 12900
rect 12575 12869 12587 12872
rect 12529 12863 12587 12869
rect 12710 12860 12716 12872
rect 12768 12900 12774 12912
rect 15470 12900 15476 12912
rect 12768 12872 15476 12900
rect 12768 12860 12774 12872
rect 9769 12835 9827 12841
rect 9769 12801 9781 12835
rect 9815 12801 9827 12835
rect 10036 12835 10094 12841
rect 10036 12832 10048 12835
rect 9769 12795 9827 12801
rect 9876 12804 10048 12832
rect 4982 12724 4988 12776
rect 5040 12764 5046 12776
rect 5077 12767 5135 12773
rect 5077 12764 5089 12767
rect 5040 12736 5089 12764
rect 5040 12724 5046 12736
rect 5077 12733 5089 12736
rect 5123 12733 5135 12767
rect 9876 12764 9904 12804
rect 10036 12801 10048 12804
rect 10082 12832 10094 12835
rect 11974 12832 11980 12844
rect 10082 12804 11980 12832
rect 10082 12801 10094 12804
rect 10036 12795 10094 12801
rect 11974 12792 11980 12804
rect 12032 12792 12038 12844
rect 12250 12792 12256 12844
rect 12308 12832 12314 12844
rect 13998 12832 14004 12844
rect 14056 12841 14062 12844
rect 14292 12841 14320 12872
rect 15470 12860 15476 12872
rect 15528 12900 15534 12912
rect 16209 12903 16267 12909
rect 16209 12900 16221 12903
rect 15528 12872 16221 12900
rect 15528 12860 15534 12872
rect 12308 12804 14004 12832
rect 12308 12792 12314 12804
rect 13998 12792 14004 12804
rect 14056 12795 14068 12841
rect 14277 12835 14335 12841
rect 14277 12801 14289 12835
rect 14323 12801 14335 12835
rect 14277 12795 14335 12801
rect 14056 12792 14062 12795
rect 14642 12792 14648 12844
rect 14700 12832 14706 12844
rect 14826 12832 14832 12844
rect 14700 12804 14832 12832
rect 14700 12792 14706 12804
rect 14826 12792 14832 12804
rect 14884 12832 14890 12844
rect 15948 12841 15976 12872
rect 16209 12869 16221 12872
rect 16255 12869 16267 12903
rect 16209 12863 16267 12869
rect 18690 12860 18696 12912
rect 18748 12900 18754 12912
rect 20162 12900 20168 12912
rect 18748 12872 20168 12900
rect 18748 12860 18754 12872
rect 20162 12860 20168 12872
rect 20220 12860 20226 12912
rect 21116 12903 21174 12909
rect 21116 12869 21128 12903
rect 21162 12900 21174 12903
rect 21634 12900 21640 12912
rect 21162 12872 21640 12900
rect 21162 12869 21174 12872
rect 21116 12863 21174 12869
rect 21634 12860 21640 12872
rect 21692 12860 21698 12912
rect 15666 12835 15724 12841
rect 15666 12832 15678 12835
rect 14884 12804 15678 12832
rect 14884 12792 14890 12804
rect 15666 12801 15678 12804
rect 15712 12801 15724 12835
rect 15666 12795 15724 12801
rect 15933 12835 15991 12841
rect 15933 12801 15945 12835
rect 15979 12801 15991 12835
rect 15933 12795 15991 12801
rect 16114 12792 16120 12844
rect 16172 12832 16178 12844
rect 17782 12835 17840 12841
rect 17782 12832 17794 12835
rect 16172 12804 17794 12832
rect 16172 12792 16178 12804
rect 17782 12801 17794 12804
rect 17828 12801 17840 12835
rect 17782 12795 17840 12801
rect 18592 12835 18650 12841
rect 18592 12801 18604 12835
rect 18638 12832 18650 12835
rect 19702 12832 19708 12844
rect 18638 12804 19708 12832
rect 18638 12801 18650 12804
rect 18592 12795 18650 12801
rect 19702 12792 19708 12804
rect 19760 12792 19766 12844
rect 21266 12792 21272 12844
rect 21324 12832 21330 12844
rect 21361 12835 21419 12841
rect 21361 12832 21373 12835
rect 21324 12804 21373 12832
rect 21324 12792 21330 12804
rect 21361 12801 21373 12804
rect 21407 12801 21419 12835
rect 21361 12795 21419 12801
rect 5077 12727 5135 12733
rect 9508 12736 9904 12764
rect 9508 12705 9536 12736
rect 10870 12724 10876 12776
rect 10928 12764 10934 12776
rect 18046 12764 18052 12776
rect 10928 12736 12940 12764
rect 18007 12736 18052 12764
rect 10928 12724 10934 12736
rect 12912 12705 12940 12736
rect 18046 12724 18052 12736
rect 18104 12764 18110 12776
rect 18325 12767 18383 12773
rect 18325 12764 18337 12767
rect 18104 12736 18337 12764
rect 18104 12724 18110 12736
rect 18325 12733 18337 12736
rect 18371 12733 18383 12767
rect 18325 12727 18383 12733
rect 9493 12699 9551 12705
rect 7760 12668 8156 12696
rect 5721 12631 5779 12637
rect 5721 12597 5733 12631
rect 5767 12628 5779 12631
rect 7760 12628 7788 12668
rect 5767 12600 7788 12628
rect 8128 12628 8156 12668
rect 9493 12665 9505 12699
rect 9539 12665 9551 12699
rect 9493 12659 9551 12665
rect 12897 12699 12955 12705
rect 12897 12665 12909 12699
rect 12943 12665 12955 12699
rect 12897 12659 12955 12665
rect 16022 12656 16028 12708
rect 16080 12696 16086 12708
rect 16669 12699 16727 12705
rect 16669 12696 16681 12699
rect 16080 12668 16681 12696
rect 16080 12656 16086 12668
rect 16669 12665 16681 12668
rect 16715 12665 16727 12699
rect 19981 12699 20039 12705
rect 19981 12696 19993 12699
rect 16669 12659 16727 12665
rect 19260 12668 19993 12696
rect 8478 12628 8484 12640
rect 8128 12600 8484 12628
rect 5767 12597 5779 12600
rect 5721 12591 5779 12597
rect 8478 12588 8484 12600
rect 8536 12588 8542 12640
rect 9030 12588 9036 12640
rect 9088 12628 9094 12640
rect 9214 12628 9220 12640
rect 9088 12600 9220 12628
rect 9088 12588 9094 12600
rect 9214 12588 9220 12600
rect 9272 12588 9278 12640
rect 11146 12628 11152 12640
rect 11107 12600 11152 12628
rect 11146 12588 11152 12600
rect 11204 12588 11210 12640
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 14274 12628 14280 12640
rect 11848 12600 14280 12628
rect 11848 12588 11854 12600
rect 14274 12588 14280 12600
rect 14332 12588 14338 12640
rect 14550 12628 14556 12640
rect 14511 12600 14556 12628
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 18690 12588 18696 12640
rect 18748 12628 18754 12640
rect 19260 12628 19288 12668
rect 19981 12665 19993 12668
rect 20027 12665 20039 12699
rect 19981 12659 20039 12665
rect 18748 12600 19288 12628
rect 19705 12631 19763 12637
rect 18748 12588 18754 12600
rect 19705 12597 19717 12631
rect 19751 12628 19763 12631
rect 19886 12628 19892 12640
rect 19751 12600 19892 12628
rect 19751 12597 19763 12600
rect 19705 12591 19763 12597
rect 19886 12588 19892 12600
rect 19944 12588 19950 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 10410 12424 10416 12436
rect 6840 12396 10416 12424
rect 5445 12291 5503 12297
rect 5445 12257 5457 12291
rect 5491 12288 5503 12291
rect 6730 12288 6736 12300
rect 5491 12260 6736 12288
rect 5491 12257 5503 12260
rect 5445 12251 5503 12257
rect 6730 12248 6736 12260
rect 6788 12248 6794 12300
rect 6840 12297 6868 12396
rect 10410 12384 10416 12396
rect 10468 12384 10474 12436
rect 12710 12384 12716 12436
rect 12768 12424 12774 12436
rect 12897 12427 12955 12433
rect 12897 12424 12909 12427
rect 12768 12396 12909 12424
rect 12768 12384 12774 12396
rect 12897 12393 12909 12396
rect 12943 12424 12955 12427
rect 13265 12427 13323 12433
rect 13265 12424 13277 12427
rect 12943 12396 13277 12424
rect 12943 12393 12955 12396
rect 12897 12387 12955 12393
rect 13265 12393 13277 12396
rect 13311 12424 13323 12427
rect 13633 12427 13691 12433
rect 13633 12424 13645 12427
rect 13311 12396 13645 12424
rect 13311 12393 13323 12396
rect 13265 12387 13323 12393
rect 13633 12393 13645 12396
rect 13679 12393 13691 12427
rect 13633 12387 13691 12393
rect 14093 12427 14151 12433
rect 14093 12393 14105 12427
rect 14139 12424 14151 12427
rect 14139 12396 15516 12424
rect 14139 12393 14151 12396
rect 14093 12387 14151 12393
rect 9030 12356 9036 12368
rect 8404 12328 9036 12356
rect 6825 12291 6883 12297
rect 6825 12257 6837 12291
rect 6871 12257 6883 12291
rect 6825 12251 6883 12257
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 5994 12220 6000 12232
rect 5684 12192 6000 12220
rect 5684 12180 5690 12192
rect 5994 12180 6000 12192
rect 6052 12180 6058 12232
rect 6546 12180 6552 12232
rect 6604 12180 6610 12232
rect 7193 12223 7251 12229
rect 7193 12189 7205 12223
rect 7239 12220 7251 12223
rect 7926 12220 7932 12232
rect 7239 12192 7932 12220
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 7926 12180 7932 12192
rect 7984 12220 7990 12232
rect 8404 12220 8432 12328
rect 9030 12316 9036 12328
rect 9088 12316 9094 12368
rect 13814 12316 13820 12368
rect 13872 12356 13878 12368
rect 14108 12356 14136 12387
rect 13872 12328 14136 12356
rect 15488 12356 15516 12396
rect 16022 12384 16028 12436
rect 16080 12424 16086 12436
rect 19613 12427 19671 12433
rect 16080 12396 19472 12424
rect 16080 12384 16086 12396
rect 16114 12356 16120 12368
rect 15488 12328 16120 12356
rect 13872 12316 13878 12328
rect 16114 12316 16120 12328
rect 16172 12316 16178 12368
rect 8956 12260 9260 12288
rect 8956 12220 8984 12260
rect 7984 12192 8432 12220
rect 8496 12192 8984 12220
rect 7984 12180 7990 12192
rect 6564 12152 6592 12180
rect 6641 12155 6699 12161
rect 6641 12152 6653 12155
rect 5000 12124 6653 12152
rect 5000 12096 5028 12124
rect 6641 12121 6653 12124
rect 6687 12121 6699 12155
rect 6641 12115 6699 12121
rect 7460 12155 7518 12161
rect 7460 12121 7472 12155
rect 7506 12152 7518 12155
rect 8496 12152 8524 12192
rect 9030 12180 9036 12232
rect 9088 12220 9094 12232
rect 9125 12223 9183 12229
rect 9125 12220 9137 12223
rect 9088 12192 9137 12220
rect 9088 12180 9094 12192
rect 9125 12189 9137 12192
rect 9171 12189 9183 12223
rect 9232 12220 9260 12260
rect 10594 12248 10600 12300
rect 10652 12288 10658 12300
rect 11146 12288 11152 12300
rect 10652 12260 11152 12288
rect 10652 12248 10658 12260
rect 11146 12248 11152 12260
rect 11204 12288 11210 12300
rect 15470 12288 15476 12300
rect 11204 12260 11376 12288
rect 15431 12260 15476 12288
rect 11204 12248 11210 12260
rect 9858 12220 9864 12232
rect 9232 12192 9864 12220
rect 9125 12183 9183 12189
rect 9858 12180 9864 12192
rect 9916 12220 9922 12232
rect 10870 12220 10876 12232
rect 9916 12192 10876 12220
rect 9916 12180 9922 12192
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 11054 12180 11060 12232
rect 11112 12220 11118 12232
rect 11241 12223 11299 12229
rect 11241 12220 11253 12223
rect 11112 12192 11253 12220
rect 11112 12180 11118 12192
rect 11241 12189 11253 12192
rect 11287 12189 11299 12223
rect 11348 12220 11376 12260
rect 15470 12248 15476 12260
rect 15528 12248 15534 12300
rect 17586 12248 17592 12300
rect 17644 12288 17650 12300
rect 17770 12288 17776 12300
rect 17644 12260 17776 12288
rect 17644 12248 17650 12260
rect 17770 12248 17776 12260
rect 17828 12248 17834 12300
rect 11497 12223 11555 12229
rect 11497 12220 11509 12223
rect 11348 12192 11509 12220
rect 11241 12183 11299 12189
rect 11497 12189 11509 12192
rect 11543 12189 11555 12223
rect 15488 12220 15516 12248
rect 17034 12220 17040 12232
rect 15488 12192 17040 12220
rect 11497 12183 11555 12189
rect 17034 12180 17040 12192
rect 17092 12220 17098 12232
rect 17129 12223 17187 12229
rect 17129 12220 17141 12223
rect 17092 12192 17141 12220
rect 17092 12180 17098 12192
rect 17129 12189 17141 12192
rect 17175 12189 17187 12223
rect 17129 12183 17187 12189
rect 18046 12180 18052 12232
rect 18104 12220 18110 12232
rect 18785 12223 18843 12229
rect 18785 12220 18797 12223
rect 18104 12192 18797 12220
rect 18104 12180 18110 12192
rect 18785 12189 18797 12192
rect 18831 12189 18843 12223
rect 18785 12183 18843 12189
rect 19058 12180 19064 12232
rect 19116 12180 19122 12232
rect 19444 12229 19472 12396
rect 19613 12393 19625 12427
rect 19659 12424 19671 12427
rect 20438 12424 20444 12436
rect 19659 12396 20444 12424
rect 19659 12393 19671 12396
rect 19613 12387 19671 12393
rect 20438 12384 20444 12396
rect 20496 12384 20502 12436
rect 19429 12223 19487 12229
rect 19429 12189 19441 12223
rect 19475 12189 19487 12223
rect 19429 12183 19487 12189
rect 21266 12180 21272 12232
rect 21324 12220 21330 12232
rect 21361 12223 21419 12229
rect 21361 12220 21373 12223
rect 21324 12192 21373 12220
rect 21324 12180 21330 12192
rect 21361 12189 21373 12192
rect 21407 12189 21419 12223
rect 21361 12183 21419 12189
rect 9392 12155 9450 12161
rect 9392 12152 9404 12155
rect 7506 12124 8524 12152
rect 8588 12124 9404 12152
rect 7506 12121 7518 12124
rect 7460 12115 7518 12121
rect 4982 12084 4988 12096
rect 4943 12056 4988 12084
rect 4982 12044 4988 12056
rect 5040 12044 5046 12096
rect 5902 12084 5908 12096
rect 5863 12056 5908 12084
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 5994 12044 6000 12096
rect 6052 12084 6058 12096
rect 6181 12087 6239 12093
rect 6181 12084 6193 12087
rect 6052 12056 6193 12084
rect 6052 12044 6058 12056
rect 6181 12053 6193 12056
rect 6227 12053 6239 12087
rect 6181 12047 6239 12053
rect 6549 12087 6607 12093
rect 6549 12053 6561 12087
rect 6595 12084 6607 12087
rect 6730 12084 6736 12096
rect 6595 12056 6736 12084
rect 6595 12053 6607 12056
rect 6549 12047 6607 12053
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 7190 12044 7196 12096
rect 7248 12084 7254 12096
rect 7650 12084 7656 12096
rect 7248 12056 7656 12084
rect 7248 12044 7254 12056
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 8588 12093 8616 12124
rect 9392 12121 9404 12124
rect 9438 12152 9450 12155
rect 9674 12152 9680 12164
rect 9438 12124 9680 12152
rect 9438 12121 9450 12124
rect 9392 12115 9450 12121
rect 9674 12112 9680 12124
rect 9732 12112 9738 12164
rect 10318 12112 10324 12164
rect 10376 12152 10382 12164
rect 12986 12152 12992 12164
rect 10376 12124 12992 12152
rect 10376 12112 10382 12124
rect 8573 12087 8631 12093
rect 8573 12053 8585 12087
rect 8619 12053 8631 12087
rect 8573 12047 8631 12053
rect 9122 12044 9128 12096
rect 9180 12084 9186 12096
rect 9490 12084 9496 12096
rect 9180 12056 9496 12084
rect 9180 12044 9186 12056
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 10520 12093 10548 12124
rect 12986 12112 12992 12124
rect 13044 12112 13050 12164
rect 15228 12155 15286 12161
rect 15228 12121 15240 12155
rect 15274 12152 15286 12155
rect 15562 12152 15568 12164
rect 15274 12124 15568 12152
rect 15274 12121 15286 12124
rect 15228 12115 15286 12121
rect 15562 12112 15568 12124
rect 15620 12152 15626 12164
rect 16942 12161 16948 12164
rect 16884 12155 16948 12161
rect 16884 12152 16896 12155
rect 15620 12124 15884 12152
rect 16855 12124 16896 12152
rect 15620 12112 15626 12124
rect 10505 12087 10563 12093
rect 10505 12053 10517 12087
rect 10551 12053 10563 12087
rect 10505 12047 10563 12053
rect 10873 12087 10931 12093
rect 10873 12053 10885 12087
rect 10919 12084 10931 12087
rect 11146 12084 11152 12096
rect 10919 12056 11152 12084
rect 10919 12053 10931 12056
rect 10873 12047 10931 12053
rect 11146 12044 11152 12056
rect 11204 12044 11210 12096
rect 12526 12044 12532 12096
rect 12584 12084 12590 12096
rect 12621 12087 12679 12093
rect 12621 12084 12633 12087
rect 12584 12056 12633 12084
rect 12584 12044 12590 12056
rect 12621 12053 12633 12056
rect 12667 12084 12679 12087
rect 12710 12084 12716 12096
rect 12667 12056 12716 12084
rect 12667 12053 12679 12056
rect 12621 12047 12679 12053
rect 12710 12044 12716 12056
rect 12768 12044 12774 12096
rect 14918 12044 14924 12096
rect 14976 12084 14982 12096
rect 15749 12087 15807 12093
rect 15749 12084 15761 12087
rect 14976 12056 15761 12084
rect 14976 12044 14982 12056
rect 15749 12053 15761 12056
rect 15795 12053 15807 12087
rect 15856 12084 15884 12124
rect 16884 12121 16896 12124
rect 16930 12121 16948 12155
rect 16884 12115 16948 12121
rect 16942 12112 16948 12115
rect 17000 12152 17006 12164
rect 17586 12152 17592 12164
rect 17000 12124 17592 12152
rect 17000 12112 17006 12124
rect 17586 12112 17592 12124
rect 17644 12112 17650 12164
rect 17954 12112 17960 12164
rect 18012 12152 18018 12164
rect 18138 12152 18144 12164
rect 18012 12124 18144 12152
rect 18012 12112 18018 12124
rect 18138 12112 18144 12124
rect 18196 12112 18202 12164
rect 18540 12155 18598 12161
rect 18540 12121 18552 12155
rect 18586 12152 18598 12155
rect 19076 12152 19104 12180
rect 18586 12124 19104 12152
rect 21116 12155 21174 12161
rect 18586 12121 18598 12124
rect 18540 12115 18598 12121
rect 18800 12096 18828 12124
rect 21116 12121 21128 12155
rect 21162 12152 21174 12155
rect 21542 12152 21548 12164
rect 21162 12124 21548 12152
rect 21162 12121 21174 12124
rect 21116 12115 21174 12121
rect 21542 12112 21548 12124
rect 21600 12152 21606 12164
rect 22094 12152 22100 12164
rect 21600 12124 22100 12152
rect 21600 12112 21606 12124
rect 22094 12112 22100 12124
rect 22152 12112 22158 12164
rect 17405 12087 17463 12093
rect 17405 12084 17417 12087
rect 15856 12056 17417 12084
rect 15749 12047 15807 12053
rect 17405 12053 17417 12056
rect 17451 12053 17463 12087
rect 17405 12047 17463 12053
rect 18782 12044 18788 12096
rect 18840 12044 18846 12096
rect 19058 12044 19064 12096
rect 19116 12084 19122 12096
rect 19518 12084 19524 12096
rect 19116 12056 19524 12084
rect 19116 12044 19122 12056
rect 19518 12044 19524 12056
rect 19576 12084 19582 12096
rect 19981 12087 20039 12093
rect 19981 12084 19993 12087
rect 19576 12056 19993 12084
rect 19576 12044 19582 12056
rect 19981 12053 19993 12056
rect 20027 12053 20039 12087
rect 19981 12047 20039 12053
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 6454 11840 6460 11892
rect 6512 11880 6518 11892
rect 6822 11880 6828 11892
rect 6512 11852 6828 11880
rect 6512 11840 6518 11852
rect 6822 11840 6828 11852
rect 6880 11840 6886 11892
rect 7006 11880 7012 11892
rect 6967 11852 7012 11880
rect 7006 11840 7012 11852
rect 7064 11840 7070 11892
rect 7469 11883 7527 11889
rect 7469 11849 7481 11883
rect 7515 11880 7527 11883
rect 8018 11880 8024 11892
rect 7515 11852 8024 11880
rect 7515 11849 7527 11852
rect 7469 11843 7527 11849
rect 8018 11840 8024 11852
rect 8076 11840 8082 11892
rect 8113 11883 8171 11889
rect 8113 11849 8125 11883
rect 8159 11880 8171 11883
rect 8202 11880 8208 11892
rect 8159 11852 8208 11880
rect 8159 11849 8171 11852
rect 8113 11843 8171 11849
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 12894 11880 12900 11892
rect 9180 11852 12434 11880
rect 12855 11852 12900 11880
rect 9180 11840 9186 11852
rect 6733 11815 6791 11821
rect 6733 11781 6745 11815
rect 6779 11812 6791 11815
rect 8481 11815 8539 11821
rect 8481 11812 8493 11815
rect 6779 11784 8493 11812
rect 6779 11781 6791 11784
rect 6733 11775 6791 11781
rect 8481 11781 8493 11784
rect 8527 11781 8539 11815
rect 11054 11812 11060 11824
rect 8481 11775 8539 11781
rect 9600 11784 11060 11812
rect 5166 11704 5172 11756
rect 5224 11744 5230 11756
rect 5537 11747 5595 11753
rect 5537 11744 5549 11747
rect 5224 11716 5549 11744
rect 5224 11704 5230 11716
rect 5537 11713 5549 11716
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 5629 11747 5687 11753
rect 5629 11713 5641 11747
rect 5675 11744 5687 11747
rect 6086 11744 6092 11756
rect 5675 11716 6092 11744
rect 5675 11713 5687 11716
rect 5629 11707 5687 11713
rect 6086 11704 6092 11716
rect 6144 11704 6150 11756
rect 6822 11704 6828 11756
rect 6880 11744 6886 11756
rect 7098 11744 7104 11756
rect 6880 11716 7104 11744
rect 6880 11704 6886 11716
rect 7098 11704 7104 11716
rect 7156 11704 7162 11756
rect 7377 11747 7435 11753
rect 7377 11713 7389 11747
rect 7423 11744 7435 11747
rect 7834 11744 7840 11756
rect 7423 11716 7840 11744
rect 7423 11713 7435 11716
rect 7377 11707 7435 11713
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 5445 11679 5503 11685
rect 5445 11645 5457 11679
rect 5491 11645 5503 11679
rect 5445 11639 5503 11645
rect 7653 11679 7711 11685
rect 7653 11645 7665 11679
rect 7699 11676 7711 11679
rect 8386 11676 8392 11688
rect 7699 11648 8392 11676
rect 7699 11645 7711 11648
rect 7653 11639 7711 11645
rect 5460 11608 5488 11639
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 8570 11676 8576 11688
rect 8531 11648 8576 11676
rect 8570 11636 8576 11648
rect 8628 11636 8634 11688
rect 8757 11679 8815 11685
rect 8757 11645 8769 11679
rect 8803 11676 8815 11679
rect 9600 11676 9628 11784
rect 11054 11772 11060 11784
rect 11112 11772 11118 11824
rect 11238 11772 11244 11824
rect 11296 11812 11302 11824
rect 12253 11815 12311 11821
rect 12253 11812 12265 11815
rect 11296 11784 12265 11812
rect 11296 11772 11302 11784
rect 12253 11781 12265 11784
rect 12299 11781 12311 11815
rect 12406 11812 12434 11852
rect 12894 11840 12900 11852
rect 12952 11840 12958 11892
rect 14366 11880 14372 11892
rect 13004 11852 13216 11880
rect 14327 11852 14372 11880
rect 13004 11812 13032 11852
rect 12406 11784 13032 11812
rect 13188 11812 13216 11852
rect 14366 11840 14372 11852
rect 14424 11840 14430 11892
rect 14734 11840 14740 11892
rect 14792 11880 14798 11892
rect 14918 11880 14924 11892
rect 14792 11852 14924 11880
rect 14792 11840 14798 11852
rect 14918 11840 14924 11852
rect 14976 11840 14982 11892
rect 15470 11840 15476 11892
rect 15528 11880 15534 11892
rect 15565 11883 15623 11889
rect 15565 11880 15577 11883
rect 15528 11852 15577 11880
rect 15528 11840 15534 11852
rect 15565 11849 15577 11852
rect 15611 11849 15623 11883
rect 15565 11843 15623 11849
rect 16114 11840 16120 11892
rect 16172 11880 16178 11892
rect 16301 11883 16359 11889
rect 16301 11880 16313 11883
rect 16172 11852 16313 11880
rect 16172 11840 16178 11852
rect 16301 11849 16313 11852
rect 16347 11880 16359 11883
rect 16942 11880 16948 11892
rect 16347 11852 16948 11880
rect 16347 11849 16359 11852
rect 16301 11843 16359 11849
rect 16942 11840 16948 11852
rect 17000 11840 17006 11892
rect 17862 11840 17868 11892
rect 17920 11880 17926 11892
rect 18690 11880 18696 11892
rect 17920 11852 18696 11880
rect 17920 11840 17926 11852
rect 15746 11812 15752 11824
rect 13188 11784 15752 11812
rect 12253 11775 12311 11781
rect 15746 11772 15752 11784
rect 15804 11772 15810 11824
rect 17034 11772 17040 11824
rect 17092 11812 17098 11824
rect 18046 11812 18052 11824
rect 17092 11784 18052 11812
rect 17092 11772 17098 11784
rect 10341 11747 10399 11753
rect 10341 11713 10353 11747
rect 10387 11744 10399 11747
rect 11790 11744 11796 11756
rect 10387 11716 11796 11744
rect 10387 11713 10399 11716
rect 10341 11707 10399 11713
rect 11790 11704 11796 11716
rect 11848 11704 11854 11756
rect 11882 11704 11888 11756
rect 11940 11744 11946 11756
rect 13265 11747 13323 11753
rect 11940 11716 11985 11744
rect 11940 11704 11946 11716
rect 13265 11713 13277 11747
rect 13311 11744 13323 11747
rect 14366 11744 14372 11756
rect 13311 11716 14372 11744
rect 13311 11713 13323 11716
rect 13265 11707 13323 11713
rect 14366 11704 14372 11716
rect 14424 11704 14430 11756
rect 14737 11747 14795 11753
rect 14737 11713 14749 11747
rect 14783 11744 14795 11747
rect 15194 11744 15200 11756
rect 14783 11716 15200 11744
rect 14783 11713 14795 11716
rect 14737 11707 14795 11713
rect 15194 11704 15200 11716
rect 15252 11704 15258 11756
rect 17218 11744 17224 11756
rect 17179 11716 17224 11744
rect 17218 11704 17224 11716
rect 17276 11704 17282 11756
rect 17972 11753 18000 11784
rect 18046 11772 18052 11784
rect 18104 11772 18110 11824
rect 18248 11821 18276 11852
rect 18690 11840 18696 11852
rect 18748 11840 18754 11892
rect 20898 11880 20904 11892
rect 19168 11852 20904 11880
rect 18224 11815 18282 11821
rect 18224 11781 18236 11815
rect 18270 11781 18282 11815
rect 18224 11775 18282 11781
rect 17957 11747 18015 11753
rect 17957 11713 17969 11747
rect 18003 11713 18015 11747
rect 19168 11744 19196 11852
rect 20898 11840 20904 11852
rect 20956 11840 20962 11892
rect 21266 11812 21272 11824
rect 19996 11784 21272 11812
rect 19996 11753 20024 11784
rect 21266 11772 21272 11784
rect 21324 11772 21330 11824
rect 17957 11707 18015 11713
rect 18064 11716 19196 11744
rect 19705 11747 19763 11753
rect 8803 11648 9628 11676
rect 10597 11679 10655 11685
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 10597 11645 10609 11679
rect 10643 11676 10655 11679
rect 10643 11648 11008 11676
rect 10643 11645 10655 11648
rect 10597 11639 10655 11645
rect 5460 11580 9674 11608
rect 4985 11543 5043 11549
rect 4985 11509 4997 11543
rect 5031 11540 5043 11543
rect 5166 11540 5172 11552
rect 5031 11512 5172 11540
rect 5031 11509 5043 11512
rect 4985 11503 5043 11509
rect 5166 11500 5172 11512
rect 5224 11500 5230 11552
rect 5997 11543 6055 11549
rect 5997 11509 6009 11543
rect 6043 11540 6055 11543
rect 7098 11540 7104 11552
rect 6043 11512 7104 11540
rect 6043 11509 6055 11512
rect 5997 11503 6055 11509
rect 7098 11500 7104 11512
rect 7156 11500 7162 11552
rect 8478 11500 8484 11552
rect 8536 11540 8542 11552
rect 8754 11540 8760 11552
rect 8536 11512 8760 11540
rect 8536 11500 8542 11512
rect 8754 11500 8760 11512
rect 8812 11500 8818 11552
rect 9217 11543 9275 11549
rect 9217 11509 9229 11543
rect 9263 11540 9275 11543
rect 9306 11540 9312 11552
rect 9263 11512 9312 11540
rect 9263 11509 9275 11512
rect 9217 11503 9275 11509
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 9646 11540 9674 11580
rect 10870 11540 10876 11552
rect 9646 11512 10876 11540
rect 10870 11500 10876 11512
rect 10928 11500 10934 11552
rect 10980 11549 11008 11648
rect 11330 11636 11336 11688
rect 11388 11676 11394 11688
rect 11900 11676 11928 11704
rect 11388 11648 11928 11676
rect 11388 11636 11394 11648
rect 12158 11636 12164 11688
rect 12216 11676 12222 11688
rect 13357 11679 13415 11685
rect 13357 11676 13369 11679
rect 12216 11648 13369 11676
rect 12216 11636 12222 11648
rect 13357 11645 13369 11648
rect 13403 11645 13415 11679
rect 13357 11639 13415 11645
rect 13449 11679 13507 11685
rect 13449 11645 13461 11679
rect 13495 11645 13507 11679
rect 14826 11676 14832 11688
rect 14787 11648 14832 11676
rect 13449 11639 13507 11645
rect 11054 11568 11060 11620
rect 11112 11608 11118 11620
rect 11112 11580 12434 11608
rect 11112 11568 11118 11580
rect 10965 11543 11023 11549
rect 10965 11509 10977 11543
rect 11011 11540 11023 11543
rect 11146 11540 11152 11552
rect 11011 11512 11152 11540
rect 11011 11509 11023 11512
rect 10965 11503 11023 11509
rect 11146 11500 11152 11512
rect 11204 11540 11210 11552
rect 11609 11543 11667 11549
rect 11609 11540 11621 11543
rect 11204 11512 11621 11540
rect 11204 11500 11210 11512
rect 11609 11509 11621 11512
rect 11655 11540 11667 11543
rect 11698 11540 11704 11552
rect 11655 11512 11704 11540
rect 11655 11509 11667 11512
rect 11609 11503 11667 11509
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 12406 11540 12434 11580
rect 12618 11568 12624 11620
rect 12676 11608 12682 11620
rect 13464 11608 13492 11639
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 15013 11679 15071 11685
rect 15013 11645 15025 11679
rect 15059 11676 15071 11679
rect 16942 11676 16948 11688
rect 15059 11648 16344 11676
rect 16903 11648 16948 11676
rect 15059 11645 15071 11648
rect 15013 11639 15071 11645
rect 15028 11608 15056 11639
rect 12676 11580 13492 11608
rect 13556 11580 15056 11608
rect 12676 11568 12682 11580
rect 13556 11540 13584 11580
rect 12406 11512 13584 11540
rect 13630 11500 13636 11552
rect 13688 11540 13694 11552
rect 13909 11543 13967 11549
rect 13909 11540 13921 11543
rect 13688 11512 13921 11540
rect 13688 11500 13694 11512
rect 13909 11509 13921 11512
rect 13955 11509 13967 11543
rect 16316 11540 16344 11648
rect 16942 11636 16948 11648
rect 17000 11636 17006 11688
rect 17497 11679 17555 11685
rect 17497 11645 17509 11679
rect 17543 11676 17555 11679
rect 18064 11676 18092 11716
rect 19705 11713 19717 11747
rect 19751 11744 19763 11747
rect 19981 11747 20039 11753
rect 19981 11744 19993 11747
rect 19751 11716 19993 11744
rect 19751 11713 19763 11716
rect 19705 11707 19763 11713
rect 19981 11713 19993 11716
rect 20027 11713 20039 11747
rect 20237 11747 20295 11753
rect 20237 11744 20249 11747
rect 19981 11707 20039 11713
rect 20088 11716 20249 11744
rect 17543 11648 18092 11676
rect 17543 11645 17555 11648
rect 17497 11639 17555 11645
rect 19886 11636 19892 11688
rect 19944 11676 19950 11688
rect 20088 11676 20116 11716
rect 20237 11713 20249 11716
rect 20283 11713 20295 11747
rect 20237 11707 20295 11713
rect 19944 11648 20116 11676
rect 19944 11636 19950 11648
rect 21542 11608 21548 11620
rect 20916 11580 21548 11608
rect 18138 11540 18144 11552
rect 16316 11512 18144 11540
rect 13909 11503 13967 11509
rect 18138 11500 18144 11512
rect 18196 11500 18202 11552
rect 19337 11543 19395 11549
rect 19337 11509 19349 11543
rect 19383 11540 19395 11543
rect 19702 11540 19708 11552
rect 19383 11512 19708 11540
rect 19383 11509 19395 11512
rect 19337 11503 19395 11509
rect 19702 11500 19708 11512
rect 19760 11540 19766 11552
rect 20916 11540 20944 11580
rect 21542 11568 21548 11580
rect 21600 11568 21606 11620
rect 19760 11512 20944 11540
rect 19760 11500 19766 11512
rect 21082 11500 21088 11552
rect 21140 11540 21146 11552
rect 21361 11543 21419 11549
rect 21361 11540 21373 11543
rect 21140 11512 21373 11540
rect 21140 11500 21146 11512
rect 21361 11509 21373 11512
rect 21407 11509 21419 11543
rect 21361 11503 21419 11509
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 5537 11339 5595 11345
rect 5537 11305 5549 11339
rect 5583 11336 5595 11339
rect 6086 11336 6092 11348
rect 5583 11308 6092 11336
rect 5583 11305 5595 11308
rect 5537 11299 5595 11305
rect 6086 11296 6092 11308
rect 6144 11296 6150 11348
rect 6549 11339 6607 11345
rect 6549 11305 6561 11339
rect 6595 11336 6607 11339
rect 7282 11336 7288 11348
rect 6595 11308 7288 11336
rect 6595 11305 6607 11308
rect 6549 11299 6607 11305
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 7558 11336 7564 11348
rect 7519 11308 7564 11336
rect 7558 11296 7564 11308
rect 7616 11296 7622 11348
rect 7834 11336 7840 11348
rect 7795 11308 7840 11336
rect 7834 11296 7840 11308
rect 7892 11296 7898 11348
rect 8128 11308 12434 11336
rect 5905 11203 5963 11209
rect 5905 11169 5917 11203
rect 5951 11169 5963 11203
rect 5905 11163 5963 11169
rect 5920 11132 5948 11163
rect 5994 11160 6000 11212
rect 6052 11200 6058 11212
rect 6089 11203 6147 11209
rect 6089 11200 6101 11203
rect 6052 11172 6101 11200
rect 6052 11160 6058 11172
rect 6089 11169 6101 11172
rect 6135 11169 6147 11203
rect 6089 11163 6147 11169
rect 7009 11203 7067 11209
rect 7009 11169 7021 11203
rect 7055 11200 7067 11203
rect 8128 11200 8156 11308
rect 9490 11268 9496 11280
rect 9451 11240 9496 11268
rect 9490 11228 9496 11240
rect 9548 11228 9554 11280
rect 10870 11228 10876 11280
rect 10928 11268 10934 11280
rect 12158 11268 12164 11280
rect 10928 11240 11560 11268
rect 12119 11240 12164 11268
rect 10928 11228 10934 11240
rect 7055 11172 8156 11200
rect 7055 11169 7067 11172
rect 7009 11163 7067 11169
rect 8202 11160 8208 11212
rect 8260 11200 8266 11212
rect 8389 11203 8447 11209
rect 8389 11200 8401 11203
rect 8260 11172 8401 11200
rect 8260 11160 8266 11172
rect 8389 11169 8401 11172
rect 8435 11169 8447 11203
rect 11054 11200 11060 11212
rect 8389 11163 8447 11169
rect 10796 11172 11060 11200
rect 7098 11132 7104 11144
rect 5920 11104 6960 11132
rect 7059 11104 7104 11132
rect 5902 11024 5908 11076
rect 5960 11064 5966 11076
rect 6181 11067 6239 11073
rect 6181 11064 6193 11067
rect 5960 11036 6193 11064
rect 5960 11024 5966 11036
rect 6181 11033 6193 11036
rect 6227 11033 6239 11067
rect 6932 11064 6960 11104
rect 7098 11092 7104 11104
rect 7156 11092 7162 11144
rect 10796 11132 10824 11172
rect 11054 11160 11060 11172
rect 11112 11200 11118 11212
rect 11422 11200 11428 11212
rect 11112 11172 11428 11200
rect 11112 11160 11118 11172
rect 11422 11160 11428 11172
rect 11480 11160 11486 11212
rect 11532 11209 11560 11240
rect 12158 11228 12164 11240
rect 12216 11228 12222 11280
rect 12406 11268 12434 11308
rect 13446 11296 13452 11348
rect 13504 11336 13510 11348
rect 14550 11336 14556 11348
rect 13504 11308 14556 11336
rect 13504 11296 13510 11308
rect 14550 11296 14556 11308
rect 14608 11296 14614 11348
rect 14826 11296 14832 11348
rect 14884 11336 14890 11348
rect 14921 11339 14979 11345
rect 14921 11336 14933 11339
rect 14884 11308 14933 11336
rect 14884 11296 14890 11308
rect 14921 11305 14933 11308
rect 14967 11305 14979 11339
rect 15194 11336 15200 11348
rect 15155 11308 15200 11336
rect 14921 11299 14979 11305
rect 15194 11296 15200 11308
rect 15252 11296 15258 11348
rect 17034 11336 17040 11348
rect 16995 11308 17040 11336
rect 17034 11296 17040 11308
rect 17092 11296 17098 11348
rect 18414 11296 18420 11348
rect 18472 11336 18478 11348
rect 19245 11339 19303 11345
rect 19245 11336 19257 11339
rect 18472 11308 19257 11336
rect 18472 11296 18478 11308
rect 19245 11305 19257 11308
rect 19291 11305 19303 11339
rect 19245 11299 19303 11305
rect 12618 11268 12624 11280
rect 12406 11240 12624 11268
rect 12618 11228 12624 11240
rect 12676 11228 12682 11280
rect 12894 11268 12900 11280
rect 12728 11240 12900 11268
rect 11517 11203 11575 11209
rect 11517 11169 11529 11203
rect 11563 11200 11575 11203
rect 12526 11200 12532 11212
rect 11563 11172 12532 11200
rect 11563 11169 11575 11172
rect 11517 11163 11575 11169
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 8128 11104 10824 11132
rect 10873 11135 10931 11141
rect 8128 11064 8156 11104
rect 10873 11101 10885 11135
rect 10919 11132 10931 11135
rect 11146 11132 11152 11144
rect 10919 11104 11152 11132
rect 10919 11101 10931 11104
rect 10873 11095 10931 11101
rect 11146 11092 11152 11104
rect 11204 11092 11210 11144
rect 11238 11092 11244 11144
rect 11296 11132 11302 11144
rect 11701 11135 11759 11141
rect 11701 11132 11713 11135
rect 11296 11104 11713 11132
rect 11296 11092 11302 11104
rect 11701 11101 11713 11104
rect 11747 11132 11759 11135
rect 12618 11132 12624 11144
rect 11747 11104 12624 11132
rect 11747 11101 11759 11104
rect 11701 11095 11759 11101
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 6932 11036 8156 11064
rect 8205 11067 8263 11073
rect 6181 11027 6239 11033
rect 8205 11033 8217 11067
rect 8251 11064 8263 11067
rect 8941 11067 8999 11073
rect 8941 11064 8953 11067
rect 8251 11036 8953 11064
rect 8251 11033 8263 11036
rect 8205 11027 8263 11033
rect 8941 11033 8953 11036
rect 8987 11033 8999 11067
rect 8941 11027 8999 11033
rect 10617 11067 10675 11073
rect 10617 11033 10629 11067
rect 10663 11033 10675 11067
rect 11330 11064 11336 11076
rect 10617 11027 10675 11033
rect 10796 11036 11336 11064
rect 6454 10956 6460 11008
rect 6512 10996 6518 11008
rect 7006 10996 7012 11008
rect 6512 10968 7012 10996
rect 6512 10956 6518 10968
rect 7006 10956 7012 10968
rect 7064 10956 7070 11008
rect 7190 10956 7196 11008
rect 7248 10996 7254 11008
rect 8297 10999 8355 11005
rect 7248 10968 7293 10996
rect 7248 10956 7254 10968
rect 8297 10965 8309 10999
rect 8343 10996 8355 10999
rect 8386 10996 8392 11008
rect 8343 10968 8392 10996
rect 8343 10965 8355 10968
rect 8297 10959 8355 10965
rect 8386 10956 8392 10968
rect 8444 10956 8450 11008
rect 10410 10956 10416 11008
rect 10468 10996 10474 11008
rect 10643 10996 10671 11027
rect 10796 10996 10824 11036
rect 11330 11024 11336 11036
rect 11388 11024 11394 11076
rect 10468 10968 10824 10996
rect 11793 10999 11851 11005
rect 10468 10956 10474 10968
rect 11793 10965 11805 10999
rect 11839 10996 11851 10999
rect 12158 10996 12164 11008
rect 11839 10968 12164 10996
rect 11839 10965 11851 10968
rect 11793 10959 11851 10965
rect 12158 10956 12164 10968
rect 12216 10956 12222 11008
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 12728 10996 12756 11240
rect 12894 11228 12900 11240
rect 12952 11228 12958 11280
rect 13280 11240 15884 11268
rect 13078 11160 13084 11212
rect 13136 11200 13142 11212
rect 13280 11200 13308 11240
rect 13136 11172 13308 11200
rect 14369 11203 14427 11209
rect 13136 11160 13142 11172
rect 14369 11169 14381 11203
rect 14415 11200 14427 11203
rect 15746 11200 15752 11212
rect 14415 11172 15752 11200
rect 14415 11169 14427 11172
rect 14369 11163 14427 11169
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 15856 11200 15884 11240
rect 16942 11228 16948 11280
rect 17000 11268 17006 11280
rect 17000 11240 18828 11268
rect 17000 11228 17006 11240
rect 17865 11203 17923 11209
rect 17865 11200 17877 11203
rect 15856 11172 17877 11200
rect 17865 11169 17877 11172
rect 17911 11169 17923 11203
rect 18690 11200 18696 11212
rect 17865 11163 17923 11169
rect 17972 11172 18696 11200
rect 14090 11092 14096 11144
rect 14148 11132 14154 11144
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 14148 11104 14473 11132
rect 14148 11092 14154 11104
rect 14461 11101 14473 11104
rect 14507 11132 14519 11135
rect 14550 11132 14556 11144
rect 14507 11104 14556 11132
rect 14507 11101 14519 11104
rect 14461 11095 14519 11101
rect 14550 11092 14556 11104
rect 14608 11092 14614 11144
rect 14642 11092 14648 11144
rect 14700 11132 14706 11144
rect 14826 11132 14832 11144
rect 14700 11104 14832 11132
rect 14700 11092 14706 11104
rect 14826 11092 14832 11104
rect 14884 11092 14890 11144
rect 15565 11135 15623 11141
rect 15565 11101 15577 11135
rect 15611 11132 15623 11135
rect 16114 11132 16120 11144
rect 15611 11104 16120 11132
rect 15611 11101 15623 11104
rect 15565 11095 15623 11101
rect 16114 11092 16120 11104
rect 16172 11092 16178 11144
rect 16206 11092 16212 11144
rect 16264 11132 16270 11144
rect 16301 11135 16359 11141
rect 16301 11132 16313 11135
rect 16264 11104 16313 11132
rect 16264 11092 16270 11104
rect 16301 11101 16313 11104
rect 16347 11132 16359 11135
rect 17972 11132 18000 11172
rect 18690 11160 18696 11172
rect 18748 11160 18754 11212
rect 18414 11132 18420 11144
rect 16347 11104 18000 11132
rect 18375 11104 18420 11132
rect 16347 11101 16359 11104
rect 16301 11095 16359 11101
rect 18414 11092 18420 11104
rect 18472 11092 18478 11144
rect 18800 11132 18828 11240
rect 19794 11200 19800 11212
rect 19755 11172 19800 11200
rect 19794 11160 19800 11172
rect 19852 11160 19858 11212
rect 20346 11160 20352 11212
rect 20404 11200 20410 11212
rect 20809 11203 20867 11209
rect 20809 11200 20821 11203
rect 20404 11172 20821 11200
rect 20404 11160 20410 11172
rect 20809 11169 20821 11172
rect 20855 11169 20867 11203
rect 20809 11163 20867 11169
rect 20625 11135 20683 11141
rect 20625 11132 20637 11135
rect 18800 11104 20637 11132
rect 20625 11101 20637 11104
rect 20671 11101 20683 11135
rect 20625 11095 20683 11101
rect 12894 11024 12900 11076
rect 12952 11064 12958 11076
rect 15654 11064 15660 11076
rect 12952 11036 12997 11064
rect 15615 11036 15660 11064
rect 12952 11024 12958 11036
rect 15654 11024 15660 11036
rect 15712 11064 15718 11076
rect 16577 11067 16635 11073
rect 16577 11064 16589 11067
rect 15712 11036 16589 11064
rect 15712 11024 15718 11036
rect 16577 11033 16589 11036
rect 16623 11033 16635 11067
rect 16577 11027 16635 11033
rect 17034 11024 17040 11076
rect 17092 11064 17098 11076
rect 17681 11067 17739 11073
rect 17681 11064 17693 11067
rect 17092 11036 17693 11064
rect 17092 11024 17098 11036
rect 17681 11033 17693 11036
rect 17727 11033 17739 11067
rect 17681 11027 17739 11033
rect 17773 11067 17831 11073
rect 17773 11033 17785 11067
rect 17819 11064 17831 11067
rect 17819 11036 17908 11064
rect 17819 11033 17831 11036
rect 17773 11027 17831 11033
rect 12805 10999 12863 11005
rect 12805 10996 12817 10999
rect 12492 10968 12537 10996
rect 12728 10968 12817 10996
rect 12492 10956 12498 10968
rect 12805 10965 12817 10968
rect 12851 10965 12863 10999
rect 12805 10959 12863 10965
rect 13078 10956 13084 11008
rect 13136 10996 13142 11008
rect 13449 10999 13507 11005
rect 13449 10996 13461 10999
rect 13136 10968 13461 10996
rect 13136 10956 13142 10968
rect 13449 10965 13461 10968
rect 13495 10965 13507 10999
rect 13449 10959 13507 10965
rect 14182 10956 14188 11008
rect 14240 10996 14246 11008
rect 14553 10999 14611 11005
rect 14553 10996 14565 10999
rect 14240 10968 14565 10996
rect 14240 10956 14246 10968
rect 14553 10965 14565 10968
rect 14599 10965 14611 10999
rect 14553 10959 14611 10965
rect 14642 10956 14648 11008
rect 14700 10996 14706 11008
rect 15010 10996 15016 11008
rect 14700 10968 15016 10996
rect 14700 10956 14706 10968
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 17310 10996 17316 11008
rect 17271 10968 17316 10996
rect 17310 10956 17316 10968
rect 17368 10956 17374 11008
rect 17880 10996 17908 11036
rect 17954 11024 17960 11076
rect 18012 11064 18018 11076
rect 18693 11067 18751 11073
rect 18693 11064 18705 11067
rect 18012 11036 18705 11064
rect 18012 11024 18018 11036
rect 18693 11033 18705 11036
rect 18739 11033 18751 11067
rect 19702 11064 19708 11076
rect 19663 11036 19708 11064
rect 18693 11027 18751 11033
rect 19702 11024 19708 11036
rect 19760 11024 19766 11076
rect 20162 11024 20168 11076
rect 20220 11064 20226 11076
rect 20530 11064 20536 11076
rect 20220 11036 20536 11064
rect 20220 11024 20226 11036
rect 20530 11024 20536 11036
rect 20588 11064 20594 11076
rect 20717 11067 20775 11073
rect 20717 11064 20729 11067
rect 20588 11036 20729 11064
rect 20588 11024 20594 11036
rect 20717 11033 20729 11036
rect 20763 11033 20775 11067
rect 21266 11064 21272 11076
rect 21227 11036 21272 11064
rect 20717 11027 20775 11033
rect 21266 11024 21272 11036
rect 21324 11024 21330 11076
rect 22002 11024 22008 11076
rect 22060 11064 22066 11076
rect 22370 11064 22376 11076
rect 22060 11036 22376 11064
rect 22060 11024 22066 11036
rect 22370 11024 22376 11036
rect 22428 11024 22434 11076
rect 18874 10996 18880 11008
rect 17880 10968 18880 10996
rect 18874 10956 18880 10968
rect 18932 10956 18938 11008
rect 19334 10956 19340 11008
rect 19392 10996 19398 11008
rect 19613 10999 19671 11005
rect 19613 10996 19625 10999
rect 19392 10968 19625 10996
rect 19392 10956 19398 10968
rect 19613 10965 19625 10968
rect 19659 10965 19671 10999
rect 19613 10959 19671 10965
rect 19794 10956 19800 11008
rect 19852 10996 19858 11008
rect 20257 10999 20315 11005
rect 20257 10996 20269 10999
rect 19852 10968 20269 10996
rect 19852 10956 19858 10968
rect 20257 10965 20269 10968
rect 20303 10965 20315 10999
rect 20257 10959 20315 10965
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 5718 10752 5724 10804
rect 5776 10792 5782 10804
rect 5902 10792 5908 10804
rect 5776 10764 5908 10792
rect 5776 10752 5782 10764
rect 5902 10752 5908 10764
rect 5960 10752 5966 10804
rect 6730 10752 6736 10804
rect 6788 10792 6794 10804
rect 6788 10764 7144 10792
rect 6788 10752 6794 10764
rect 7116 10724 7144 10764
rect 7190 10752 7196 10804
rect 7248 10792 7254 10804
rect 7377 10795 7435 10801
rect 7377 10792 7389 10795
rect 7248 10764 7389 10792
rect 7248 10752 7254 10764
rect 7377 10761 7389 10764
rect 7423 10761 7435 10795
rect 7926 10792 7932 10804
rect 7887 10764 7932 10792
rect 7377 10755 7435 10761
rect 7926 10752 7932 10764
rect 7984 10752 7990 10804
rect 8297 10795 8355 10801
rect 8297 10761 8309 10795
rect 8343 10792 8355 10795
rect 8570 10792 8576 10804
rect 8343 10764 8576 10792
rect 8343 10761 8355 10764
rect 8297 10755 8355 10761
rect 8570 10752 8576 10764
rect 8628 10752 8634 10804
rect 10134 10792 10140 10804
rect 10095 10764 10140 10792
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 10410 10752 10416 10804
rect 10468 10792 10474 10804
rect 10686 10792 10692 10804
rect 10468 10764 10692 10792
rect 10468 10752 10474 10764
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 11149 10795 11207 10801
rect 11149 10761 11161 10795
rect 11195 10792 11207 10795
rect 12158 10792 12164 10804
rect 11195 10764 12164 10792
rect 11195 10761 11207 10764
rect 11149 10755 11207 10761
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 12805 10795 12863 10801
rect 12805 10792 12817 10795
rect 12492 10764 12817 10792
rect 12492 10752 12498 10764
rect 12805 10761 12817 10764
rect 12851 10761 12863 10795
rect 12805 10755 12863 10761
rect 13630 10752 13636 10804
rect 13688 10792 13694 10804
rect 13906 10792 13912 10804
rect 13688 10764 13912 10792
rect 13688 10752 13694 10764
rect 13906 10752 13912 10764
rect 13964 10752 13970 10804
rect 14366 10792 14372 10804
rect 14327 10764 14372 10792
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 17310 10792 17316 10804
rect 14660 10764 17316 10792
rect 7116 10696 7972 10724
rect 7944 10668 7972 10696
rect 8386 10684 8392 10736
rect 8444 10724 8450 10736
rect 8757 10727 8815 10733
rect 8757 10724 8769 10727
rect 8444 10696 8769 10724
rect 8444 10684 8450 10696
rect 8757 10693 8769 10696
rect 8803 10693 8815 10727
rect 8757 10687 8815 10693
rect 9769 10727 9827 10733
rect 9769 10693 9781 10727
rect 9815 10724 9827 10727
rect 11606 10724 11612 10736
rect 9815 10696 11612 10724
rect 9815 10693 9827 10696
rect 9769 10687 9827 10693
rect 11606 10684 11612 10696
rect 11664 10684 11670 10736
rect 12713 10727 12771 10733
rect 12713 10693 12725 10727
rect 12759 10724 12771 10727
rect 14660 10724 14688 10764
rect 17310 10752 17316 10764
rect 17368 10752 17374 10804
rect 17497 10795 17555 10801
rect 17497 10761 17509 10795
rect 17543 10792 17555 10795
rect 17678 10792 17684 10804
rect 17543 10764 17684 10792
rect 17543 10761 17555 10764
rect 17497 10755 17555 10761
rect 17678 10752 17684 10764
rect 17736 10752 17742 10804
rect 18138 10752 18144 10804
rect 18196 10792 18202 10804
rect 18233 10795 18291 10801
rect 18233 10792 18245 10795
rect 18196 10764 18245 10792
rect 18196 10752 18202 10764
rect 18233 10761 18245 10764
rect 18279 10792 18291 10795
rect 18414 10792 18420 10804
rect 18279 10764 18420 10792
rect 18279 10761 18291 10764
rect 18233 10755 18291 10761
rect 18414 10752 18420 10764
rect 18472 10752 18478 10804
rect 18693 10795 18751 10801
rect 18693 10761 18705 10795
rect 18739 10792 18751 10795
rect 19334 10792 19340 10804
rect 18739 10764 19340 10792
rect 18739 10761 18751 10764
rect 18693 10755 18751 10761
rect 19334 10752 19340 10764
rect 19392 10752 19398 10804
rect 19521 10795 19579 10801
rect 19521 10761 19533 10795
rect 19567 10792 19579 10795
rect 20257 10795 20315 10801
rect 20257 10792 20269 10795
rect 19567 10764 20269 10792
rect 19567 10761 19579 10764
rect 19521 10755 19579 10761
rect 20257 10761 20269 10764
rect 20303 10761 20315 10795
rect 20257 10755 20315 10761
rect 20622 10752 20628 10804
rect 20680 10792 20686 10804
rect 21269 10795 21327 10801
rect 21269 10792 21281 10795
rect 20680 10764 21281 10792
rect 20680 10752 20686 10764
rect 21269 10761 21281 10764
rect 21315 10761 21327 10795
rect 21269 10755 21327 10761
rect 12759 10696 14688 10724
rect 14829 10727 14887 10733
rect 12759 10693 12771 10696
rect 12713 10687 12771 10693
rect 14829 10693 14841 10727
rect 14875 10724 14887 10727
rect 16117 10727 16175 10733
rect 14875 10696 16068 10724
rect 14875 10693 14887 10696
rect 14829 10687 14887 10693
rect 6730 10656 6736 10668
rect 6691 10628 6736 10656
rect 6730 10616 6736 10628
rect 6788 10616 6794 10668
rect 7926 10616 7932 10668
rect 7984 10616 7990 10668
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10656 8723 10659
rect 8846 10656 8852 10668
rect 8711 10628 8852 10656
rect 8711 10625 8723 10628
rect 8665 10619 8723 10625
rect 8846 10616 8852 10628
rect 8904 10616 8910 10668
rect 9858 10656 9864 10668
rect 9600 10628 9864 10656
rect 6457 10591 6515 10597
rect 6457 10557 6469 10591
rect 6503 10557 6515 10591
rect 6457 10551 6515 10557
rect 6472 10520 6500 10551
rect 6546 10548 6552 10600
rect 6604 10588 6610 10600
rect 6641 10591 6699 10597
rect 6641 10588 6653 10591
rect 6604 10560 6653 10588
rect 6604 10548 6610 10560
rect 6641 10557 6653 10560
rect 6687 10557 6699 10591
rect 6641 10551 6699 10557
rect 6914 10548 6920 10600
rect 6972 10588 6978 10600
rect 8941 10591 8999 10597
rect 6972 10560 8708 10588
rect 6972 10548 6978 10560
rect 7466 10520 7472 10532
rect 6472 10492 7472 10520
rect 7466 10480 7472 10492
rect 7524 10480 7530 10532
rect 5718 10412 5724 10464
rect 5776 10452 5782 10464
rect 5905 10455 5963 10461
rect 5905 10452 5917 10455
rect 5776 10424 5917 10452
rect 5776 10412 5782 10424
rect 5905 10421 5917 10424
rect 5951 10421 5963 10455
rect 7098 10452 7104 10464
rect 7059 10424 7104 10452
rect 5905 10415 5963 10421
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 8680 10452 8708 10560
rect 8941 10557 8953 10591
rect 8987 10588 8999 10591
rect 9122 10588 9128 10600
rect 8987 10560 9128 10588
rect 8987 10557 8999 10560
rect 8941 10551 8999 10557
rect 9122 10548 9128 10560
rect 9180 10548 9186 10600
rect 9600 10597 9628 10628
rect 9858 10616 9864 10628
rect 9916 10616 9922 10668
rect 10781 10659 10839 10665
rect 10781 10625 10793 10659
rect 10827 10656 10839 10659
rect 11146 10656 11152 10668
rect 10827 10628 11152 10656
rect 10827 10625 10839 10628
rect 10781 10619 10839 10625
rect 11146 10616 11152 10628
rect 11204 10616 11210 10668
rect 11238 10616 11244 10668
rect 11296 10656 11302 10668
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 11296 10628 11529 10656
rect 11296 10616 11302 10628
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 13722 10656 13728 10668
rect 13683 10628 13728 10656
rect 11517 10619 11575 10625
rect 13722 10616 13728 10628
rect 13780 10616 13786 10668
rect 13814 10616 13820 10668
rect 13872 10616 13878 10668
rect 14737 10659 14795 10665
rect 14737 10625 14749 10659
rect 14783 10656 14795 10659
rect 14783 10628 15056 10656
rect 14783 10625 14795 10628
rect 14737 10619 14795 10625
rect 9585 10591 9643 10597
rect 9585 10557 9597 10591
rect 9631 10557 9643 10591
rect 9585 10551 9643 10557
rect 9677 10591 9735 10597
rect 9677 10557 9689 10591
rect 9723 10588 9735 10591
rect 10318 10588 10324 10600
rect 9723 10560 10324 10588
rect 9723 10557 9735 10560
rect 9677 10551 9735 10557
rect 10318 10548 10324 10560
rect 10376 10548 10382 10600
rect 10594 10588 10600 10600
rect 10555 10560 10600 10588
rect 10594 10548 10600 10560
rect 10652 10548 10658 10600
rect 10689 10591 10747 10597
rect 10689 10557 10701 10591
rect 10735 10588 10747 10591
rect 11054 10588 11060 10600
rect 10735 10560 11060 10588
rect 10735 10557 10747 10560
rect 10689 10551 10747 10557
rect 11054 10548 11060 10560
rect 11112 10548 11118 10600
rect 12069 10591 12127 10597
rect 12069 10557 12081 10591
rect 12115 10588 12127 10591
rect 12250 10588 12256 10600
rect 12115 10560 12256 10588
rect 12115 10557 12127 10560
rect 12069 10551 12127 10557
rect 12250 10548 12256 10560
rect 12308 10548 12314 10600
rect 12897 10591 12955 10597
rect 12897 10557 12909 10591
rect 12943 10557 12955 10591
rect 12897 10551 12955 10557
rect 13449 10591 13507 10597
rect 13449 10557 13461 10591
rect 13495 10557 13507 10591
rect 13630 10588 13636 10600
rect 13591 10560 13636 10588
rect 13449 10551 13507 10557
rect 10962 10480 10968 10532
rect 11020 10520 11026 10532
rect 12912 10520 12940 10551
rect 11020 10492 12940 10520
rect 13464 10520 13492 10551
rect 13630 10548 13636 10560
rect 13688 10548 13694 10600
rect 13832 10520 13860 10616
rect 14918 10588 14924 10600
rect 14879 10560 14924 10588
rect 14918 10548 14924 10560
rect 14976 10548 14982 10600
rect 15028 10588 15056 10628
rect 15194 10616 15200 10668
rect 15252 10656 15258 10668
rect 15841 10659 15899 10665
rect 15841 10656 15853 10659
rect 15252 10628 15853 10656
rect 15252 10616 15258 10628
rect 15841 10625 15853 10628
rect 15887 10625 15899 10659
rect 16040 10656 16068 10696
rect 16117 10693 16129 10727
rect 16163 10724 16175 10727
rect 16298 10724 16304 10736
rect 16163 10696 16304 10724
rect 16163 10693 16175 10696
rect 16117 10687 16175 10693
rect 16298 10684 16304 10696
rect 16356 10684 16362 10736
rect 19613 10727 19671 10733
rect 19613 10693 19625 10727
rect 19659 10724 19671 10727
rect 19794 10724 19800 10736
rect 19659 10696 19800 10724
rect 19659 10693 19671 10696
rect 19613 10687 19671 10693
rect 19794 10684 19800 10696
rect 19852 10684 19858 10736
rect 16666 10656 16672 10668
rect 16040 10628 16574 10656
rect 16627 10628 16672 10656
rect 15841 10619 15899 10625
rect 16546 10600 16574 10628
rect 16666 10616 16672 10628
rect 16724 10616 16730 10668
rect 16945 10659 17003 10665
rect 16945 10625 16957 10659
rect 16991 10656 17003 10659
rect 17494 10656 17500 10668
rect 16991 10628 17500 10656
rect 16991 10625 17003 10628
rect 16945 10619 17003 10625
rect 17494 10616 17500 10628
rect 17552 10616 17558 10668
rect 17681 10659 17739 10665
rect 17681 10625 17693 10659
rect 17727 10656 17739 10659
rect 17954 10656 17960 10668
rect 17727 10628 17960 10656
rect 17727 10625 17739 10628
rect 17681 10619 17739 10625
rect 17954 10616 17960 10628
rect 18012 10616 18018 10668
rect 18325 10659 18383 10665
rect 18325 10625 18337 10659
rect 18371 10656 18383 10659
rect 18690 10656 18696 10668
rect 18371 10628 18696 10656
rect 18371 10625 18383 10628
rect 18325 10619 18383 10625
rect 18690 10616 18696 10628
rect 18748 10616 18754 10668
rect 20070 10616 20076 10668
rect 20128 10656 20134 10668
rect 20622 10656 20628 10668
rect 20128 10628 20628 10656
rect 20128 10616 20134 10628
rect 20622 10616 20628 10628
rect 20680 10616 20686 10668
rect 22002 10616 22008 10668
rect 22060 10656 22066 10668
rect 22278 10656 22284 10668
rect 22060 10628 22284 10656
rect 22060 10616 22066 10628
rect 22278 10616 22284 10628
rect 22336 10616 22342 10668
rect 16206 10588 16212 10600
rect 15028 10560 16212 10588
rect 16206 10548 16212 10560
rect 16264 10548 16270 10600
rect 16546 10560 16580 10600
rect 16574 10548 16580 10560
rect 16632 10548 16638 10600
rect 18138 10588 18144 10600
rect 18099 10560 18144 10588
rect 18138 10548 18144 10560
rect 18196 10548 18202 10600
rect 18966 10548 18972 10600
rect 19024 10588 19030 10600
rect 19337 10591 19395 10597
rect 19337 10588 19349 10591
rect 19024 10560 19349 10588
rect 19024 10548 19030 10560
rect 19337 10557 19349 10560
rect 19383 10557 19395 10591
rect 20438 10588 20444 10600
rect 19337 10551 19395 10557
rect 19628 10560 20444 10588
rect 13464 10492 13860 10520
rect 14093 10523 14151 10529
rect 11020 10480 11026 10492
rect 14093 10489 14105 10523
rect 14139 10520 14151 10523
rect 19518 10520 19524 10532
rect 14139 10492 19524 10520
rect 14139 10489 14151 10492
rect 14093 10483 14151 10489
rect 19518 10480 19524 10492
rect 19576 10480 19582 10532
rect 12345 10455 12403 10461
rect 12345 10452 12357 10455
rect 8680 10424 12357 10452
rect 12345 10421 12357 10424
rect 12391 10421 12403 10455
rect 12345 10415 12403 10421
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12802 10452 12808 10464
rect 12492 10424 12808 10452
rect 12492 10412 12498 10424
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 13814 10412 13820 10464
rect 13872 10452 13878 10464
rect 13906 10452 13912 10464
rect 13872 10424 13912 10452
rect 13872 10412 13878 10424
rect 13906 10412 13912 10424
rect 13964 10412 13970 10464
rect 14182 10412 14188 10464
rect 14240 10452 14246 10464
rect 15473 10455 15531 10461
rect 15473 10452 15485 10455
rect 14240 10424 15485 10452
rect 14240 10412 14246 10424
rect 15473 10421 15485 10424
rect 15519 10452 15531 10455
rect 15746 10452 15752 10464
rect 15519 10424 15752 10452
rect 15519 10421 15531 10424
rect 15473 10415 15531 10421
rect 15746 10412 15752 10424
rect 15804 10412 15810 10464
rect 17494 10412 17500 10464
rect 17552 10452 17558 10464
rect 18046 10452 18052 10464
rect 17552 10424 18052 10452
rect 17552 10412 17558 10424
rect 18046 10412 18052 10424
rect 18104 10412 18110 10464
rect 18966 10412 18972 10464
rect 19024 10452 19030 10464
rect 19628 10452 19656 10560
rect 20438 10548 20444 10560
rect 20496 10588 20502 10600
rect 20717 10591 20775 10597
rect 20717 10588 20729 10591
rect 20496 10560 20729 10588
rect 20496 10548 20502 10560
rect 20717 10557 20729 10560
rect 20763 10557 20775 10591
rect 20717 10551 20775 10557
rect 20809 10591 20867 10597
rect 20809 10557 20821 10591
rect 20855 10557 20867 10591
rect 20809 10551 20867 10557
rect 20346 10480 20352 10532
rect 20404 10520 20410 10532
rect 20824 10520 20852 10551
rect 20404 10492 20852 10520
rect 20404 10480 20410 10492
rect 19024 10424 19656 10452
rect 19981 10455 20039 10461
rect 19024 10412 19030 10424
rect 19981 10421 19993 10455
rect 20027 10452 20039 10455
rect 20162 10452 20168 10464
rect 20027 10424 20168 10452
rect 20027 10421 20039 10424
rect 19981 10415 20039 10421
rect 20162 10412 20168 10424
rect 20220 10412 20226 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 7282 10208 7288 10260
rect 7340 10248 7346 10260
rect 7377 10251 7435 10257
rect 7377 10248 7389 10251
rect 7340 10220 7389 10248
rect 7340 10208 7346 10220
rect 7377 10217 7389 10220
rect 7423 10248 7435 10251
rect 8202 10248 8208 10260
rect 7423 10220 8208 10248
rect 7423 10217 7435 10220
rect 7377 10211 7435 10217
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 13081 10251 13139 10257
rect 13081 10248 13093 10251
rect 12860 10220 13093 10248
rect 12860 10208 12866 10220
rect 13081 10217 13093 10220
rect 13127 10217 13139 10251
rect 14550 10248 14556 10260
rect 14511 10220 14556 10248
rect 13081 10211 13139 10217
rect 14550 10208 14556 10220
rect 14608 10208 14614 10260
rect 17402 10208 17408 10260
rect 17460 10248 17466 10260
rect 17681 10251 17739 10257
rect 17681 10248 17693 10251
rect 17460 10220 17693 10248
rect 17460 10208 17466 10220
rect 17681 10217 17693 10220
rect 17727 10217 17739 10251
rect 21174 10248 21180 10260
rect 21135 10220 21180 10248
rect 17681 10211 17739 10217
rect 21174 10208 21180 10220
rect 21232 10208 21238 10260
rect 5534 10140 5540 10192
rect 5592 10180 5598 10192
rect 6365 10183 6423 10189
rect 6365 10180 6377 10183
rect 5592 10152 6377 10180
rect 5592 10140 5598 10152
rect 6365 10149 6377 10152
rect 6411 10149 6423 10183
rect 6365 10143 6423 10149
rect 7098 10140 7104 10192
rect 7156 10180 7162 10192
rect 16666 10180 16672 10192
rect 7156 10152 16672 10180
rect 7156 10140 7162 10152
rect 16666 10140 16672 10152
rect 16724 10140 16730 10192
rect 5258 10072 5264 10124
rect 5316 10112 5322 10124
rect 5442 10112 5448 10124
rect 5316 10084 5448 10112
rect 5316 10072 5322 10084
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 5629 10115 5687 10121
rect 5629 10081 5641 10115
rect 5675 10112 5687 10115
rect 5902 10112 5908 10124
rect 5675 10084 5908 10112
rect 5675 10081 5687 10084
rect 5629 10075 5687 10081
rect 5902 10072 5908 10084
rect 5960 10072 5966 10124
rect 6822 10112 6828 10124
rect 6656 10084 6828 10112
rect 4982 10004 4988 10056
rect 5040 10044 5046 10056
rect 6656 10044 6684 10084
rect 6822 10072 6828 10084
rect 6880 10112 6886 10124
rect 6917 10115 6975 10121
rect 6917 10112 6929 10115
rect 6880 10084 6929 10112
rect 6880 10072 6886 10084
rect 6917 10081 6929 10084
rect 6963 10081 6975 10115
rect 9214 10112 9220 10124
rect 9175 10084 9220 10112
rect 6917 10075 6975 10081
rect 9214 10072 9220 10084
rect 9272 10072 9278 10124
rect 9306 10072 9312 10124
rect 9364 10112 9370 10124
rect 10229 10115 10287 10121
rect 10229 10112 10241 10115
rect 9364 10084 10241 10112
rect 9364 10072 9370 10084
rect 10229 10081 10241 10084
rect 10275 10081 10287 10115
rect 11146 10112 11152 10124
rect 11107 10084 11152 10112
rect 10229 10075 10287 10081
rect 11146 10072 11152 10084
rect 11204 10072 11210 10124
rect 11606 10112 11612 10124
rect 11567 10084 11612 10112
rect 11606 10072 11612 10084
rect 11664 10072 11670 10124
rect 12529 10115 12587 10121
rect 12529 10081 12541 10115
rect 12575 10112 12587 10115
rect 13538 10112 13544 10124
rect 12575 10084 13544 10112
rect 12575 10081 12587 10084
rect 12529 10075 12587 10081
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 13722 10072 13728 10124
rect 13780 10112 13786 10124
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 13780 10084 14105 10112
rect 13780 10072 13786 10084
rect 14093 10081 14105 10084
rect 14139 10081 14151 10115
rect 14093 10075 14151 10081
rect 15749 10115 15807 10121
rect 15749 10081 15761 10115
rect 15795 10112 15807 10115
rect 15930 10112 15936 10124
rect 15795 10084 15936 10112
rect 15795 10081 15807 10084
rect 15749 10075 15807 10081
rect 15930 10072 15936 10084
rect 15988 10072 15994 10124
rect 17954 10112 17960 10124
rect 16776 10084 17960 10112
rect 5040 10016 6684 10044
rect 6733 10047 6791 10053
rect 5040 10004 5046 10016
rect 6733 10013 6745 10047
rect 6779 10044 6791 10047
rect 7282 10044 7288 10056
rect 6779 10016 7288 10044
rect 6779 10013 6791 10016
rect 6733 10007 6791 10013
rect 7282 10004 7288 10016
rect 7340 10004 7346 10056
rect 7926 10004 7932 10056
rect 7984 10044 7990 10056
rect 9401 10047 9459 10053
rect 9401 10044 9413 10047
rect 7984 10016 9413 10044
rect 7984 10004 7990 10016
rect 9401 10013 9413 10016
rect 9447 10044 9459 10047
rect 10502 10044 10508 10056
rect 9447 10016 10508 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 10502 10004 10508 10016
rect 10560 10004 10566 10056
rect 12250 10004 12256 10056
rect 12308 10044 12314 10056
rect 12713 10047 12771 10053
rect 12713 10044 12725 10047
rect 12308 10016 12725 10044
rect 12308 10004 12314 10016
rect 12713 10013 12725 10016
rect 12759 10013 12771 10047
rect 12713 10007 12771 10013
rect 15194 10004 15200 10056
rect 15252 10004 15258 10056
rect 15473 10047 15531 10053
rect 15473 10013 15485 10047
rect 15519 10044 15531 10047
rect 16776 10044 16804 10084
rect 17954 10072 17960 10084
rect 18012 10072 18018 10124
rect 18322 10112 18328 10124
rect 18283 10084 18328 10112
rect 18322 10072 18328 10084
rect 18380 10072 18386 10124
rect 18690 10112 18696 10124
rect 18651 10084 18696 10112
rect 18690 10072 18696 10084
rect 18748 10072 18754 10124
rect 19444 10084 21036 10112
rect 16942 10044 16948 10056
rect 15519 10016 16804 10044
rect 16903 10016 16948 10044
rect 15519 10013 15531 10016
rect 15473 10007 15531 10013
rect 5350 9936 5356 9988
rect 5408 9976 5414 9988
rect 7745 9979 7803 9985
rect 7745 9976 7757 9979
rect 5408 9948 7757 9976
rect 5408 9936 5414 9948
rect 7745 9945 7757 9948
rect 7791 9976 7803 9979
rect 8386 9976 8392 9988
rect 7791 9948 8392 9976
rect 7791 9945 7803 9948
rect 7745 9939 7803 9945
rect 8386 9936 8392 9948
rect 8444 9936 8450 9988
rect 9950 9936 9956 9988
rect 10008 9976 10014 9988
rect 15212 9976 15240 10004
rect 15948 9988 15976 10016
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 17221 10047 17279 10053
rect 17221 10013 17233 10047
rect 17267 10044 17279 10047
rect 19444 10044 19472 10084
rect 17267 10016 19472 10044
rect 17267 10013 17279 10016
rect 17221 10007 17279 10013
rect 19518 10004 19524 10056
rect 19576 10044 19582 10056
rect 20254 10044 20260 10056
rect 19576 10016 19621 10044
rect 20215 10016 20260 10044
rect 19576 10004 19582 10016
rect 20254 10004 20260 10016
rect 20312 10004 20318 10056
rect 21008 10053 21036 10084
rect 20993 10047 21051 10053
rect 20993 10013 21005 10047
rect 21039 10013 21051 10047
rect 20993 10007 21051 10013
rect 10008 9948 15240 9976
rect 10008 9936 10014 9948
rect 15930 9936 15936 9988
rect 15988 9936 15994 9988
rect 16209 9979 16267 9985
rect 16209 9945 16221 9979
rect 16255 9976 16267 9979
rect 16574 9976 16580 9988
rect 16255 9948 16580 9976
rect 16255 9945 16267 9948
rect 16209 9939 16267 9945
rect 16574 9936 16580 9948
rect 16632 9976 16638 9988
rect 17402 9976 17408 9988
rect 16632 9948 17408 9976
rect 16632 9936 16638 9948
rect 17402 9936 17408 9948
rect 17460 9936 17466 9988
rect 19797 9979 19855 9985
rect 19797 9945 19809 9979
rect 19843 9945 19855 9979
rect 19797 9939 19855 9945
rect 5718 9908 5724 9920
rect 5679 9880 5724 9908
rect 5718 9868 5724 9880
rect 5776 9868 5782 9920
rect 5994 9868 6000 9920
rect 6052 9908 6058 9920
rect 6089 9911 6147 9917
rect 6089 9908 6101 9911
rect 6052 9880 6101 9908
rect 6052 9868 6058 9880
rect 6089 9877 6101 9880
rect 6135 9877 6147 9911
rect 6089 9871 6147 9877
rect 6825 9911 6883 9917
rect 6825 9877 6837 9911
rect 6871 9908 6883 9911
rect 7006 9908 7012 9920
rect 6871 9880 7012 9908
rect 6871 9877 6883 9880
rect 6825 9871 6883 9877
rect 7006 9868 7012 9880
rect 7064 9908 7070 9920
rect 7466 9908 7472 9920
rect 7064 9880 7472 9908
rect 7064 9868 7070 9880
rect 7466 9868 7472 9880
rect 7524 9868 7530 9920
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 8113 9911 8171 9917
rect 8113 9908 8125 9911
rect 7984 9880 8125 9908
rect 7984 9868 7990 9880
rect 8113 9877 8125 9880
rect 8159 9877 8171 9911
rect 8570 9908 8576 9920
rect 8531 9880 8576 9908
rect 8113 9871 8171 9877
rect 8570 9868 8576 9880
rect 8628 9868 8634 9920
rect 9493 9911 9551 9917
rect 9493 9877 9505 9911
rect 9539 9908 9551 9911
rect 9674 9908 9680 9920
rect 9539 9880 9680 9908
rect 9539 9877 9551 9880
rect 9493 9871 9551 9877
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 9858 9908 9864 9920
rect 9819 9880 9864 9908
rect 9858 9868 9864 9880
rect 9916 9868 9922 9920
rect 10410 9908 10416 9920
rect 10371 9880 10416 9908
rect 10410 9868 10416 9880
rect 10468 9868 10474 9920
rect 10502 9868 10508 9920
rect 10560 9908 10566 9920
rect 10873 9911 10931 9917
rect 10560 9880 10605 9908
rect 10560 9868 10566 9880
rect 10873 9877 10885 9911
rect 10919 9908 10931 9911
rect 11238 9908 11244 9920
rect 10919 9880 11244 9908
rect 10919 9877 10931 9880
rect 10873 9871 10931 9877
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 12618 9908 12624 9920
rect 12579 9880 12624 9908
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 13354 9868 13360 9920
rect 13412 9908 13418 9920
rect 13449 9911 13507 9917
rect 13449 9908 13461 9911
rect 13412 9880 13461 9908
rect 13412 9868 13418 9880
rect 13449 9877 13461 9880
rect 13495 9908 13507 9911
rect 13722 9908 13728 9920
rect 13495 9880 13728 9908
rect 13495 9877 13507 9880
rect 13449 9871 13507 9877
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 15102 9908 15108 9920
rect 15063 9880 15108 9908
rect 15102 9868 15108 9880
rect 15160 9868 15166 9920
rect 15194 9868 15200 9920
rect 15252 9908 15258 9920
rect 15565 9911 15623 9917
rect 15565 9908 15577 9911
rect 15252 9880 15577 9908
rect 15252 9868 15258 9880
rect 15565 9877 15577 9880
rect 15611 9877 15623 9911
rect 15565 9871 15623 9877
rect 16669 9911 16727 9917
rect 16669 9877 16681 9911
rect 16715 9908 16727 9911
rect 17034 9908 17040 9920
rect 16715 9880 17040 9908
rect 16715 9877 16727 9880
rect 16669 9871 16727 9877
rect 17034 9868 17040 9880
rect 17092 9868 17098 9920
rect 18046 9908 18052 9920
rect 18007 9880 18052 9908
rect 18046 9868 18052 9880
rect 18104 9868 18110 9920
rect 18138 9868 18144 9920
rect 18196 9908 18202 9920
rect 19812 9908 19840 9939
rect 19886 9936 19892 9988
rect 19944 9976 19950 9988
rect 20533 9979 20591 9985
rect 20533 9976 20545 9979
rect 19944 9948 20545 9976
rect 19944 9936 19950 9948
rect 20533 9945 20545 9948
rect 20579 9945 20591 9979
rect 20533 9939 20591 9945
rect 20806 9908 20812 9920
rect 18196 9880 18241 9908
rect 19812 9880 20812 9908
rect 18196 9868 18202 9880
rect 20806 9868 20812 9880
rect 20864 9868 20870 9920
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 5994 9664 6000 9716
rect 6052 9704 6058 9716
rect 6733 9707 6791 9713
rect 6733 9704 6745 9707
rect 6052 9676 6745 9704
rect 6052 9664 6058 9676
rect 6733 9673 6745 9676
rect 6779 9673 6791 9707
rect 6733 9667 6791 9673
rect 9858 9664 9864 9716
rect 9916 9704 9922 9716
rect 10229 9707 10287 9713
rect 10229 9704 10241 9707
rect 9916 9676 10241 9704
rect 9916 9664 9922 9676
rect 10229 9673 10241 9676
rect 10275 9673 10287 9707
rect 10229 9667 10287 9673
rect 10502 9664 10508 9716
rect 10560 9704 10566 9716
rect 10873 9707 10931 9713
rect 10873 9704 10885 9707
rect 10560 9676 10885 9704
rect 10560 9664 10566 9676
rect 10873 9673 10885 9676
rect 10919 9673 10931 9707
rect 10873 9667 10931 9673
rect 11238 9664 11244 9716
rect 11296 9704 11302 9716
rect 14737 9707 14795 9713
rect 11296 9676 12434 9704
rect 11296 9664 11302 9676
rect 6638 9636 6644 9648
rect 6599 9608 6644 9636
rect 6638 9596 6644 9608
rect 6696 9596 6702 9648
rect 8662 9636 8668 9648
rect 7576 9608 8064 9636
rect 8623 9608 8668 9636
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 5629 9571 5687 9577
rect 5629 9568 5641 9571
rect 5031 9540 5641 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5629 9537 5641 9540
rect 5675 9568 5687 9571
rect 5718 9568 5724 9580
rect 5675 9540 5724 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 5718 9528 5724 9540
rect 5776 9568 5782 9580
rect 7576 9568 7604 9608
rect 7742 9568 7748 9580
rect 5776 9540 7604 9568
rect 7703 9540 7748 9568
rect 5776 9528 5782 9540
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 8036 9568 8064 9608
rect 8662 9596 8668 9608
rect 8720 9596 8726 9648
rect 11609 9639 11667 9645
rect 11609 9605 11621 9639
rect 11655 9636 11667 9639
rect 11698 9636 11704 9648
rect 11655 9608 11704 9636
rect 11655 9605 11667 9608
rect 11609 9599 11667 9605
rect 11698 9596 11704 9608
rect 11756 9596 11762 9648
rect 12406 9636 12434 9676
rect 14737 9673 14749 9707
rect 14783 9704 14795 9707
rect 15102 9704 15108 9716
rect 14783 9676 15108 9704
rect 14783 9673 14795 9676
rect 14737 9667 14795 9673
rect 15102 9664 15108 9676
rect 15160 9664 15166 9716
rect 17034 9704 17040 9716
rect 16995 9676 17040 9704
rect 17034 9664 17040 9676
rect 17092 9664 17098 9716
rect 18138 9664 18144 9716
rect 18196 9704 18202 9716
rect 18417 9707 18475 9713
rect 18417 9704 18429 9707
rect 18196 9676 18429 9704
rect 18196 9664 18202 9676
rect 18417 9673 18429 9676
rect 18463 9673 18475 9707
rect 18417 9667 18475 9673
rect 20530 9664 20536 9716
rect 20588 9664 20594 9716
rect 12406 9608 18736 9636
rect 8754 9568 8760 9580
rect 8036 9540 8760 9568
rect 8754 9528 8760 9540
rect 8812 9528 8818 9580
rect 9306 9528 9312 9580
rect 9364 9568 9370 9580
rect 9401 9571 9459 9577
rect 9401 9568 9413 9571
rect 9364 9540 9413 9568
rect 9364 9528 9370 9540
rect 9401 9537 9413 9540
rect 9447 9537 9459 9571
rect 11974 9568 11980 9580
rect 9401 9531 9459 9537
rect 10060 9540 11980 9568
rect 4798 9460 4804 9512
rect 4856 9500 4862 9512
rect 5353 9503 5411 9509
rect 5353 9500 5365 9503
rect 4856 9472 5365 9500
rect 4856 9460 4862 9472
rect 5353 9469 5365 9472
rect 5399 9469 5411 9503
rect 5353 9463 5411 9469
rect 5537 9503 5595 9509
rect 5537 9469 5549 9503
rect 5583 9500 5595 9503
rect 5902 9500 5908 9512
rect 5583 9472 5908 9500
rect 5583 9469 5595 9472
rect 5537 9463 5595 9469
rect 5368 9432 5396 9463
rect 5718 9432 5724 9444
rect 5368 9404 5724 9432
rect 5718 9392 5724 9404
rect 5776 9392 5782 9444
rect 4617 9367 4675 9373
rect 4617 9333 4629 9367
rect 4663 9364 4675 9367
rect 5828 9364 5856 9472
rect 5902 9460 5908 9472
rect 5960 9500 5966 9512
rect 6270 9500 6276 9512
rect 5960 9472 6276 9500
rect 5960 9460 5966 9472
rect 6270 9460 6276 9472
rect 6328 9460 6334 9512
rect 6549 9503 6607 9509
rect 6549 9469 6561 9503
rect 6595 9500 6607 9503
rect 6638 9500 6644 9512
rect 6595 9472 6644 9500
rect 6595 9469 6607 9472
rect 6549 9463 6607 9469
rect 6638 9460 6644 9472
rect 6696 9460 6702 9512
rect 7558 9500 7564 9512
rect 7519 9472 7564 9500
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 7653 9503 7711 9509
rect 7653 9469 7665 9503
rect 7699 9469 7711 9503
rect 7653 9463 7711 9469
rect 8573 9503 8631 9509
rect 8573 9469 8585 9503
rect 8619 9500 8631 9503
rect 9214 9500 9220 9512
rect 8619 9472 9220 9500
rect 8619 9469 8631 9472
rect 8573 9463 8631 9469
rect 7101 9435 7159 9441
rect 7101 9401 7113 9435
rect 7147 9432 7159 9435
rect 7668 9432 7696 9463
rect 9214 9460 9220 9472
rect 9272 9460 9278 9512
rect 10060 9509 10088 9540
rect 11974 9528 11980 9540
rect 12032 9528 12038 9580
rect 12529 9571 12587 9577
rect 12529 9537 12541 9571
rect 12575 9537 12587 9571
rect 12529 9531 12587 9537
rect 12621 9571 12679 9577
rect 12621 9537 12633 9571
rect 12667 9568 12679 9571
rect 12667 9540 13216 9568
rect 12667 9537 12679 9540
rect 12621 9531 12679 9537
rect 10045 9503 10103 9509
rect 10045 9469 10057 9503
rect 10091 9469 10103 9503
rect 10045 9463 10103 9469
rect 10137 9503 10195 9509
rect 10137 9469 10149 9503
rect 10183 9469 10195 9503
rect 10137 9463 10195 9469
rect 8110 9432 8116 9444
rect 7147 9404 7696 9432
rect 8071 9404 8116 9432
rect 7147 9401 7159 9404
rect 7101 9395 7159 9401
rect 8110 9392 8116 9404
rect 8168 9392 8174 9444
rect 9125 9435 9183 9441
rect 9125 9401 9137 9435
rect 9171 9432 9183 9435
rect 10152 9432 10180 9463
rect 12158 9432 12164 9444
rect 9171 9404 10180 9432
rect 10428 9404 12020 9432
rect 12119 9404 12164 9432
rect 9171 9401 9183 9404
rect 9125 9395 9183 9401
rect 4663 9336 5856 9364
rect 5997 9367 6055 9373
rect 4663 9333 4675 9336
rect 4617 9327 4675 9333
rect 5997 9333 6009 9367
rect 6043 9364 6055 9367
rect 7190 9364 7196 9376
rect 6043 9336 7196 9364
rect 6043 9333 6055 9336
rect 5997 9327 6055 9333
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 10428 9364 10456 9404
rect 7340 9336 10456 9364
rect 10597 9367 10655 9373
rect 7340 9324 7346 9336
rect 10597 9333 10609 9367
rect 10643 9364 10655 9367
rect 11882 9364 11888 9376
rect 10643 9336 11888 9364
rect 10643 9333 10655 9336
rect 10597 9327 10655 9333
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 11992 9364 12020 9404
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 12544 9432 12572 9531
rect 12802 9500 12808 9512
rect 12763 9472 12808 9500
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 13188 9500 13216 9540
rect 13262 9528 13268 9580
rect 13320 9568 13326 9580
rect 13541 9571 13599 9577
rect 13541 9568 13553 9571
rect 13320 9540 13553 9568
rect 13320 9528 13326 9540
rect 13541 9537 13553 9540
rect 13587 9537 13599 9571
rect 13541 9531 13599 9537
rect 14645 9571 14703 9577
rect 14645 9537 14657 9571
rect 14691 9568 14703 9571
rect 14918 9568 14924 9580
rect 14691 9540 14924 9568
rect 14691 9537 14703 9540
rect 14645 9531 14703 9537
rect 14918 9528 14924 9540
rect 14976 9528 14982 9580
rect 15654 9568 15660 9580
rect 15615 9540 15660 9568
rect 15654 9528 15660 9540
rect 15712 9528 15718 9580
rect 17126 9568 17132 9580
rect 16868 9540 17132 9568
rect 13633 9503 13691 9509
rect 13188 9472 13492 9500
rect 13173 9435 13231 9441
rect 13173 9432 13185 9435
rect 12544 9404 13185 9432
rect 13173 9401 13185 9404
rect 13219 9401 13231 9435
rect 13464 9432 13492 9472
rect 13633 9469 13645 9503
rect 13679 9500 13691 9503
rect 13722 9500 13728 9512
rect 13679 9472 13728 9500
rect 13679 9469 13691 9472
rect 13633 9463 13691 9469
rect 13722 9460 13728 9472
rect 13780 9460 13786 9512
rect 13817 9503 13875 9509
rect 13817 9469 13829 9503
rect 13863 9500 13875 9503
rect 14550 9500 14556 9512
rect 13863 9472 14556 9500
rect 13863 9469 13875 9472
rect 13817 9463 13875 9469
rect 14550 9460 14556 9472
rect 14608 9500 14614 9512
rect 14829 9503 14887 9509
rect 14829 9500 14841 9503
rect 14608 9472 14841 9500
rect 14608 9460 14614 9472
rect 14829 9469 14841 9472
rect 14875 9469 14887 9503
rect 14829 9463 14887 9469
rect 15102 9460 15108 9512
rect 15160 9500 15166 9512
rect 15381 9503 15439 9509
rect 15381 9500 15393 9503
rect 15160 9472 15393 9500
rect 15160 9460 15166 9472
rect 15381 9469 15393 9472
rect 15427 9469 15439 9503
rect 15381 9463 15439 9469
rect 15565 9503 15623 9509
rect 15565 9469 15577 9503
rect 15611 9500 15623 9503
rect 15746 9500 15752 9512
rect 15611 9472 15752 9500
rect 15611 9469 15623 9472
rect 15565 9463 15623 9469
rect 15746 9460 15752 9472
rect 15804 9500 15810 9512
rect 16390 9500 16396 9512
rect 15804 9472 16396 9500
rect 15804 9460 15810 9472
rect 16390 9460 16396 9472
rect 16448 9460 16454 9512
rect 16574 9460 16580 9512
rect 16632 9500 16638 9512
rect 16868 9509 16896 9540
rect 17126 9528 17132 9540
rect 17184 9528 17190 9580
rect 17678 9528 17684 9580
rect 17736 9568 17742 9580
rect 18708 9577 18736 9608
rect 20254 9596 20260 9648
rect 20312 9636 20318 9648
rect 20548 9636 20576 9664
rect 20625 9639 20683 9645
rect 20625 9636 20637 9639
rect 20312 9608 20637 9636
rect 20312 9596 20318 9608
rect 20625 9605 20637 9608
rect 20671 9605 20683 9639
rect 20625 9599 20683 9605
rect 18049 9571 18107 9577
rect 18049 9568 18061 9571
rect 17736 9540 18061 9568
rect 17736 9528 17742 9540
rect 18049 9537 18061 9540
rect 18095 9537 18107 9571
rect 18049 9531 18107 9537
rect 18693 9571 18751 9577
rect 18693 9537 18705 9571
rect 18739 9537 18751 9571
rect 19886 9568 19892 9580
rect 19847 9540 19892 9568
rect 18693 9531 18751 9537
rect 19886 9528 19892 9540
rect 19944 9528 19950 9580
rect 20533 9571 20591 9577
rect 20533 9537 20545 9571
rect 20579 9568 20591 9571
rect 21177 9571 21235 9577
rect 21177 9568 21189 9571
rect 20579 9540 21189 9568
rect 20579 9537 20591 9540
rect 20533 9531 20591 9537
rect 21177 9537 21189 9540
rect 21223 9537 21235 9571
rect 21177 9531 21235 9537
rect 16853 9503 16911 9509
rect 16853 9500 16865 9503
rect 16632 9472 16865 9500
rect 16632 9460 16638 9472
rect 16853 9469 16865 9472
rect 16899 9469 16911 9503
rect 16853 9463 16911 9469
rect 16942 9460 16948 9512
rect 17000 9500 17006 9512
rect 17865 9503 17923 9509
rect 17000 9472 17045 9500
rect 17000 9460 17006 9472
rect 17865 9469 17877 9503
rect 17911 9469 17923 9503
rect 17865 9463 17923 9469
rect 17957 9503 18015 9509
rect 17957 9469 17969 9503
rect 18003 9500 18015 9503
rect 18138 9500 18144 9512
rect 18003 9472 18144 9500
rect 18003 9469 18015 9472
rect 17957 9463 18015 9469
rect 14277 9435 14335 9441
rect 14277 9432 14289 9435
rect 13464 9404 14289 9432
rect 13173 9395 13231 9401
rect 14277 9401 14289 9404
rect 14323 9401 14335 9435
rect 14277 9395 14335 9401
rect 16025 9435 16083 9441
rect 16025 9401 16037 9435
rect 16071 9432 16083 9435
rect 17126 9432 17132 9444
rect 16071 9404 17132 9432
rect 16071 9401 16083 9404
rect 16025 9395 16083 9401
rect 17126 9392 17132 9404
rect 17184 9392 17190 9444
rect 17880 9432 17908 9463
rect 18138 9460 18144 9472
rect 18196 9460 18202 9512
rect 18874 9500 18880 9512
rect 18835 9472 18880 9500
rect 18874 9460 18880 9472
rect 18932 9460 18938 9512
rect 19334 9460 19340 9512
rect 19392 9500 19398 9512
rect 20717 9503 20775 9509
rect 19392 9472 20392 9500
rect 19392 9460 19398 9472
rect 20364 9444 20392 9472
rect 20717 9469 20729 9503
rect 20763 9469 20775 9503
rect 20717 9463 20775 9469
rect 17880 9404 18000 9432
rect 14550 9364 14556 9376
rect 11992 9336 14556 9364
rect 14550 9324 14556 9336
rect 14608 9324 14614 9376
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 16942 9364 16948 9376
rect 16356 9336 16948 9364
rect 16356 9324 16362 9336
rect 16942 9324 16948 9336
rect 17000 9324 17006 9376
rect 17034 9324 17040 9376
rect 17092 9364 17098 9376
rect 17405 9367 17463 9373
rect 17405 9364 17417 9367
rect 17092 9336 17417 9364
rect 17092 9324 17098 9336
rect 17405 9333 17417 9336
rect 17451 9333 17463 9367
rect 17972 9364 18000 9404
rect 18046 9392 18052 9444
rect 18104 9432 18110 9444
rect 20165 9435 20223 9441
rect 20165 9432 20177 9435
rect 18104 9404 20177 9432
rect 18104 9392 18110 9404
rect 20165 9401 20177 9404
rect 20211 9401 20223 9435
rect 20165 9395 20223 9401
rect 20346 9392 20352 9444
rect 20404 9432 20410 9444
rect 20732 9432 20760 9463
rect 20404 9404 20760 9432
rect 20404 9392 20410 9404
rect 19334 9364 19340 9376
rect 17972 9336 19340 9364
rect 17405 9327 17463 9333
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 19705 9367 19763 9373
rect 19705 9333 19717 9367
rect 19751 9364 19763 9367
rect 19978 9364 19984 9376
rect 19751 9336 19984 9364
rect 19751 9333 19763 9336
rect 19705 9327 19763 9333
rect 19978 9324 19984 9336
rect 20036 9324 20042 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 5905 9163 5963 9169
rect 5905 9129 5917 9163
rect 5951 9160 5963 9163
rect 6546 9160 6552 9172
rect 5951 9132 6552 9160
rect 5951 9129 5963 9132
rect 5905 9123 5963 9129
rect 6546 9120 6552 9132
rect 6604 9120 6610 9172
rect 6638 9120 6644 9172
rect 6696 9160 6702 9172
rect 9582 9160 9588 9172
rect 6696 9132 9588 9160
rect 6696 9120 6702 9132
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 9950 9160 9956 9172
rect 9911 9132 9956 9160
rect 9950 9120 9956 9132
rect 10008 9120 10014 9172
rect 10410 9120 10416 9172
rect 10468 9160 10474 9172
rect 11885 9163 11943 9169
rect 11885 9160 11897 9163
rect 10468 9132 11897 9160
rect 10468 9120 10474 9132
rect 11885 9129 11897 9132
rect 11931 9129 11943 9163
rect 11885 9123 11943 9129
rect 11974 9120 11980 9172
rect 12032 9160 12038 9172
rect 13998 9160 14004 9172
rect 12032 9132 14004 9160
rect 12032 9120 12038 9132
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 14182 9160 14188 9172
rect 14095 9132 14188 9160
rect 14182 9120 14188 9132
rect 14240 9160 14246 9172
rect 14918 9160 14924 9172
rect 14240 9132 14924 9160
rect 14240 9120 14246 9132
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 15102 9160 15108 9172
rect 15063 9132 15108 9160
rect 15102 9120 15108 9132
rect 15160 9120 15166 9172
rect 15746 9120 15752 9172
rect 15804 9160 15810 9172
rect 16206 9160 16212 9172
rect 15804 9132 16212 9160
rect 15804 9120 15810 9132
rect 16206 9120 16212 9132
rect 16264 9120 16270 9172
rect 17678 9160 17684 9172
rect 17639 9132 17684 9160
rect 17678 9120 17684 9132
rect 17736 9120 17742 9172
rect 18782 9160 18788 9172
rect 18156 9132 18788 9160
rect 7834 9092 7840 9104
rect 6104 9064 7840 9092
rect 5353 9027 5411 9033
rect 5353 8993 5365 9027
rect 5399 9024 5411 9027
rect 5994 9024 6000 9036
rect 5399 8996 6000 9024
rect 5399 8993 5411 8996
rect 5353 8987 5411 8993
rect 5994 8984 6000 8996
rect 6052 9024 6058 9036
rect 6104 9024 6132 9064
rect 7834 9052 7840 9064
rect 7892 9052 7898 9104
rect 10870 9092 10876 9104
rect 9232 9064 10876 9092
rect 6052 8996 6132 9024
rect 7009 9027 7067 9033
rect 6052 8984 6058 8996
rect 7009 8993 7021 9027
rect 7055 9024 7067 9027
rect 9232 9024 9260 9064
rect 10870 9052 10876 9064
rect 10928 9052 10934 9104
rect 15654 9052 15660 9104
rect 15712 9092 15718 9104
rect 17954 9092 17960 9104
rect 15712 9064 17960 9092
rect 15712 9052 15718 9064
rect 17954 9052 17960 9064
rect 18012 9052 18018 9104
rect 9398 9024 9404 9036
rect 7055 8996 9260 9024
rect 9359 8996 9404 9024
rect 7055 8993 7067 8996
rect 7009 8987 7067 8993
rect 9398 8984 9404 8996
rect 9456 8984 9462 9036
rect 9674 8984 9680 9036
rect 9732 9024 9738 9036
rect 10229 9027 10287 9033
rect 10229 9024 10241 9027
rect 9732 8996 10241 9024
rect 9732 8984 9738 8996
rect 10229 8993 10241 8996
rect 10275 8993 10287 9027
rect 12526 9024 12532 9036
rect 12487 8996 12532 9024
rect 10229 8987 10287 8993
rect 12526 8984 12532 8996
rect 12584 8984 12590 9036
rect 13262 9024 13268 9036
rect 13223 8996 13268 9024
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 15933 9027 15991 9033
rect 15933 8993 15945 9027
rect 15979 9024 15991 9027
rect 16574 9024 16580 9036
rect 15979 8996 16580 9024
rect 15979 8993 15991 8996
rect 15933 8987 15991 8993
rect 16574 8984 16580 8996
rect 16632 8984 16638 9036
rect 18156 9033 18184 9132
rect 18782 9120 18788 9132
rect 18840 9160 18846 9172
rect 19426 9160 19432 9172
rect 18840 9132 19432 9160
rect 18840 9120 18846 9132
rect 19426 9120 19432 9132
rect 19484 9120 19490 9172
rect 19702 9120 19708 9172
rect 19760 9160 19766 9172
rect 20441 9163 20499 9169
rect 20441 9160 20453 9163
rect 19760 9132 20453 9160
rect 19760 9120 19766 9132
rect 20441 9129 20453 9132
rect 20487 9129 20499 9163
rect 20441 9123 20499 9129
rect 18230 9052 18236 9104
rect 18288 9092 18294 9104
rect 18288 9064 21036 9092
rect 18288 9052 18294 9064
rect 18141 9027 18199 9033
rect 18141 8993 18153 9027
rect 18187 8993 18199 9027
rect 18141 8987 18199 8993
rect 18325 9027 18383 9033
rect 18325 8993 18337 9027
rect 18371 9024 18383 9027
rect 18506 9024 18512 9036
rect 18371 8996 18512 9024
rect 18371 8993 18383 8996
rect 18325 8987 18383 8993
rect 18506 8984 18512 8996
rect 18564 8984 18570 9036
rect 18966 8984 18972 9036
rect 19024 9024 19030 9036
rect 21008 9033 21036 9064
rect 19981 9027 20039 9033
rect 19981 9024 19993 9027
rect 19024 8996 19993 9024
rect 19024 8984 19030 8996
rect 19981 8993 19993 8996
rect 20027 8993 20039 9027
rect 19981 8987 20039 8993
rect 20993 9027 21051 9033
rect 20993 8993 21005 9027
rect 21039 8993 21051 9027
rect 20993 8987 21051 8993
rect 5534 8956 5540 8968
rect 5495 8928 5540 8956
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 7190 8956 7196 8968
rect 7151 8928 7196 8956
rect 7190 8916 7196 8928
rect 7248 8916 7254 8968
rect 9585 8959 9643 8965
rect 9585 8925 9597 8959
rect 9631 8956 9643 8959
rect 10134 8956 10140 8968
rect 9631 8928 10140 8956
rect 9631 8925 9643 8928
rect 9585 8919 9643 8925
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 12253 8959 12311 8965
rect 12253 8956 12265 8959
rect 11204 8928 12265 8956
rect 11204 8916 11210 8928
rect 12253 8925 12265 8928
rect 12299 8925 12311 8959
rect 12253 8919 12311 8925
rect 13998 8916 14004 8968
rect 14056 8956 14062 8968
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 14056 8928 16865 8956
rect 14056 8916 14062 8928
rect 16853 8925 16865 8928
rect 16899 8925 16911 8959
rect 18046 8956 18052 8968
rect 18007 8928 18052 8956
rect 16853 8919 16911 8925
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 18230 8916 18236 8968
rect 18288 8956 18294 8968
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 18288 8928 19257 8956
rect 18288 8916 18294 8928
rect 19245 8925 19257 8928
rect 19291 8925 19303 8959
rect 20806 8956 20812 8968
rect 19245 8919 19303 8925
rect 19352 8928 20812 8956
rect 4706 8848 4712 8900
rect 4764 8888 4770 8900
rect 5445 8891 5503 8897
rect 5445 8888 5457 8891
rect 4764 8860 5457 8888
rect 4764 8848 4770 8860
rect 5445 8857 5457 8860
rect 5491 8857 5503 8891
rect 5445 8851 5503 8857
rect 5810 8848 5816 8900
rect 5868 8888 5874 8900
rect 7101 8891 7159 8897
rect 7101 8888 7113 8891
rect 5868 8860 7113 8888
rect 5868 8848 5874 8860
rect 7101 8857 7113 8860
rect 7147 8857 7159 8891
rect 9493 8891 9551 8897
rect 9493 8888 9505 8891
rect 7101 8851 7159 8857
rect 7576 8860 9505 8888
rect 6270 8820 6276 8832
rect 6183 8792 6276 8820
rect 6270 8780 6276 8792
rect 6328 8820 6334 8832
rect 7282 8820 7288 8832
rect 6328 8792 7288 8820
rect 6328 8780 6334 8792
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 7576 8829 7604 8860
rect 9493 8857 9505 8860
rect 9539 8857 9551 8891
rect 9493 8851 9551 8857
rect 9646 8860 12112 8888
rect 7561 8823 7619 8829
rect 7561 8789 7573 8823
rect 7607 8789 7619 8823
rect 7561 8783 7619 8789
rect 7650 8780 7656 8832
rect 7708 8820 7714 8832
rect 7834 8820 7840 8832
rect 7708 8792 7840 8820
rect 7708 8780 7714 8792
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 8573 8823 8631 8829
rect 8573 8789 8585 8823
rect 8619 8820 8631 8823
rect 8662 8820 8668 8832
rect 8619 8792 8668 8820
rect 8619 8789 8631 8792
rect 8573 8783 8631 8789
rect 8662 8780 8668 8792
rect 8720 8820 8726 8832
rect 9646 8820 9674 8860
rect 10686 8820 10692 8832
rect 8720 8792 9674 8820
rect 10647 8792 10692 8820
rect 8720 8780 8726 8792
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 11146 8780 11152 8832
rect 11204 8820 11210 8832
rect 11517 8823 11575 8829
rect 11517 8820 11529 8823
rect 11204 8792 11529 8820
rect 11204 8780 11210 8792
rect 11517 8789 11529 8792
rect 11563 8789 11575 8823
rect 12084 8820 12112 8860
rect 16390 8848 16396 8900
rect 16448 8888 16454 8900
rect 17129 8891 17187 8897
rect 16448 8860 17080 8888
rect 16448 8848 16454 8860
rect 12345 8823 12403 8829
rect 12345 8820 12357 8823
rect 12084 8792 12357 8820
rect 11517 8783 11575 8789
rect 12345 8789 12357 8792
rect 12391 8820 12403 8823
rect 13633 8823 13691 8829
rect 13633 8820 13645 8823
rect 12391 8792 13645 8820
rect 12391 8789 12403 8792
rect 12345 8783 12403 8789
rect 13633 8789 13645 8792
rect 13679 8820 13691 8823
rect 13814 8820 13820 8832
rect 13679 8792 13820 8820
rect 13679 8789 13691 8792
rect 13633 8783 13691 8789
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 14829 8823 14887 8829
rect 14829 8789 14841 8823
rect 14875 8820 14887 8823
rect 15194 8820 15200 8832
rect 14875 8792 15200 8820
rect 14875 8789 14887 8792
rect 14829 8783 14887 8789
rect 15194 8780 15200 8792
rect 15252 8820 15258 8832
rect 15378 8820 15384 8832
rect 15252 8792 15384 8820
rect 15252 8780 15258 8792
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 15562 8780 15568 8832
rect 15620 8820 15626 8832
rect 16025 8823 16083 8829
rect 16025 8820 16037 8823
rect 15620 8792 16037 8820
rect 15620 8780 15626 8792
rect 16025 8789 16037 8792
rect 16071 8789 16083 8823
rect 16025 8783 16083 8789
rect 16117 8823 16175 8829
rect 16117 8789 16129 8823
rect 16163 8820 16175 8823
rect 16298 8820 16304 8832
rect 16163 8792 16304 8820
rect 16163 8789 16175 8792
rect 16117 8783 16175 8789
rect 16298 8780 16304 8792
rect 16356 8780 16362 8832
rect 16485 8823 16543 8829
rect 16485 8789 16497 8823
rect 16531 8820 16543 8823
rect 16942 8820 16948 8832
rect 16531 8792 16948 8820
rect 16531 8789 16543 8792
rect 16485 8783 16543 8789
rect 16942 8780 16948 8792
rect 17000 8780 17006 8832
rect 17052 8820 17080 8860
rect 17129 8857 17141 8891
rect 17175 8888 17187 8891
rect 19352 8888 19380 8928
rect 20806 8916 20812 8928
rect 20864 8916 20870 8968
rect 19518 8888 19524 8900
rect 17175 8860 19380 8888
rect 19479 8860 19524 8888
rect 17175 8857 17187 8860
rect 17129 8851 17187 8857
rect 19518 8848 19524 8860
rect 19576 8848 19582 8900
rect 22278 8888 22284 8900
rect 20824 8860 22284 8888
rect 18785 8823 18843 8829
rect 18785 8820 18797 8823
rect 17052 8792 18797 8820
rect 18785 8789 18797 8792
rect 18831 8820 18843 8823
rect 18874 8820 18880 8832
rect 18831 8792 18880 8820
rect 18831 8789 18843 8792
rect 18785 8783 18843 8789
rect 18874 8780 18880 8792
rect 18932 8780 18938 8832
rect 20824 8829 20852 8860
rect 22278 8848 22284 8860
rect 22336 8848 22342 8900
rect 20809 8823 20867 8829
rect 20809 8789 20821 8823
rect 20855 8789 20867 8823
rect 20809 8783 20867 8789
rect 20898 8780 20904 8832
rect 20956 8820 20962 8832
rect 20956 8792 21001 8820
rect 20956 8780 20962 8792
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 9398 8576 9404 8628
rect 9456 8616 9462 8628
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 9456 8588 9505 8616
rect 9456 8576 9462 8588
rect 9493 8585 9505 8588
rect 9539 8585 9551 8619
rect 10134 8616 10140 8628
rect 10095 8588 10140 8616
rect 9493 8579 9551 8585
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 12802 8576 12808 8628
rect 12860 8616 12866 8628
rect 13081 8619 13139 8625
rect 13081 8616 13093 8619
rect 12860 8588 13093 8616
rect 12860 8576 12866 8588
rect 13081 8585 13093 8588
rect 13127 8616 13139 8619
rect 13538 8616 13544 8628
rect 13127 8588 13544 8616
rect 13127 8585 13139 8588
rect 13081 8579 13139 8585
rect 13538 8576 13544 8588
rect 13596 8616 13602 8628
rect 13633 8619 13691 8625
rect 13633 8616 13645 8619
rect 13596 8588 13645 8616
rect 13596 8576 13602 8588
rect 13633 8585 13645 8588
rect 13679 8585 13691 8619
rect 15194 8616 15200 8628
rect 15155 8588 15200 8616
rect 13633 8579 13691 8585
rect 15194 8576 15200 8588
rect 15252 8576 15258 8628
rect 15565 8619 15623 8625
rect 15565 8585 15577 8619
rect 15611 8616 15623 8619
rect 15930 8616 15936 8628
rect 15611 8588 15936 8616
rect 15611 8585 15623 8588
rect 15565 8579 15623 8585
rect 15930 8576 15936 8588
rect 15988 8576 15994 8628
rect 16942 8616 16948 8628
rect 16903 8588 16948 8616
rect 16942 8576 16948 8588
rect 17000 8576 17006 8628
rect 17034 8576 17040 8628
rect 17092 8616 17098 8628
rect 17405 8619 17463 8625
rect 17092 8588 17137 8616
rect 17092 8576 17098 8588
rect 17405 8585 17417 8619
rect 17451 8585 17463 8619
rect 17405 8579 17463 8585
rect 17773 8619 17831 8625
rect 17773 8585 17785 8619
rect 17819 8616 17831 8619
rect 17954 8616 17960 8628
rect 17819 8588 17960 8616
rect 17819 8585 17831 8588
rect 17773 8579 17831 8585
rect 4982 8508 4988 8560
rect 5040 8548 5046 8560
rect 7285 8551 7343 8557
rect 5040 8520 6868 8548
rect 5040 8508 5046 8520
rect 5350 8412 5356 8424
rect 5311 8384 5356 8412
rect 5350 8372 5356 8384
rect 5408 8372 5414 8424
rect 5534 8372 5540 8424
rect 5592 8412 5598 8424
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 5592 8384 6377 8412
rect 5592 8372 5598 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 6840 8412 6868 8520
rect 7285 8517 7297 8551
rect 7331 8548 7343 8551
rect 7929 8551 7987 8557
rect 7929 8548 7941 8551
rect 7331 8520 7941 8548
rect 7331 8517 7343 8520
rect 7285 8511 7343 8517
rect 7929 8517 7941 8520
rect 7975 8548 7987 8551
rect 8662 8548 8668 8560
rect 7975 8520 8668 8548
rect 7975 8517 7987 8520
rect 7929 8511 7987 8517
rect 8662 8508 8668 8520
rect 8720 8508 8726 8560
rect 8772 8520 9674 8548
rect 7377 8483 7435 8489
rect 7377 8449 7389 8483
rect 7423 8480 7435 8483
rect 8389 8483 8447 8489
rect 8389 8480 8401 8483
rect 7423 8452 8401 8480
rect 7423 8449 7435 8452
rect 7377 8443 7435 8449
rect 8389 8449 8401 8452
rect 8435 8480 8447 8483
rect 8772 8480 8800 8520
rect 8435 8452 8800 8480
rect 9646 8480 9674 8520
rect 9766 8508 9772 8560
rect 9824 8548 9830 8560
rect 10505 8551 10563 8557
rect 10505 8548 10517 8551
rect 9824 8520 10517 8548
rect 9824 8508 9830 8520
rect 10505 8517 10517 8520
rect 10551 8517 10563 8551
rect 14274 8548 14280 8560
rect 10505 8511 10563 8517
rect 13556 8520 14280 8548
rect 11974 8480 11980 8492
rect 9646 8452 11980 8480
rect 8435 8449 8447 8452
rect 8389 8443 8447 8449
rect 11974 8440 11980 8452
rect 12032 8480 12038 8492
rect 12032 8452 13400 8480
rect 12032 8440 12038 8452
rect 7469 8415 7527 8421
rect 7469 8412 7481 8415
rect 6840 8384 7481 8412
rect 6365 8375 6423 8381
rect 7469 8381 7481 8384
rect 7515 8381 7527 8415
rect 7469 8375 7527 8381
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8412 9643 8415
rect 9674 8412 9680 8424
rect 9631 8384 9680 8412
rect 9631 8381 9643 8384
rect 9585 8375 9643 8381
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 9769 8415 9827 8421
rect 9769 8381 9781 8415
rect 9815 8412 9827 8415
rect 10594 8412 10600 8424
rect 9815 8384 9904 8412
rect 10555 8384 10600 8412
rect 9815 8381 9827 8384
rect 9769 8375 9827 8381
rect 5258 8304 5264 8356
rect 5316 8344 5322 8356
rect 5316 8316 9674 8344
rect 5316 8304 5322 8316
rect 6914 8276 6920 8288
rect 6875 8248 6920 8276
rect 6914 8236 6920 8248
rect 6972 8236 6978 8288
rect 9122 8276 9128 8288
rect 9083 8248 9128 8276
rect 9122 8236 9128 8248
rect 9180 8236 9186 8288
rect 9646 8276 9674 8316
rect 9876 8276 9904 8384
rect 10594 8372 10600 8384
rect 10652 8372 10658 8424
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8412 10839 8415
rect 10870 8412 10876 8424
rect 10827 8384 10876 8412
rect 10827 8381 10839 8384
rect 10781 8375 10839 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 10962 8372 10968 8424
rect 11020 8412 11026 8424
rect 12437 8415 12495 8421
rect 12437 8412 12449 8415
rect 11020 8384 12449 8412
rect 11020 8372 11026 8384
rect 12437 8381 12449 8384
rect 12483 8412 12495 8415
rect 13262 8412 13268 8424
rect 12483 8384 13268 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 11882 8304 11888 8356
rect 11940 8344 11946 8356
rect 11977 8347 12035 8353
rect 11977 8344 11989 8347
rect 11940 8316 11989 8344
rect 11940 8304 11946 8316
rect 11977 8313 11989 8316
rect 12023 8344 12035 8347
rect 12023 8316 12434 8344
rect 12023 8313 12035 8316
rect 11977 8307 12035 8313
rect 9646 8248 9904 8276
rect 11238 8236 11244 8288
rect 11296 8276 11302 8288
rect 11609 8279 11667 8285
rect 11609 8276 11621 8279
rect 11296 8248 11621 8276
rect 11296 8236 11302 8248
rect 11609 8245 11621 8248
rect 11655 8245 11667 8279
rect 12406 8276 12434 8316
rect 12526 8276 12532 8288
rect 12406 8248 12532 8276
rect 11609 8239 11667 8245
rect 12526 8236 12532 8248
rect 12584 8236 12590 8288
rect 13372 8276 13400 8452
rect 13556 8421 13584 8520
rect 14274 8508 14280 8520
rect 14332 8508 14338 8560
rect 16022 8548 16028 8560
rect 15983 8520 16028 8548
rect 16022 8508 16028 8520
rect 16080 8508 16086 8560
rect 16850 8548 16856 8560
rect 16316 8520 16856 8548
rect 16316 8489 16344 8520
rect 16850 8508 16856 8520
rect 16908 8508 16914 8560
rect 17420 8548 17448 8579
rect 17954 8576 17960 8588
rect 18012 8576 18018 8628
rect 18138 8616 18144 8628
rect 18099 8588 18144 8616
rect 18138 8576 18144 8588
rect 18196 8576 18202 8628
rect 18414 8576 18420 8628
rect 18472 8616 18478 8628
rect 19153 8619 19211 8625
rect 19153 8616 19165 8619
rect 18472 8588 19165 8616
rect 18472 8576 18478 8588
rect 19153 8585 19165 8588
rect 19199 8585 19211 8619
rect 19153 8579 19211 8585
rect 19610 8576 19616 8628
rect 19668 8616 19674 8628
rect 19705 8619 19763 8625
rect 19705 8616 19717 8619
rect 19668 8588 19717 8616
rect 19668 8576 19674 8588
rect 19705 8585 19717 8588
rect 19751 8585 19763 8619
rect 20254 8616 20260 8628
rect 20215 8588 20260 8616
rect 19705 8579 19763 8585
rect 20254 8576 20260 8588
rect 20312 8576 20318 8628
rect 20625 8619 20683 8625
rect 20625 8585 20637 8619
rect 20671 8616 20683 8619
rect 20898 8616 20904 8628
rect 20671 8588 20904 8616
rect 20671 8585 20683 8588
rect 20625 8579 20683 8585
rect 20898 8576 20904 8588
rect 20956 8576 20962 8628
rect 20990 8576 20996 8628
rect 21048 8616 21054 8628
rect 21174 8616 21180 8628
rect 21048 8588 21180 8616
rect 21048 8576 21054 8588
rect 21174 8576 21180 8588
rect 21232 8576 21238 8628
rect 17420 8520 18184 8548
rect 13725 8483 13783 8489
rect 13725 8449 13737 8483
rect 13771 8449 13783 8483
rect 13725 8443 13783 8449
rect 16301 8483 16359 8489
rect 16301 8449 16313 8483
rect 16347 8449 16359 8483
rect 18156 8480 18184 8520
rect 18230 8508 18236 8560
rect 18288 8548 18294 8560
rect 18509 8551 18567 8557
rect 18509 8548 18521 8551
rect 18288 8520 18521 8548
rect 18288 8508 18294 8520
rect 18509 8517 18521 8520
rect 18555 8548 18567 8551
rect 18690 8548 18696 8560
rect 18555 8520 18696 8548
rect 18555 8517 18567 8520
rect 18509 8511 18567 8517
rect 18690 8508 18696 8520
rect 18748 8508 18754 8560
rect 18322 8480 18328 8492
rect 18156 8452 18328 8480
rect 16301 8443 16359 8449
rect 13541 8415 13599 8421
rect 13541 8381 13553 8415
rect 13587 8381 13599 8415
rect 13541 8375 13599 8381
rect 13740 8344 13768 8443
rect 18322 8440 18328 8452
rect 18380 8440 18386 8492
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8480 18659 8483
rect 18782 8480 18788 8492
rect 18647 8452 18788 8480
rect 18647 8449 18659 8452
rect 18601 8443 18659 8449
rect 18782 8440 18788 8452
rect 18840 8440 18846 8492
rect 19518 8480 19524 8492
rect 19479 8452 19524 8480
rect 19518 8440 19524 8452
rect 19576 8440 19582 8492
rect 19978 8440 19984 8492
rect 20036 8480 20042 8492
rect 20073 8483 20131 8489
rect 20073 8480 20085 8483
rect 20036 8452 20085 8480
rect 20036 8440 20042 8452
rect 20073 8449 20085 8452
rect 20119 8449 20131 8483
rect 20073 8443 20131 8449
rect 20898 8440 20904 8492
rect 20956 8480 20962 8492
rect 20993 8483 21051 8489
rect 20993 8480 21005 8483
rect 20956 8452 21005 8480
rect 20956 8440 20962 8452
rect 20993 8449 21005 8452
rect 21039 8449 21051 8483
rect 20993 8443 21051 8449
rect 13906 8372 13912 8424
rect 13964 8412 13970 8424
rect 15194 8412 15200 8424
rect 13964 8384 15200 8412
rect 13964 8372 13970 8384
rect 15194 8372 15200 8384
rect 15252 8372 15258 8424
rect 16853 8415 16911 8421
rect 16853 8381 16865 8415
rect 16899 8412 16911 8415
rect 17218 8412 17224 8424
rect 16899 8384 17224 8412
rect 16899 8381 16911 8384
rect 16853 8375 16911 8381
rect 17218 8372 17224 8384
rect 17276 8372 17282 8424
rect 18693 8415 18751 8421
rect 18693 8381 18705 8415
rect 18739 8381 18751 8415
rect 18693 8375 18751 8381
rect 21085 8415 21143 8421
rect 21085 8381 21097 8415
rect 21131 8412 21143 8415
rect 21174 8412 21180 8424
rect 21131 8384 21180 8412
rect 21131 8381 21143 8384
rect 21085 8375 21143 8381
rect 14369 8347 14427 8353
rect 14369 8344 14381 8347
rect 13740 8316 14381 8344
rect 13538 8276 13544 8288
rect 13372 8248 13544 8276
rect 13538 8236 13544 8248
rect 13596 8276 13602 8288
rect 13740 8276 13768 8316
rect 14369 8313 14381 8316
rect 14415 8313 14427 8347
rect 14826 8344 14832 8356
rect 14787 8316 14832 8344
rect 14369 8307 14427 8313
rect 14826 8304 14832 8316
rect 14884 8304 14890 8356
rect 15378 8304 15384 8356
rect 15436 8344 15442 8356
rect 15436 8316 16574 8344
rect 15436 8304 15442 8316
rect 13596 8248 13768 8276
rect 14093 8279 14151 8285
rect 13596 8236 13602 8248
rect 14093 8245 14105 8279
rect 14139 8276 14151 8279
rect 14274 8276 14280 8288
rect 14139 8248 14280 8276
rect 14139 8245 14151 8248
rect 14093 8239 14151 8245
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 16546 8276 16574 8316
rect 18506 8304 18512 8356
rect 18564 8344 18570 8356
rect 18708 8344 18736 8375
rect 21174 8372 21180 8384
rect 21232 8372 21238 8424
rect 21269 8415 21327 8421
rect 21269 8381 21281 8415
rect 21315 8412 21327 8415
rect 21450 8412 21456 8424
rect 21315 8384 21456 8412
rect 21315 8381 21327 8384
rect 21269 8375 21327 8381
rect 21450 8372 21456 8384
rect 21508 8372 21514 8424
rect 18564 8316 18736 8344
rect 18564 8304 18570 8316
rect 18322 8276 18328 8288
rect 16546 8248 18328 8276
rect 18322 8236 18328 8248
rect 18380 8236 18386 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 6730 8032 6736 8084
rect 6788 8072 6794 8084
rect 6825 8075 6883 8081
rect 6825 8072 6837 8075
rect 6788 8044 6837 8072
rect 6788 8032 6794 8044
rect 6825 8041 6837 8044
rect 6871 8041 6883 8075
rect 6825 8035 6883 8041
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 7800 8044 8953 8072
rect 7800 8032 7806 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 10134 8072 10140 8084
rect 10095 8044 10140 8072
rect 8941 8035 8999 8041
rect 10134 8032 10140 8044
rect 10192 8032 10198 8084
rect 10318 8032 10324 8084
rect 10376 8072 10382 8084
rect 10873 8075 10931 8081
rect 10873 8072 10885 8075
rect 10376 8044 10885 8072
rect 10376 8032 10382 8044
rect 10873 8041 10885 8044
rect 10919 8041 10931 8075
rect 10873 8035 10931 8041
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 12897 8075 12955 8081
rect 12897 8072 12909 8075
rect 12676 8044 12909 8072
rect 12676 8032 12682 8044
rect 12897 8041 12909 8044
rect 12943 8041 12955 8075
rect 13722 8072 13728 8084
rect 13683 8044 13728 8072
rect 12897 8035 12955 8041
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 14550 8032 14556 8084
rect 14608 8072 14614 8084
rect 15378 8072 15384 8084
rect 14608 8044 15384 8072
rect 14608 8032 14614 8044
rect 15378 8032 15384 8044
rect 15436 8032 15442 8084
rect 16850 8032 16856 8084
rect 16908 8072 16914 8084
rect 18049 8075 18107 8081
rect 18049 8072 18061 8075
rect 16908 8044 18061 8072
rect 16908 8032 16914 8044
rect 18049 8041 18061 8044
rect 18095 8041 18107 8075
rect 18049 8035 18107 8041
rect 21085 8075 21143 8081
rect 21085 8041 21097 8075
rect 21131 8072 21143 8075
rect 21358 8072 21364 8084
rect 21131 8044 21364 8072
rect 21131 8041 21143 8044
rect 21085 8035 21143 8041
rect 21358 8032 21364 8044
rect 21416 8032 21422 8084
rect 8662 7964 8668 8016
rect 8720 8004 8726 8016
rect 10410 8004 10416 8016
rect 8720 7976 10416 8004
rect 8720 7964 8726 7976
rect 10410 7964 10416 7976
rect 10468 8004 10474 8016
rect 10962 8004 10968 8016
rect 10468 7976 10968 8004
rect 10468 7964 10474 7976
rect 10962 7964 10968 7976
rect 11020 8004 11026 8016
rect 11020 7976 11376 8004
rect 11020 7964 11026 7976
rect 5258 7936 5264 7948
rect 5219 7908 5264 7936
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 5994 7896 6000 7948
rect 6052 7936 6058 7948
rect 6181 7939 6239 7945
rect 6181 7936 6193 7939
rect 6052 7908 6193 7936
rect 6052 7896 6058 7908
rect 6181 7905 6193 7908
rect 6227 7905 6239 7939
rect 6181 7899 6239 7905
rect 6365 7939 6423 7945
rect 6365 7905 6377 7939
rect 6411 7936 6423 7939
rect 6914 7936 6920 7948
rect 6411 7908 6920 7936
rect 6411 7905 6423 7908
rect 6365 7899 6423 7905
rect 6914 7896 6920 7908
rect 6972 7896 6978 7948
rect 9122 7896 9128 7948
rect 9180 7936 9186 7948
rect 9401 7939 9459 7945
rect 9401 7936 9413 7939
rect 9180 7908 9413 7936
rect 9180 7896 9186 7908
rect 9401 7905 9413 7908
rect 9447 7905 9459 7939
rect 9582 7936 9588 7948
rect 9543 7908 9588 7936
rect 9401 7899 9459 7905
rect 9582 7896 9588 7908
rect 9640 7896 9646 7948
rect 11348 7945 11376 7976
rect 12434 7964 12440 8016
rect 12492 8004 12498 8016
rect 13265 8007 13323 8013
rect 13265 8004 13277 8007
rect 12492 7976 13277 8004
rect 12492 7964 12498 7976
rect 13265 7973 13277 7976
rect 13311 8004 13323 8007
rect 16206 8004 16212 8016
rect 13311 7976 16212 8004
rect 13311 7973 13323 7976
rect 13265 7967 13323 7973
rect 16206 7964 16212 7976
rect 16264 7964 16270 8016
rect 17954 7964 17960 8016
rect 18012 8004 18018 8016
rect 22186 8004 22192 8016
rect 18012 7976 22192 8004
rect 18012 7964 18018 7976
rect 22186 7964 22192 7976
rect 22244 7964 22250 8016
rect 11333 7939 11391 7945
rect 11333 7905 11345 7939
rect 11379 7905 11391 7939
rect 11333 7899 11391 7905
rect 11517 7939 11575 7945
rect 11517 7905 11529 7939
rect 11563 7936 11575 7939
rect 12158 7936 12164 7948
rect 11563 7908 12164 7936
rect 11563 7905 11575 7908
rect 11517 7899 11575 7905
rect 12158 7896 12164 7908
rect 12216 7896 12222 7948
rect 12345 7939 12403 7945
rect 12345 7905 12357 7939
rect 12391 7936 12403 7939
rect 12710 7936 12716 7948
rect 12391 7908 12716 7936
rect 12391 7905 12403 7908
rect 12345 7899 12403 7905
rect 12710 7896 12716 7908
rect 12768 7896 12774 7948
rect 14277 7939 14335 7945
rect 14277 7905 14289 7939
rect 14323 7936 14335 7939
rect 14366 7936 14372 7948
rect 14323 7908 14372 7936
rect 14323 7905 14335 7908
rect 14277 7899 14335 7905
rect 14366 7896 14372 7908
rect 14424 7896 14430 7948
rect 17037 7939 17095 7945
rect 17037 7936 17049 7939
rect 14476 7908 17049 7936
rect 5445 7871 5503 7877
rect 5445 7837 5457 7871
rect 5491 7868 5503 7871
rect 5534 7868 5540 7880
rect 5491 7840 5540 7868
rect 5491 7837 5503 7840
rect 5445 7831 5503 7837
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 12526 7868 12532 7880
rect 12487 7840 12532 7868
rect 12526 7828 12532 7840
rect 12584 7828 12590 7880
rect 14476 7868 14504 7908
rect 17037 7905 17049 7908
rect 17083 7905 17095 7939
rect 17037 7899 17095 7905
rect 17221 7939 17279 7945
rect 17221 7905 17233 7939
rect 17267 7936 17279 7939
rect 17494 7936 17500 7948
rect 17267 7908 17500 7936
rect 17267 7905 17279 7908
rect 17221 7899 17279 7905
rect 17494 7896 17500 7908
rect 17552 7896 17558 7948
rect 18690 7936 18696 7948
rect 18651 7908 18696 7936
rect 18690 7896 18696 7908
rect 18748 7896 18754 7948
rect 20441 7939 20499 7945
rect 20441 7905 20453 7939
rect 20487 7936 20499 7939
rect 20714 7936 20720 7948
rect 20487 7908 20720 7936
rect 20487 7905 20499 7908
rect 20441 7899 20499 7905
rect 20714 7896 20720 7908
rect 20772 7896 20778 7948
rect 13372 7840 14504 7868
rect 9309 7803 9367 7809
rect 9309 7800 9321 7803
rect 5828 7772 9321 7800
rect 4246 7692 4252 7744
rect 4304 7732 4310 7744
rect 4709 7735 4767 7741
rect 4709 7732 4721 7735
rect 4304 7704 4721 7732
rect 4304 7692 4310 7704
rect 4709 7701 4721 7704
rect 4755 7732 4767 7735
rect 5353 7735 5411 7741
rect 5353 7732 5365 7735
rect 4755 7704 5365 7732
rect 4755 7701 4767 7704
rect 4709 7695 4767 7701
rect 5353 7701 5365 7704
rect 5399 7732 5411 7735
rect 5442 7732 5448 7744
rect 5399 7704 5448 7732
rect 5399 7701 5411 7704
rect 5353 7695 5411 7701
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 5828 7741 5856 7772
rect 9309 7769 9321 7772
rect 9355 7769 9367 7803
rect 9309 7763 9367 7769
rect 10686 7760 10692 7812
rect 10744 7800 10750 7812
rect 12434 7800 12440 7812
rect 10744 7772 12440 7800
rect 10744 7760 10750 7772
rect 12434 7760 12440 7772
rect 12492 7760 12498 7812
rect 12618 7760 12624 7812
rect 12676 7800 12682 7812
rect 13372 7800 13400 7840
rect 14918 7828 14924 7880
rect 14976 7868 14982 7880
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 14976 7840 19257 7868
rect 14976 7828 14982 7840
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 20162 7868 20168 7880
rect 20123 7840 20168 7868
rect 19245 7831 19303 7837
rect 20162 7828 20168 7840
rect 20220 7828 20226 7880
rect 20806 7828 20812 7880
rect 20864 7868 20870 7880
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 20864 7840 20913 7868
rect 20864 7828 20870 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 12676 7772 13400 7800
rect 12676 7760 12682 7772
rect 13722 7760 13728 7812
rect 13780 7800 13786 7812
rect 14369 7803 14427 7809
rect 14369 7800 14381 7803
rect 13780 7772 14381 7800
rect 13780 7760 13786 7772
rect 14369 7769 14381 7772
rect 14415 7769 14427 7803
rect 14369 7763 14427 7769
rect 14461 7803 14519 7809
rect 14461 7769 14473 7803
rect 14507 7800 14519 7803
rect 15105 7803 15163 7809
rect 15105 7800 15117 7803
rect 14507 7772 15117 7800
rect 14507 7769 14519 7772
rect 14461 7763 14519 7769
rect 15105 7769 15117 7772
rect 15151 7769 15163 7803
rect 15105 7763 15163 7769
rect 16945 7803 17003 7809
rect 16945 7769 16957 7803
rect 16991 7800 17003 7803
rect 17126 7800 17132 7812
rect 16991 7772 17132 7800
rect 16991 7769 17003 7772
rect 16945 7763 17003 7769
rect 17126 7760 17132 7772
rect 17184 7760 17190 7812
rect 19518 7800 19524 7812
rect 19479 7772 19524 7800
rect 19518 7760 19524 7772
rect 19576 7760 19582 7812
rect 5813 7735 5871 7741
rect 5813 7701 5825 7735
rect 5859 7701 5871 7735
rect 5813 7695 5871 7701
rect 5902 7692 5908 7744
rect 5960 7732 5966 7744
rect 6457 7735 6515 7741
rect 6457 7732 6469 7735
rect 5960 7704 6469 7732
rect 5960 7692 5966 7704
rect 6457 7701 6469 7704
rect 6503 7701 6515 7735
rect 6457 7695 6515 7701
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 10505 7735 10563 7741
rect 10505 7732 10517 7735
rect 8720 7704 10517 7732
rect 8720 7692 8726 7704
rect 10505 7701 10517 7704
rect 10551 7732 10563 7735
rect 11241 7735 11299 7741
rect 11241 7732 11253 7735
rect 10551 7704 11253 7732
rect 10551 7701 10563 7704
rect 10505 7695 10563 7701
rect 11241 7701 11253 7704
rect 11287 7701 11299 7735
rect 11241 7695 11299 7701
rect 11974 7692 11980 7744
rect 12032 7732 12038 7744
rect 12158 7732 12164 7744
rect 12032 7704 12164 7732
rect 12032 7692 12038 7704
rect 12158 7692 12164 7704
rect 12216 7692 12222 7744
rect 13078 7692 13084 7744
rect 13136 7732 13142 7744
rect 13446 7732 13452 7744
rect 13136 7704 13452 7732
rect 13136 7692 13142 7704
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 14550 7692 14556 7744
rect 14608 7732 14614 7744
rect 14829 7735 14887 7741
rect 14829 7732 14841 7735
rect 14608 7704 14841 7732
rect 14608 7692 14614 7704
rect 14829 7701 14841 7704
rect 14875 7701 14887 7735
rect 14829 7695 14887 7701
rect 15841 7735 15899 7741
rect 15841 7701 15853 7735
rect 15887 7732 15899 7735
rect 15930 7732 15936 7744
rect 15887 7704 15936 7732
rect 15887 7701 15899 7704
rect 15841 7695 15899 7701
rect 15930 7692 15936 7704
rect 15988 7692 15994 7744
rect 16298 7732 16304 7744
rect 16259 7704 16304 7732
rect 16298 7692 16304 7704
rect 16356 7692 16362 7744
rect 16390 7692 16396 7744
rect 16448 7732 16454 7744
rect 16577 7735 16635 7741
rect 16577 7732 16589 7735
rect 16448 7704 16589 7732
rect 16448 7692 16454 7704
rect 16577 7701 16589 7704
rect 16623 7701 16635 7735
rect 17770 7732 17776 7744
rect 17731 7704 17776 7732
rect 16577 7695 16635 7701
rect 17770 7692 17776 7704
rect 17828 7692 17834 7744
rect 18414 7732 18420 7744
rect 18375 7704 18420 7732
rect 18414 7692 18420 7704
rect 18472 7692 18478 7744
rect 18506 7692 18512 7744
rect 18564 7732 18570 7744
rect 18564 7704 18609 7732
rect 18564 7692 18570 7704
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 5261 7531 5319 7537
rect 5261 7497 5273 7531
rect 5307 7528 5319 7531
rect 5350 7528 5356 7540
rect 5307 7500 5356 7528
rect 5307 7497 5319 7500
rect 5261 7491 5319 7497
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 5629 7531 5687 7537
rect 5629 7497 5641 7531
rect 5675 7528 5687 7531
rect 5902 7528 5908 7540
rect 5675 7500 5908 7528
rect 5675 7497 5687 7500
rect 5629 7491 5687 7497
rect 5902 7488 5908 7500
rect 5960 7488 5966 7540
rect 7101 7531 7159 7537
rect 7101 7497 7113 7531
rect 7147 7528 7159 7531
rect 9582 7528 9588 7540
rect 7147 7500 9588 7528
rect 7147 7497 7159 7500
rect 7101 7491 7159 7497
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 9769 7531 9827 7537
rect 9769 7497 9781 7531
rect 9815 7528 9827 7531
rect 10594 7528 10600 7540
rect 9815 7500 10600 7528
rect 9815 7497 9827 7500
rect 9769 7491 9827 7497
rect 10594 7488 10600 7500
rect 10652 7488 10658 7540
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 11112 7500 11529 7528
rect 11112 7488 11118 7500
rect 11517 7497 11529 7500
rect 11563 7497 11575 7531
rect 11974 7528 11980 7540
rect 11935 7500 11980 7528
rect 11517 7491 11575 7497
rect 11974 7488 11980 7500
rect 12032 7488 12038 7540
rect 12084 7500 13492 7528
rect 9398 7460 9404 7472
rect 6472 7432 6868 7460
rect 9359 7432 9404 7460
rect 4982 7324 4988 7336
rect 4943 7296 4988 7324
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 5166 7324 5172 7336
rect 5127 7296 5172 7324
rect 5166 7284 5172 7296
rect 5224 7284 5230 7336
rect 5718 7284 5724 7336
rect 5776 7324 5782 7336
rect 6472 7333 6500 7432
rect 6730 7392 6736 7404
rect 6691 7364 6736 7392
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 6457 7327 6515 7333
rect 6457 7324 6469 7327
rect 5776 7296 6469 7324
rect 5776 7284 5782 7296
rect 6457 7293 6469 7296
rect 6503 7293 6515 7327
rect 6638 7324 6644 7336
rect 6599 7296 6644 7324
rect 6457 7287 6515 7293
rect 6638 7284 6644 7296
rect 6696 7284 6702 7336
rect 6840 7324 6868 7432
rect 9398 7420 9404 7432
rect 9456 7460 9462 7472
rect 10134 7460 10140 7472
rect 9456 7432 10140 7460
rect 9456 7420 9462 7432
rect 10134 7420 10140 7432
rect 10192 7420 10198 7472
rect 10505 7463 10563 7469
rect 10505 7429 10517 7463
rect 10551 7460 10563 7463
rect 10686 7460 10692 7472
rect 10551 7432 10692 7460
rect 10551 7429 10563 7432
rect 10505 7423 10563 7429
rect 8202 7352 8208 7404
rect 8260 7392 8266 7404
rect 9309 7395 9367 7401
rect 8260 7364 9260 7392
rect 8260 7352 8266 7364
rect 9125 7327 9183 7333
rect 9125 7324 9137 7327
rect 6840 7296 9137 7324
rect 9125 7293 9137 7296
rect 9171 7293 9183 7327
rect 9232 7324 9260 7364
rect 9309 7361 9321 7395
rect 9355 7392 9367 7395
rect 10520 7392 10548 7423
rect 10686 7420 10692 7432
rect 10744 7420 10750 7472
rect 12084 7460 12112 7500
rect 10980 7432 12112 7460
rect 9355 7364 10548 7392
rect 9355 7361 9367 7364
rect 9309 7355 9367 7361
rect 10980 7324 11008 7432
rect 12158 7420 12164 7472
rect 12216 7460 12222 7472
rect 13464 7469 13492 7500
rect 13630 7488 13636 7540
rect 13688 7528 13694 7540
rect 13909 7531 13967 7537
rect 13909 7528 13921 7531
rect 13688 7500 13921 7528
rect 13688 7488 13694 7500
rect 13909 7497 13921 7500
rect 13955 7497 13967 7531
rect 14550 7528 14556 7540
rect 14511 7500 14556 7528
rect 13909 7491 13967 7497
rect 14550 7488 14556 7500
rect 14608 7488 14614 7540
rect 14918 7528 14924 7540
rect 14879 7500 14924 7528
rect 14918 7488 14924 7500
rect 14976 7488 14982 7540
rect 16298 7488 16304 7540
rect 16356 7528 16362 7540
rect 17037 7531 17095 7537
rect 17037 7528 17049 7531
rect 16356 7500 17049 7528
rect 16356 7488 16362 7500
rect 17037 7497 17049 7500
rect 17083 7497 17095 7531
rect 17037 7491 17095 7497
rect 17770 7488 17776 7540
rect 17828 7528 17834 7540
rect 18233 7531 18291 7537
rect 18233 7528 18245 7531
rect 17828 7500 18245 7528
rect 17828 7488 17834 7500
rect 18233 7497 18245 7500
rect 18279 7497 18291 7531
rect 18233 7491 18291 7497
rect 18414 7488 18420 7540
rect 18472 7528 18478 7540
rect 18601 7531 18659 7537
rect 18601 7528 18613 7531
rect 18472 7500 18613 7528
rect 18472 7488 18478 7500
rect 18601 7497 18613 7500
rect 18647 7497 18659 7531
rect 18601 7491 18659 7497
rect 12529 7463 12587 7469
rect 12529 7460 12541 7463
rect 12216 7432 12541 7460
rect 12216 7420 12222 7432
rect 12529 7429 12541 7432
rect 12575 7429 12587 7463
rect 12529 7423 12587 7429
rect 13449 7463 13507 7469
rect 13449 7429 13461 7463
rect 13495 7460 13507 7463
rect 13495 7432 13860 7460
rect 13495 7429 13507 7432
rect 13449 7423 13507 7429
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 9232 7296 11008 7324
rect 11072 7364 11897 7392
rect 9125 7287 9183 7293
rect 2590 7216 2596 7268
rect 2648 7256 2654 7268
rect 11072 7265 11100 7364
rect 11885 7361 11897 7364
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 13078 7352 13084 7404
rect 13136 7392 13142 7404
rect 13541 7395 13599 7401
rect 13541 7392 13553 7395
rect 13136 7364 13553 7392
rect 13136 7352 13142 7364
rect 13541 7361 13553 7364
rect 13587 7361 13599 7395
rect 13832 7392 13860 7432
rect 14274 7420 14280 7472
rect 14332 7460 14338 7472
rect 14461 7463 14519 7469
rect 14461 7460 14473 7463
rect 14332 7432 14473 7460
rect 14332 7420 14338 7432
rect 14461 7429 14473 7432
rect 14507 7429 14519 7463
rect 14461 7423 14519 7429
rect 15657 7463 15715 7469
rect 15657 7429 15669 7463
rect 15703 7460 15715 7463
rect 16390 7460 16396 7472
rect 15703 7432 16396 7460
rect 15703 7429 15715 7432
rect 15657 7423 15715 7429
rect 16390 7420 16396 7432
rect 16448 7420 16454 7472
rect 19153 7463 19211 7469
rect 19153 7429 19165 7463
rect 19199 7460 19211 7463
rect 21082 7460 21088 7472
rect 19199 7432 21088 7460
rect 19199 7429 19211 7432
rect 19153 7423 19211 7429
rect 21082 7420 21088 7432
rect 21140 7420 21146 7472
rect 14826 7392 14832 7404
rect 13832 7364 14832 7392
rect 13541 7355 13599 7361
rect 14826 7352 14832 7364
rect 14884 7352 14890 7404
rect 15562 7392 15568 7404
rect 15523 7364 15568 7392
rect 15562 7352 15568 7364
rect 15620 7352 15626 7404
rect 17310 7392 17316 7404
rect 16776 7364 17316 7392
rect 12066 7324 12072 7336
rect 12027 7296 12072 7324
rect 12066 7284 12072 7296
rect 12124 7284 12130 7336
rect 13357 7327 13415 7333
rect 13357 7293 13369 7327
rect 13403 7324 13415 7327
rect 13814 7324 13820 7336
rect 13403 7296 13820 7324
rect 13403 7293 13415 7296
rect 13357 7287 13415 7293
rect 13814 7284 13820 7296
rect 13872 7284 13878 7336
rect 14369 7327 14427 7333
rect 14369 7293 14381 7327
rect 14415 7324 14427 7327
rect 14458 7324 14464 7336
rect 14415 7296 14464 7324
rect 14415 7293 14427 7296
rect 14369 7287 14427 7293
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 15838 7324 15844 7336
rect 15799 7296 15844 7324
rect 15838 7284 15844 7296
rect 15896 7284 15902 7336
rect 16776 7333 16804 7364
rect 17310 7352 17316 7364
rect 17368 7352 17374 7404
rect 17770 7352 17776 7404
rect 17828 7392 17834 7404
rect 18322 7392 18328 7404
rect 17828 7364 18328 7392
rect 17828 7352 17834 7364
rect 18322 7352 18328 7364
rect 18380 7352 18386 7404
rect 18877 7395 18935 7401
rect 18877 7361 18889 7395
rect 18923 7361 18935 7395
rect 18877 7355 18935 7361
rect 16761 7327 16819 7333
rect 16761 7293 16773 7327
rect 16807 7293 16819 7327
rect 16942 7324 16948 7336
rect 16903 7296 16948 7324
rect 16761 7287 16819 7293
rect 16942 7284 16948 7296
rect 17000 7284 17006 7336
rect 17954 7324 17960 7336
rect 17915 7296 17960 7324
rect 17954 7284 17960 7296
rect 18012 7284 18018 7336
rect 18138 7324 18144 7336
rect 18099 7296 18144 7324
rect 18138 7284 18144 7296
rect 18196 7284 18202 7336
rect 11057 7259 11115 7265
rect 11057 7256 11069 7259
rect 2648 7228 11069 7256
rect 2648 7216 2654 7228
rect 11057 7225 11069 7228
rect 11103 7225 11115 7259
rect 15197 7259 15255 7265
rect 15197 7256 15209 7259
rect 11057 7219 11115 7225
rect 12084 7228 12848 7256
rect 12084 7200 12112 7228
rect 4154 7148 4160 7200
rect 4212 7188 4218 7200
rect 4525 7191 4583 7197
rect 4525 7188 4537 7191
rect 4212 7160 4537 7188
rect 4212 7148 4218 7160
rect 4525 7157 4537 7160
rect 4571 7188 4583 7191
rect 5166 7188 5172 7200
rect 4571 7160 5172 7188
rect 4571 7157 4583 7160
rect 4525 7151 4583 7157
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 5902 7188 5908 7200
rect 5863 7160 5908 7188
rect 5902 7148 5908 7160
rect 5960 7188 5966 7200
rect 6638 7188 6644 7200
rect 5960 7160 6644 7188
rect 5960 7148 5966 7160
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 12066 7148 12072 7200
rect 12124 7148 12130 7200
rect 12820 7188 12848 7228
rect 13648 7228 15209 7256
rect 13648 7188 13676 7228
rect 15197 7225 15209 7228
rect 15243 7225 15255 7259
rect 15197 7219 15255 7225
rect 17405 7259 17463 7265
rect 17405 7225 17417 7259
rect 17451 7256 17463 7259
rect 18892 7256 18920 7355
rect 19518 7352 19524 7404
rect 19576 7392 19582 7404
rect 20165 7395 20223 7401
rect 20165 7392 20177 7395
rect 19576 7364 20177 7392
rect 19576 7352 19582 7364
rect 20165 7361 20177 7364
rect 20211 7361 20223 7395
rect 20714 7392 20720 7404
rect 20675 7364 20720 7392
rect 20165 7355 20223 7361
rect 20714 7352 20720 7364
rect 20772 7352 20778 7404
rect 19610 7324 19616 7336
rect 19571 7296 19616 7324
rect 19610 7284 19616 7296
rect 19668 7284 19674 7336
rect 20806 7284 20812 7336
rect 20864 7324 20870 7336
rect 20901 7327 20959 7333
rect 20901 7324 20913 7327
rect 20864 7296 20913 7324
rect 20864 7284 20870 7296
rect 20901 7293 20913 7296
rect 20947 7293 20959 7327
rect 20901 7287 20959 7293
rect 17451 7228 18920 7256
rect 17451 7225 17463 7228
rect 17405 7219 17463 7225
rect 12820 7160 13676 7188
rect 13814 7148 13820 7200
rect 13872 7188 13878 7200
rect 15654 7188 15660 7200
rect 13872 7160 15660 7188
rect 13872 7148 13878 7160
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 16206 7148 16212 7200
rect 16264 7188 16270 7200
rect 16301 7191 16359 7197
rect 16301 7188 16313 7191
rect 16264 7160 16313 7188
rect 16264 7148 16270 7160
rect 16301 7157 16313 7160
rect 16347 7188 16359 7191
rect 18322 7188 18328 7200
rect 16347 7160 18328 7188
rect 16347 7157 16359 7160
rect 16301 7151 16359 7157
rect 18322 7148 18328 7160
rect 18380 7148 18386 7200
rect 18598 7148 18604 7200
rect 18656 7188 18662 7200
rect 20349 7191 20407 7197
rect 20349 7188 20361 7191
rect 18656 7160 20361 7188
rect 18656 7148 18662 7160
rect 20349 7157 20361 7160
rect 20395 7157 20407 7191
rect 20349 7151 20407 7157
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 15562 6984 15568 6996
rect 8444 6956 15240 6984
rect 15523 6956 15568 6984
rect 8444 6944 8450 6956
rect 6638 6876 6644 6928
rect 6696 6916 6702 6928
rect 10870 6916 10876 6928
rect 6696 6888 10876 6916
rect 6696 6876 6702 6888
rect 10870 6876 10876 6888
rect 10928 6876 10934 6928
rect 13078 6876 13084 6928
rect 13136 6876 13142 6928
rect 15212 6916 15240 6956
rect 15562 6944 15568 6956
rect 15620 6944 15626 6996
rect 16942 6944 16948 6996
rect 17000 6984 17006 6996
rect 17313 6987 17371 6993
rect 17313 6984 17325 6987
rect 17000 6956 17325 6984
rect 17000 6944 17006 6956
rect 17313 6953 17325 6956
rect 17359 6953 17371 6987
rect 17313 6947 17371 6953
rect 18506 6944 18512 6996
rect 18564 6984 18570 6996
rect 18601 6987 18659 6993
rect 18601 6984 18613 6987
rect 18564 6956 18613 6984
rect 18564 6944 18570 6956
rect 18601 6953 18613 6956
rect 18647 6953 18659 6987
rect 18601 6947 18659 6953
rect 15930 6916 15936 6928
rect 15212 6888 15936 6916
rect 15930 6876 15936 6888
rect 15988 6876 15994 6928
rect 17494 6916 17500 6928
rect 16224 6888 17500 6916
rect 6181 6851 6239 6857
rect 6181 6817 6193 6851
rect 6227 6848 6239 6851
rect 6730 6848 6736 6860
rect 6227 6820 6736 6848
rect 6227 6817 6239 6820
rect 6181 6811 6239 6817
rect 6730 6808 6736 6820
rect 6788 6808 6794 6860
rect 9858 6808 9864 6860
rect 9916 6848 9922 6860
rect 10686 6848 10692 6860
rect 9916 6820 10692 6848
rect 9916 6808 9922 6820
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 11146 6848 11152 6860
rect 11107 6820 11152 6848
rect 11146 6808 11152 6820
rect 11204 6808 11210 6860
rect 11974 6848 11980 6860
rect 11935 6820 11980 6848
rect 11974 6808 11980 6820
rect 12032 6808 12038 6860
rect 12526 6808 12532 6860
rect 12584 6848 12590 6860
rect 12989 6851 13047 6857
rect 12989 6848 13001 6851
rect 12584 6820 13001 6848
rect 12584 6808 12590 6820
rect 12989 6817 13001 6820
rect 13035 6817 13047 6851
rect 13096 6848 13124 6876
rect 13265 6851 13323 6857
rect 13265 6848 13277 6851
rect 13096 6820 13277 6848
rect 12989 6811 13047 6817
rect 13265 6817 13277 6820
rect 13311 6817 13323 6851
rect 13265 6811 13323 6817
rect 13538 6808 13544 6860
rect 13596 6848 13602 6860
rect 14737 6851 14795 6857
rect 14737 6848 14749 6851
rect 13596 6820 14749 6848
rect 13596 6808 13602 6820
rect 14737 6817 14749 6820
rect 14783 6848 14795 6851
rect 15010 6848 15016 6860
rect 14783 6820 15016 6848
rect 14783 6817 14795 6820
rect 14737 6811 14795 6817
rect 15010 6808 15016 6820
rect 15068 6808 15074 6860
rect 16025 6851 16083 6857
rect 16025 6817 16037 6851
rect 16071 6848 16083 6851
rect 16114 6848 16120 6860
rect 16071 6820 16120 6848
rect 16071 6817 16083 6820
rect 16025 6811 16083 6817
rect 16114 6808 16120 6820
rect 16172 6808 16178 6860
rect 16224 6857 16252 6888
rect 17494 6876 17500 6888
rect 17552 6876 17558 6928
rect 16209 6851 16267 6857
rect 16209 6817 16221 6851
rect 16255 6817 16267 6851
rect 16209 6811 16267 6817
rect 16761 6851 16819 6857
rect 16761 6817 16773 6851
rect 16807 6848 16819 6851
rect 17678 6848 17684 6860
rect 16807 6820 17684 6848
rect 16807 6817 16819 6820
rect 16761 6811 16819 6817
rect 17678 6808 17684 6820
rect 17736 6808 17742 6860
rect 17954 6848 17960 6860
rect 17915 6820 17960 6848
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 19334 6848 19340 6860
rect 19247 6820 19340 6848
rect 19334 6808 19340 6820
rect 19392 6848 19398 6860
rect 19518 6848 19524 6860
rect 19392 6820 19524 6848
rect 19392 6808 19398 6820
rect 19518 6808 19524 6820
rect 19576 6808 19582 6860
rect 20438 6848 20444 6860
rect 20399 6820 20444 6848
rect 20438 6808 20444 6820
rect 20496 6808 20502 6860
rect 10594 6740 10600 6792
rect 10652 6780 10658 6792
rect 11238 6780 11244 6792
rect 10652 6752 11244 6780
rect 10652 6740 10658 6752
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 12069 6783 12127 6789
rect 12069 6749 12081 6783
rect 12115 6780 12127 6783
rect 16132 6780 16160 6808
rect 18046 6780 18052 6792
rect 12115 6752 13124 6780
rect 16132 6752 18052 6780
rect 12115 6749 12127 6752
rect 12069 6743 12127 6749
rect 9309 6715 9367 6721
rect 9309 6681 9321 6715
rect 9355 6712 9367 6715
rect 12710 6712 12716 6724
rect 9355 6684 12716 6712
rect 9355 6681 9367 6684
rect 9309 6675 9367 6681
rect 12710 6672 12716 6684
rect 12768 6672 12774 6724
rect 9585 6647 9643 6653
rect 9585 6613 9597 6647
rect 9631 6644 9643 6647
rect 9674 6644 9680 6656
rect 9631 6616 9680 6644
rect 9631 6613 9643 6616
rect 9585 6607 9643 6613
rect 9674 6604 9680 6616
rect 9732 6604 9738 6656
rect 10413 6647 10471 6653
rect 10413 6613 10425 6647
rect 10459 6644 10471 6647
rect 10594 6644 10600 6656
rect 10459 6616 10600 6644
rect 10459 6613 10471 6616
rect 10413 6607 10471 6613
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 10870 6604 10876 6656
rect 10928 6644 10934 6656
rect 11425 6647 11483 6653
rect 11425 6644 11437 6647
rect 10928 6616 11437 6644
rect 10928 6604 10934 6616
rect 11425 6613 11437 6616
rect 11471 6644 11483 6647
rect 12161 6647 12219 6653
rect 12161 6644 12173 6647
rect 11471 6616 12173 6644
rect 11471 6613 11483 6616
rect 11425 6607 11483 6613
rect 12161 6613 12173 6616
rect 12207 6613 12219 6647
rect 12161 6607 12219 6613
rect 12526 6604 12532 6656
rect 12584 6644 12590 6656
rect 13096 6644 13124 6752
rect 18046 6740 18052 6752
rect 18104 6740 18110 6792
rect 18141 6783 18199 6789
rect 18141 6749 18153 6783
rect 18187 6780 18199 6783
rect 20070 6780 20076 6792
rect 18187 6752 20076 6780
rect 18187 6749 18199 6752
rect 18141 6743 18199 6749
rect 20070 6740 20076 6752
rect 20128 6740 20134 6792
rect 20806 6780 20812 6792
rect 20767 6752 20812 6780
rect 20806 6740 20812 6752
rect 20864 6740 20870 6792
rect 13725 6715 13783 6721
rect 13725 6681 13737 6715
rect 13771 6712 13783 6715
rect 14274 6712 14280 6724
rect 13771 6684 14280 6712
rect 13771 6681 13783 6684
rect 13725 6675 13783 6681
rect 13740 6644 13768 6675
rect 14274 6672 14280 6684
rect 14332 6672 14338 6724
rect 14461 6715 14519 6721
rect 14461 6681 14473 6715
rect 14507 6712 14519 6715
rect 14918 6712 14924 6724
rect 14507 6684 14924 6712
rect 14507 6681 14519 6684
rect 14461 6675 14519 6681
rect 14918 6672 14924 6684
rect 14976 6672 14982 6724
rect 15378 6672 15384 6724
rect 15436 6712 15442 6724
rect 16298 6712 16304 6724
rect 15436 6684 16304 6712
rect 15436 6672 15442 6684
rect 16298 6672 16304 6684
rect 16356 6712 16362 6724
rect 16853 6715 16911 6721
rect 16853 6712 16865 6715
rect 16356 6684 16865 6712
rect 16356 6672 16362 6684
rect 16853 6681 16865 6684
rect 16899 6681 16911 6715
rect 19613 6715 19671 6721
rect 19613 6712 19625 6715
rect 16853 6675 16911 6681
rect 16960 6684 19625 6712
rect 16960 6656 16988 6684
rect 19613 6681 19625 6684
rect 19659 6681 19671 6715
rect 19613 6675 19671 6681
rect 12584 6616 12629 6644
rect 13096 6616 13768 6644
rect 12584 6604 12590 6616
rect 13814 6604 13820 6656
rect 13872 6644 13878 6656
rect 14093 6647 14151 6653
rect 14093 6644 14105 6647
rect 13872 6616 14105 6644
rect 13872 6604 13878 6616
rect 14093 6613 14105 6616
rect 14139 6613 14151 6647
rect 14093 6607 14151 6613
rect 14553 6647 14611 6653
rect 14553 6613 14565 6647
rect 14599 6644 14611 6647
rect 15010 6644 15016 6656
rect 14599 6616 15016 6644
rect 14599 6613 14611 6616
rect 14553 6607 14611 6613
rect 15010 6604 15016 6616
rect 15068 6604 15074 6656
rect 15289 6647 15347 6653
rect 15289 6613 15301 6647
rect 15335 6644 15347 6647
rect 15933 6647 15991 6653
rect 15933 6644 15945 6647
rect 15335 6616 15945 6644
rect 15335 6613 15347 6616
rect 15289 6607 15347 6613
rect 15933 6613 15945 6616
rect 15979 6613 15991 6647
rect 15933 6607 15991 6613
rect 16942 6604 16948 6656
rect 17000 6644 17006 6656
rect 18233 6647 18291 6653
rect 17000 6616 17045 6644
rect 17000 6604 17006 6616
rect 18233 6613 18245 6647
rect 18279 6644 18291 6647
rect 18598 6644 18604 6656
rect 18279 6616 18604 6644
rect 18279 6613 18291 6616
rect 18233 6607 18291 6613
rect 18598 6604 18604 6616
rect 18656 6604 18662 6656
rect 20165 6647 20223 6653
rect 20165 6613 20177 6647
rect 20211 6644 20223 6647
rect 20346 6644 20352 6656
rect 20211 6616 20352 6644
rect 20211 6613 20223 6616
rect 20165 6607 20223 6613
rect 20346 6604 20352 6616
rect 20404 6604 20410 6656
rect 20993 6647 21051 6653
rect 20993 6613 21005 6647
rect 21039 6644 21051 6647
rect 22554 6644 22560 6656
rect 21039 6616 22560 6644
rect 21039 6613 21051 6616
rect 20993 6607 21051 6613
rect 22554 6604 22560 6616
rect 22612 6604 22618 6656
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 9493 6443 9551 6449
rect 9493 6409 9505 6443
rect 9539 6440 9551 6443
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 9539 6412 10057 6440
rect 9539 6409 9551 6412
rect 9493 6403 9551 6409
rect 10045 6409 10057 6412
rect 10091 6409 10103 6443
rect 10502 6440 10508 6452
rect 10463 6412 10508 6440
rect 10045 6403 10103 6409
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 11146 6400 11152 6452
rect 11204 6440 11210 6452
rect 12069 6443 12127 6449
rect 12069 6440 12081 6443
rect 11204 6412 12081 6440
rect 11204 6400 11210 6412
rect 12069 6409 12081 6412
rect 12115 6440 12127 6443
rect 12434 6440 12440 6452
rect 12115 6412 12440 6440
rect 12115 6409 12127 6412
rect 12069 6403 12127 6409
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 12529 6443 12587 6449
rect 12529 6409 12541 6443
rect 12575 6440 12587 6443
rect 12618 6440 12624 6452
rect 12575 6412 12624 6440
rect 12575 6409 12587 6412
rect 12529 6403 12587 6409
rect 12618 6400 12624 6412
rect 12676 6400 12682 6452
rect 13170 6440 13176 6452
rect 13131 6412 13176 6440
rect 13170 6400 13176 6412
rect 13228 6400 13234 6452
rect 14553 6443 14611 6449
rect 14553 6409 14565 6443
rect 14599 6440 14611 6443
rect 16669 6443 16727 6449
rect 16669 6440 16681 6443
rect 14599 6412 16681 6440
rect 14599 6409 14611 6412
rect 14553 6403 14611 6409
rect 16669 6409 16681 6412
rect 16715 6409 16727 6443
rect 16669 6403 16727 6409
rect 17037 6443 17095 6449
rect 17037 6409 17049 6443
rect 17083 6440 17095 6443
rect 17494 6440 17500 6452
rect 17083 6412 17500 6440
rect 17083 6409 17095 6412
rect 17037 6403 17095 6409
rect 17494 6400 17500 6412
rect 17552 6400 17558 6452
rect 18141 6443 18199 6449
rect 18141 6409 18153 6443
rect 18187 6440 18199 6443
rect 18782 6440 18788 6452
rect 18187 6412 18788 6440
rect 18187 6409 18199 6412
rect 18141 6403 18199 6409
rect 18782 6400 18788 6412
rect 18840 6440 18846 6452
rect 18966 6440 18972 6452
rect 18840 6412 18972 6440
rect 18840 6400 18846 6412
rect 18966 6400 18972 6412
rect 19024 6440 19030 6452
rect 19242 6440 19248 6452
rect 19024 6412 19248 6440
rect 19024 6400 19030 6412
rect 19242 6400 19248 6412
rect 19300 6400 19306 6452
rect 12710 6332 12716 6384
rect 12768 6372 12774 6384
rect 12894 6372 12900 6384
rect 12768 6344 12900 6372
rect 12768 6332 12774 6344
rect 12894 6332 12900 6344
rect 12952 6372 12958 6384
rect 13538 6372 13544 6384
rect 12952 6344 13544 6372
rect 12952 6332 12958 6344
rect 13538 6332 13544 6344
rect 13596 6332 13602 6384
rect 14918 6332 14924 6384
rect 14976 6372 14982 6384
rect 18049 6375 18107 6381
rect 14976 6344 17172 6372
rect 14976 6332 14982 6344
rect 9122 6304 9128 6316
rect 9083 6276 9128 6304
rect 9122 6264 9128 6276
rect 9180 6264 9186 6316
rect 10134 6304 10140 6316
rect 10095 6276 10140 6304
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6304 11207 6307
rect 12158 6304 12164 6316
rect 11195 6276 12164 6304
rect 11195 6273 11207 6276
rect 11149 6267 11207 6273
rect 12158 6264 12164 6276
rect 12216 6264 12222 6316
rect 12986 6264 12992 6316
rect 13044 6304 13050 6316
rect 13044 6276 13400 6304
rect 13044 6264 13050 6276
rect 8941 6239 8999 6245
rect 8941 6205 8953 6239
rect 8987 6205 8999 6239
rect 8941 6199 8999 6205
rect 9033 6239 9091 6245
rect 9033 6205 9045 6239
rect 9079 6236 9091 6239
rect 9766 6236 9772 6248
rect 9079 6208 9772 6236
rect 9079 6205 9091 6208
rect 9033 6199 9091 6205
rect 8956 6168 8984 6199
rect 9766 6196 9772 6208
rect 9824 6196 9830 6248
rect 9953 6239 10011 6245
rect 9953 6205 9965 6239
rect 9999 6236 10011 6239
rect 10226 6236 10232 6248
rect 9999 6208 10232 6236
rect 9999 6205 10011 6208
rect 9953 6199 10011 6205
rect 10226 6196 10232 6208
rect 10284 6196 10290 6248
rect 10686 6196 10692 6248
rect 10744 6236 10750 6248
rect 11885 6239 11943 6245
rect 11885 6236 11897 6239
rect 10744 6208 11897 6236
rect 10744 6196 10750 6208
rect 11885 6205 11897 6208
rect 11931 6205 11943 6239
rect 11885 6199 11943 6205
rect 12894 6196 12900 6248
rect 12952 6236 12958 6248
rect 13372 6245 13400 6276
rect 13722 6264 13728 6316
rect 13780 6304 13786 6316
rect 14458 6304 14464 6316
rect 13780 6276 14464 6304
rect 13780 6264 13786 6276
rect 14458 6264 14464 6276
rect 14516 6264 14522 6316
rect 15473 6307 15531 6313
rect 15473 6273 15485 6307
rect 15519 6304 15531 6307
rect 15930 6304 15936 6316
rect 15519 6276 15936 6304
rect 15519 6273 15531 6276
rect 15473 6267 15531 6273
rect 15930 6264 15936 6276
rect 15988 6264 15994 6316
rect 16114 6264 16120 6316
rect 16172 6304 16178 6316
rect 17034 6304 17040 6316
rect 16172 6276 17040 6304
rect 16172 6264 16178 6276
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 17144 6304 17172 6344
rect 18049 6341 18061 6375
rect 18095 6372 18107 6375
rect 18230 6372 18236 6384
rect 18095 6344 18236 6372
rect 18095 6341 18107 6344
rect 18049 6335 18107 6341
rect 18230 6332 18236 6344
rect 18288 6372 18294 6384
rect 19518 6372 19524 6384
rect 18288 6344 19524 6372
rect 18288 6332 18294 6344
rect 19518 6332 19524 6344
rect 19576 6332 19582 6384
rect 19978 6372 19984 6384
rect 19939 6344 19984 6372
rect 19978 6332 19984 6344
rect 20036 6332 20042 6384
rect 20898 6332 20904 6384
rect 20956 6372 20962 6384
rect 20993 6375 21051 6381
rect 20993 6372 21005 6375
rect 20956 6344 21005 6372
rect 20956 6332 20962 6344
rect 20993 6341 21005 6344
rect 21039 6341 21051 6375
rect 20993 6335 21051 6341
rect 19702 6304 19708 6316
rect 17144 6276 18828 6304
rect 19663 6276 19708 6304
rect 13265 6239 13323 6245
rect 13265 6236 13277 6239
rect 12952 6208 13277 6236
rect 12952 6196 12958 6208
rect 13265 6205 13277 6208
rect 13311 6205 13323 6239
rect 13265 6199 13323 6205
rect 13357 6239 13415 6245
rect 13357 6205 13369 6239
rect 13403 6205 13415 6239
rect 14734 6236 14740 6248
rect 14695 6208 14740 6236
rect 13357 6199 13415 6205
rect 14734 6196 14740 6208
rect 14792 6196 14798 6248
rect 15286 6236 15292 6248
rect 15247 6208 15292 6236
rect 15286 6196 15292 6208
rect 15344 6196 15350 6248
rect 15381 6239 15439 6245
rect 15381 6205 15393 6239
rect 15427 6236 15439 6239
rect 16942 6236 16948 6248
rect 15427 6208 16948 6236
rect 15427 6205 15439 6208
rect 15381 6199 15439 6205
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 17129 6239 17187 6245
rect 17129 6205 17141 6239
rect 17175 6236 17187 6239
rect 17218 6236 17224 6248
rect 17175 6208 17224 6236
rect 17175 6205 17187 6208
rect 17129 6199 17187 6205
rect 17218 6196 17224 6208
rect 17276 6196 17282 6248
rect 17313 6239 17371 6245
rect 17313 6205 17325 6239
rect 17359 6236 17371 6239
rect 17586 6236 17592 6248
rect 17359 6208 17592 6236
rect 17359 6205 17371 6208
rect 17313 6199 17371 6205
rect 17586 6196 17592 6208
rect 17644 6196 17650 6248
rect 17770 6196 17776 6248
rect 17828 6236 17834 6248
rect 18800 6245 18828 6276
rect 19702 6264 19708 6276
rect 19760 6264 19766 6316
rect 18233 6239 18291 6245
rect 18233 6236 18245 6239
rect 17828 6208 18245 6236
rect 17828 6196 17834 6208
rect 18233 6205 18245 6208
rect 18279 6205 18291 6239
rect 18233 6199 18291 6205
rect 18785 6239 18843 6245
rect 18785 6205 18797 6239
rect 18831 6236 18843 6239
rect 19610 6236 19616 6248
rect 18831 6208 19616 6236
rect 18831 6205 18843 6208
rect 18785 6199 18843 6205
rect 19610 6196 19616 6208
rect 19668 6236 19674 6248
rect 19886 6236 19892 6248
rect 19668 6208 19892 6236
rect 19668 6196 19674 6208
rect 19886 6196 19892 6208
rect 19944 6196 19950 6248
rect 21082 6236 21088 6248
rect 21043 6208 21088 6236
rect 21082 6196 21088 6208
rect 21140 6196 21146 6248
rect 21174 6196 21180 6248
rect 21232 6236 21238 6248
rect 21542 6236 21548 6248
rect 21232 6208 21548 6236
rect 21232 6196 21238 6208
rect 21542 6196 21548 6208
rect 21600 6196 21606 6248
rect 9490 6168 9496 6180
rect 8956 6140 9496 6168
rect 9490 6128 9496 6140
rect 9548 6128 9554 6180
rect 11146 6128 11152 6180
rect 11204 6168 11210 6180
rect 12805 6171 12863 6177
rect 12805 6168 12817 6171
rect 11204 6140 12817 6168
rect 11204 6128 11210 6140
rect 12805 6137 12817 6140
rect 12851 6137 12863 6171
rect 12805 6131 12863 6137
rect 15841 6171 15899 6177
rect 15841 6137 15853 6171
rect 15887 6168 15899 6171
rect 16758 6168 16764 6180
rect 15887 6140 16764 6168
rect 15887 6137 15899 6140
rect 15841 6131 15899 6137
rect 16758 6128 16764 6140
rect 16816 6128 16822 6180
rect 17954 6168 17960 6180
rect 17052 6140 17960 6168
rect 8018 6060 8024 6112
rect 8076 6100 8082 6112
rect 11882 6100 11888 6112
rect 8076 6072 11888 6100
rect 8076 6060 8082 6072
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 13446 6060 13452 6112
rect 13504 6100 13510 6112
rect 14093 6103 14151 6109
rect 14093 6100 14105 6103
rect 13504 6072 14105 6100
rect 13504 6060 13510 6072
rect 14093 6069 14105 6072
rect 14139 6069 14151 6103
rect 14093 6063 14151 6069
rect 15010 6060 15016 6112
rect 15068 6100 15074 6112
rect 16209 6103 16267 6109
rect 16209 6100 16221 6103
rect 15068 6072 16221 6100
rect 15068 6060 15074 6072
rect 16209 6069 16221 6072
rect 16255 6100 16267 6103
rect 17052 6100 17080 6140
rect 17954 6128 17960 6140
rect 18012 6128 18018 6180
rect 18046 6128 18052 6180
rect 18104 6168 18110 6180
rect 19061 6171 19119 6177
rect 19061 6168 19073 6171
rect 18104 6140 19073 6168
rect 18104 6128 18110 6140
rect 19061 6137 19073 6140
rect 19107 6137 19119 6171
rect 19061 6131 19119 6137
rect 16255 6072 17080 6100
rect 16255 6069 16267 6072
rect 16209 6063 16267 6069
rect 17126 6060 17132 6112
rect 17184 6100 17190 6112
rect 17681 6103 17739 6109
rect 17681 6100 17693 6103
rect 17184 6072 17693 6100
rect 17184 6060 17190 6072
rect 17681 6069 17693 6072
rect 17727 6069 17739 6103
rect 17681 6063 17739 6069
rect 18138 6060 18144 6112
rect 18196 6100 18202 6112
rect 19334 6100 19340 6112
rect 18196 6072 19340 6100
rect 18196 6060 18202 6072
rect 19334 6060 19340 6072
rect 19392 6060 19398 6112
rect 19886 6060 19892 6112
rect 19944 6100 19950 6112
rect 20625 6103 20683 6109
rect 20625 6100 20637 6103
rect 19944 6072 20637 6100
rect 19944 6060 19950 6072
rect 20625 6069 20637 6072
rect 20671 6069 20683 6103
rect 20625 6063 20683 6069
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 3510 5856 3516 5908
rect 3568 5896 3574 5908
rect 8294 5896 8300 5908
rect 3568 5868 8300 5896
rect 3568 5856 3574 5868
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 9033 5899 9091 5905
rect 9033 5865 9045 5899
rect 9079 5896 9091 5899
rect 9214 5896 9220 5908
rect 9079 5868 9220 5896
rect 9079 5865 9091 5868
rect 9033 5859 9091 5865
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 10045 5899 10103 5905
rect 10045 5865 10057 5899
rect 10091 5896 10103 5899
rect 10134 5896 10140 5908
rect 10091 5868 10140 5896
rect 10091 5865 10103 5868
rect 10045 5859 10103 5865
rect 10134 5856 10140 5868
rect 10192 5856 10198 5908
rect 10410 5896 10416 5908
rect 10371 5868 10416 5896
rect 10410 5856 10416 5868
rect 10468 5856 10474 5908
rect 11882 5896 11888 5908
rect 11843 5868 11888 5896
rect 11882 5856 11888 5868
rect 11940 5856 11946 5908
rect 12894 5896 12900 5908
rect 12855 5868 12900 5896
rect 12894 5856 12900 5868
rect 12952 5856 12958 5908
rect 13814 5896 13820 5908
rect 13096 5868 13820 5896
rect 8478 5788 8484 5840
rect 8536 5828 8542 5840
rect 8536 5800 9628 5828
rect 8536 5788 8542 5800
rect 9490 5760 9496 5772
rect 9451 5732 9496 5760
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 9600 5760 9628 5800
rect 9950 5788 9956 5840
rect 10008 5828 10014 5840
rect 10428 5828 10456 5856
rect 10008 5800 10456 5828
rect 10008 5788 10014 5800
rect 11241 5763 11299 5769
rect 11241 5760 11253 5763
rect 9600 5732 11253 5760
rect 11241 5729 11253 5732
rect 11287 5729 11299 5763
rect 11241 5723 11299 5729
rect 12342 5720 12348 5772
rect 12400 5760 12406 5772
rect 12437 5763 12495 5769
rect 12437 5760 12449 5763
rect 12400 5732 12449 5760
rect 12400 5720 12406 5732
rect 12437 5729 12449 5732
rect 12483 5729 12495 5763
rect 12437 5723 12495 5729
rect 9674 5692 9680 5704
rect 9635 5664 9680 5692
rect 9674 5652 9680 5664
rect 9732 5652 9738 5704
rect 11057 5695 11115 5701
rect 11057 5661 11069 5695
rect 11103 5692 11115 5695
rect 11146 5692 11152 5704
rect 11103 5664 11152 5692
rect 11103 5661 11115 5664
rect 11057 5655 11115 5661
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 12253 5695 12311 5701
rect 12253 5661 12265 5695
rect 12299 5692 12311 5695
rect 12526 5692 12532 5704
rect 12299 5664 12532 5692
rect 12299 5661 12311 5664
rect 12253 5655 12311 5661
rect 12526 5652 12532 5664
rect 12584 5652 12590 5704
rect 8294 5584 8300 5636
rect 8352 5624 8358 5636
rect 12345 5627 12403 5633
rect 8352 5596 12020 5624
rect 8352 5584 8358 5596
rect 9582 5556 9588 5568
rect 9543 5528 9588 5556
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 10689 5559 10747 5565
rect 10689 5525 10701 5559
rect 10735 5556 10747 5559
rect 10962 5556 10968 5568
rect 10735 5528 10968 5556
rect 10735 5525 10747 5528
rect 10689 5519 10747 5525
rect 10962 5516 10968 5528
rect 11020 5516 11026 5568
rect 11146 5516 11152 5568
rect 11204 5556 11210 5568
rect 11992 5556 12020 5596
rect 12345 5593 12357 5627
rect 12391 5624 12403 5627
rect 13096 5624 13124 5868
rect 13814 5856 13820 5868
rect 13872 5856 13878 5908
rect 15194 5856 15200 5908
rect 15252 5896 15258 5908
rect 15930 5896 15936 5908
rect 15252 5868 15608 5896
rect 15891 5868 15936 5896
rect 15252 5856 15258 5868
rect 13722 5788 13728 5840
rect 13780 5828 13786 5840
rect 14921 5831 14979 5837
rect 14921 5828 14933 5831
rect 13780 5800 14933 5828
rect 13780 5788 13786 5800
rect 14921 5797 14933 5800
rect 14967 5797 14979 5831
rect 14921 5791 14979 5797
rect 15378 5788 15384 5840
rect 15436 5828 15442 5840
rect 15580 5828 15608 5868
rect 15930 5856 15936 5868
rect 15988 5856 15994 5908
rect 16942 5896 16948 5908
rect 16903 5868 16948 5896
rect 16942 5856 16948 5868
rect 17000 5856 17006 5908
rect 17034 5856 17040 5908
rect 17092 5896 17098 5908
rect 18138 5896 18144 5908
rect 17092 5868 18144 5896
rect 17092 5856 17098 5868
rect 18138 5856 18144 5868
rect 18196 5856 18202 5908
rect 17310 5828 17316 5840
rect 15436 5800 15516 5828
rect 15580 5800 17316 5828
rect 15436 5788 15442 5800
rect 13538 5760 13544 5772
rect 13499 5732 13544 5760
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 15488 5769 15516 5800
rect 17310 5788 17316 5800
rect 17368 5828 17374 5840
rect 17770 5828 17776 5840
rect 17368 5800 17776 5828
rect 17368 5788 17374 5800
rect 17770 5788 17776 5800
rect 17828 5788 17834 5840
rect 19058 5828 19064 5840
rect 18340 5800 19064 5828
rect 15473 5763 15531 5769
rect 15473 5729 15485 5763
rect 15519 5760 15531 5763
rect 15654 5760 15660 5772
rect 15519 5732 15660 5760
rect 15519 5729 15531 5732
rect 15473 5723 15531 5729
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 16022 5720 16028 5772
rect 16080 5760 16086 5772
rect 16206 5760 16212 5772
rect 16080 5732 16212 5760
rect 16080 5720 16086 5732
rect 16206 5720 16212 5732
rect 16264 5760 16270 5772
rect 16393 5763 16451 5769
rect 16393 5760 16405 5763
rect 16264 5732 16405 5760
rect 16264 5720 16270 5732
rect 16393 5729 16405 5732
rect 16439 5729 16451 5763
rect 16393 5723 16451 5729
rect 16577 5763 16635 5769
rect 16577 5729 16589 5763
rect 16623 5760 16635 5763
rect 17494 5760 17500 5772
rect 16623 5732 17500 5760
rect 16623 5729 16635 5732
rect 16577 5723 16635 5729
rect 17494 5720 17500 5732
rect 17552 5720 17558 5772
rect 17586 5720 17592 5772
rect 17644 5760 17650 5772
rect 18138 5760 18144 5772
rect 17644 5732 18144 5760
rect 17644 5720 17650 5732
rect 18138 5720 18144 5732
rect 18196 5720 18202 5772
rect 18340 5769 18368 5800
rect 19058 5788 19064 5800
rect 19116 5828 19122 5840
rect 19978 5828 19984 5840
rect 19116 5800 19984 5828
rect 19116 5788 19122 5800
rect 19978 5788 19984 5800
rect 20036 5788 20042 5840
rect 18325 5763 18383 5769
rect 18325 5729 18337 5763
rect 18371 5729 18383 5763
rect 18325 5723 18383 5729
rect 18414 5720 18420 5772
rect 18472 5760 18478 5772
rect 19705 5763 19763 5769
rect 18472 5732 18517 5760
rect 18472 5720 18478 5732
rect 19705 5729 19717 5763
rect 19751 5760 19763 5763
rect 19794 5760 19800 5772
rect 19751 5732 19800 5760
rect 19751 5729 19763 5732
rect 19705 5723 19763 5729
rect 19794 5720 19800 5732
rect 19852 5760 19858 5772
rect 21085 5763 21143 5769
rect 21085 5760 21097 5763
rect 19852 5732 21097 5760
rect 19852 5720 19858 5732
rect 21085 5729 21097 5732
rect 21131 5729 21143 5763
rect 21085 5723 21143 5729
rect 13170 5652 13176 5704
rect 13228 5692 13234 5704
rect 13357 5695 13415 5701
rect 13357 5692 13369 5695
rect 13228 5664 13369 5692
rect 13228 5652 13234 5664
rect 13357 5661 13369 5664
rect 13403 5692 13415 5695
rect 13814 5692 13820 5704
rect 13403 5664 13820 5692
rect 13403 5661 13415 5664
rect 13357 5655 13415 5661
rect 13814 5652 13820 5664
rect 13872 5652 13878 5704
rect 15194 5652 15200 5704
rect 15252 5692 15258 5704
rect 15289 5695 15347 5701
rect 15289 5692 15301 5695
rect 15252 5664 15301 5692
rect 15252 5652 15258 5664
rect 15289 5661 15301 5664
rect 15335 5661 15347 5695
rect 17402 5692 17408 5704
rect 17363 5664 17408 5692
rect 15289 5655 15347 5661
rect 17402 5652 17408 5664
rect 17460 5652 17466 5704
rect 18506 5692 18512 5704
rect 18419 5664 18512 5692
rect 18506 5652 18512 5664
rect 18564 5692 18570 5704
rect 18874 5692 18880 5704
rect 18564 5664 18880 5692
rect 18564 5652 18570 5664
rect 18874 5652 18880 5664
rect 18932 5652 18938 5704
rect 19886 5692 19892 5704
rect 19847 5664 19892 5692
rect 19886 5652 19892 5664
rect 19944 5652 19950 5704
rect 20898 5652 20904 5704
rect 20956 5692 20962 5704
rect 20993 5695 21051 5701
rect 20993 5692 21005 5695
rect 20956 5664 21005 5692
rect 20956 5652 20962 5664
rect 20993 5661 21005 5664
rect 21039 5692 21051 5695
rect 22278 5692 22284 5704
rect 21039 5664 22284 5692
rect 21039 5661 21051 5664
rect 20993 5655 21051 5661
rect 22278 5652 22284 5664
rect 22336 5652 22342 5704
rect 12391 5596 13124 5624
rect 14645 5627 14703 5633
rect 12391 5593 12403 5596
rect 12345 5587 12403 5593
rect 14645 5593 14657 5627
rect 14691 5624 14703 5627
rect 16301 5627 16359 5633
rect 16301 5624 16313 5627
rect 14691 5596 16313 5624
rect 14691 5593 14703 5596
rect 14645 5587 14703 5593
rect 16301 5593 16313 5596
rect 16347 5593 16359 5627
rect 16301 5587 16359 5593
rect 16482 5584 16488 5636
rect 16540 5624 16546 5636
rect 19797 5627 19855 5633
rect 19797 5624 19809 5627
rect 16540 5596 19809 5624
rect 16540 5584 16546 5596
rect 19797 5593 19809 5596
rect 19843 5593 19855 5627
rect 19797 5587 19855 5593
rect 13265 5559 13323 5565
rect 13265 5556 13277 5559
rect 11204 5528 11249 5556
rect 11992 5528 13277 5556
rect 11204 5516 11210 5528
rect 13265 5525 13277 5528
rect 13311 5556 13323 5559
rect 14185 5559 14243 5565
rect 14185 5556 14197 5559
rect 13311 5528 14197 5556
rect 13311 5525 13323 5528
rect 13265 5519 13323 5525
rect 14185 5525 14197 5528
rect 14231 5556 14243 5559
rect 15194 5556 15200 5568
rect 14231 5528 15200 5556
rect 14231 5525 14243 5528
rect 14185 5519 14243 5525
rect 15194 5516 15200 5528
rect 15252 5516 15258 5568
rect 15381 5559 15439 5565
rect 15381 5525 15393 5559
rect 15427 5556 15439 5559
rect 16114 5556 16120 5568
rect 15427 5528 16120 5556
rect 15427 5525 15439 5528
rect 15381 5519 15439 5525
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 16758 5516 16764 5568
rect 16816 5556 16822 5568
rect 17034 5556 17040 5568
rect 16816 5528 17040 5556
rect 16816 5516 16822 5528
rect 17034 5516 17040 5528
rect 17092 5516 17098 5568
rect 17313 5559 17371 5565
rect 17313 5525 17325 5559
rect 17359 5556 17371 5559
rect 17494 5556 17500 5568
rect 17359 5528 17500 5556
rect 17359 5525 17371 5528
rect 17313 5519 17371 5525
rect 17494 5516 17500 5528
rect 17552 5556 17558 5568
rect 17678 5556 17684 5568
rect 17552 5528 17684 5556
rect 17552 5516 17558 5528
rect 17678 5516 17684 5528
rect 17736 5516 17742 5568
rect 18874 5556 18880 5568
rect 18835 5528 18880 5556
rect 18874 5516 18880 5528
rect 18932 5516 18938 5568
rect 20254 5556 20260 5568
rect 20215 5528 20260 5556
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 20530 5556 20536 5568
rect 20491 5528 20536 5556
rect 20530 5516 20536 5528
rect 20588 5516 20594 5568
rect 20898 5556 20904 5568
rect 20859 5528 20904 5556
rect 20898 5516 20904 5528
rect 20956 5516 20962 5568
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 8570 5352 8576 5364
rect 8168 5324 8576 5352
rect 8168 5312 8174 5324
rect 8570 5312 8576 5324
rect 8628 5312 8634 5364
rect 8754 5312 8760 5364
rect 8812 5352 8818 5364
rect 9493 5355 9551 5361
rect 8812 5324 9444 5352
rect 8812 5312 8818 5324
rect 5074 5244 5080 5296
rect 5132 5284 5138 5296
rect 5132 5256 8892 5284
rect 5132 5244 5138 5256
rect 6822 5176 6828 5228
rect 6880 5216 6886 5228
rect 8754 5216 8760 5228
rect 6880 5188 8760 5216
rect 6880 5176 6886 5188
rect 8754 5176 8760 5188
rect 8812 5176 8818 5228
rect 8864 5216 8892 5256
rect 8938 5244 8944 5296
rect 8996 5284 9002 5296
rect 9306 5284 9312 5296
rect 8996 5256 9312 5284
rect 8996 5244 9002 5256
rect 9306 5244 9312 5256
rect 9364 5244 9370 5296
rect 9416 5284 9444 5324
rect 9493 5321 9505 5355
rect 9539 5352 9551 5355
rect 9582 5352 9588 5364
rect 9539 5324 9588 5352
rect 9539 5321 9551 5324
rect 9493 5315 9551 5321
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 9950 5352 9956 5364
rect 9911 5324 9956 5352
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 10597 5355 10655 5361
rect 10597 5321 10609 5355
rect 10643 5352 10655 5355
rect 10778 5352 10784 5364
rect 10643 5324 10784 5352
rect 10643 5321 10655 5324
rect 10597 5315 10655 5321
rect 10134 5284 10140 5296
rect 9416 5256 10140 5284
rect 10134 5244 10140 5256
rect 10192 5244 10198 5296
rect 9125 5219 9183 5225
rect 9125 5216 9137 5219
rect 8864 5188 9137 5216
rect 9125 5185 9137 5188
rect 9171 5216 9183 5219
rect 9861 5219 9919 5225
rect 9861 5216 9873 5219
rect 9171 5188 9873 5216
rect 9171 5185 9183 5188
rect 9125 5179 9183 5185
rect 9861 5185 9873 5188
rect 9907 5185 9919 5219
rect 9861 5179 9919 5185
rect 7834 5108 7840 5160
rect 7892 5148 7898 5160
rect 7892 5120 9674 5148
rect 7892 5108 7898 5120
rect 9646 5080 9674 5120
rect 10042 5108 10048 5160
rect 10100 5148 10106 5160
rect 10137 5151 10195 5157
rect 10137 5148 10149 5151
rect 10100 5120 10149 5148
rect 10100 5108 10106 5120
rect 10137 5117 10149 5120
rect 10183 5148 10195 5151
rect 10612 5148 10640 5315
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 11701 5355 11759 5361
rect 11701 5352 11713 5355
rect 11204 5324 11713 5352
rect 11204 5312 11210 5324
rect 11701 5321 11713 5324
rect 11747 5321 11759 5355
rect 13446 5352 13452 5364
rect 13407 5324 13452 5352
rect 11701 5315 11759 5321
rect 13446 5312 13452 5324
rect 13504 5312 13510 5364
rect 13906 5352 13912 5364
rect 13867 5324 13912 5352
rect 13906 5312 13912 5324
rect 13964 5312 13970 5364
rect 14918 5352 14924 5364
rect 14879 5324 14924 5352
rect 14918 5312 14924 5324
rect 14976 5312 14982 5364
rect 15194 5312 15200 5364
rect 15252 5352 15258 5364
rect 15378 5352 15384 5364
rect 15252 5324 15384 5352
rect 15252 5312 15258 5324
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 15838 5352 15844 5364
rect 15799 5324 15844 5352
rect 15838 5312 15844 5324
rect 15896 5312 15902 5364
rect 16301 5355 16359 5361
rect 16301 5321 16313 5355
rect 16347 5352 16359 5355
rect 16390 5352 16396 5364
rect 16347 5324 16396 5352
rect 16347 5321 16359 5324
rect 16301 5315 16359 5321
rect 16390 5312 16396 5324
rect 16448 5312 16454 5364
rect 16758 5312 16764 5364
rect 16816 5352 16822 5364
rect 17773 5355 17831 5361
rect 16816 5324 17724 5352
rect 16816 5312 16822 5324
rect 12069 5287 12127 5293
rect 12069 5253 12081 5287
rect 12115 5284 12127 5287
rect 17126 5284 17132 5296
rect 12115 5256 17132 5284
rect 12115 5253 12127 5256
rect 12069 5247 12127 5253
rect 17126 5244 17132 5256
rect 17184 5244 17190 5296
rect 17696 5284 17724 5324
rect 17773 5321 17785 5355
rect 17819 5352 17831 5355
rect 18325 5355 18383 5361
rect 18325 5352 18337 5355
rect 17819 5324 18337 5352
rect 17819 5321 17831 5324
rect 17773 5315 17831 5321
rect 18325 5321 18337 5324
rect 18371 5321 18383 5355
rect 18325 5315 18383 5321
rect 18693 5355 18751 5361
rect 18693 5321 18705 5355
rect 18739 5352 18751 5355
rect 18874 5352 18880 5364
rect 18739 5324 18880 5352
rect 18739 5321 18751 5324
rect 18693 5315 18751 5321
rect 18874 5312 18880 5324
rect 18932 5312 18938 5364
rect 19260 5324 20208 5352
rect 19260 5284 19288 5324
rect 17696 5256 19288 5284
rect 13538 5216 13544 5228
rect 13499 5188 13544 5216
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 14829 5219 14887 5225
rect 14829 5185 14841 5219
rect 14875 5216 14887 5219
rect 15010 5216 15016 5228
rect 14875 5188 15016 5216
rect 14875 5185 14887 5188
rect 14829 5179 14887 5185
rect 15010 5176 15016 5188
rect 15068 5176 15074 5228
rect 15933 5219 15991 5225
rect 15933 5185 15945 5219
rect 15979 5185 15991 5219
rect 15933 5179 15991 5185
rect 16669 5219 16727 5225
rect 16669 5185 16681 5219
rect 16715 5216 16727 5219
rect 17402 5216 17408 5228
rect 16715 5188 17408 5216
rect 16715 5185 16727 5188
rect 16669 5179 16727 5185
rect 12158 5148 12164 5160
rect 10183 5120 10640 5148
rect 12119 5120 12164 5148
rect 10183 5117 10195 5120
rect 10137 5111 10195 5117
rect 12158 5108 12164 5120
rect 12216 5108 12222 5160
rect 12345 5151 12403 5157
rect 12345 5117 12357 5151
rect 12391 5148 12403 5151
rect 12802 5148 12808 5160
rect 12391 5120 12808 5148
rect 12391 5117 12403 5120
rect 12345 5111 12403 5117
rect 12802 5108 12808 5120
rect 12860 5108 12866 5160
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5148 12955 5151
rect 12986 5148 12992 5160
rect 12943 5120 12992 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 12986 5108 12992 5120
rect 13044 5108 13050 5160
rect 13354 5148 13360 5160
rect 13315 5120 13360 5148
rect 13354 5108 13360 5120
rect 13412 5108 13418 5160
rect 14642 5148 14648 5160
rect 14603 5120 14648 5148
rect 14642 5108 14648 5120
rect 14700 5108 14706 5160
rect 15749 5151 15807 5157
rect 15749 5117 15761 5151
rect 15795 5117 15807 5151
rect 15948 5148 15976 5179
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 17678 5216 17684 5228
rect 17639 5188 17684 5216
rect 17678 5176 17684 5188
rect 17736 5176 17742 5228
rect 19705 5219 19763 5225
rect 19705 5185 19717 5219
rect 19751 5216 19763 5219
rect 20180 5216 20208 5324
rect 20530 5312 20536 5364
rect 20588 5352 20594 5364
rect 20717 5355 20775 5361
rect 20717 5352 20729 5355
rect 20588 5324 20729 5352
rect 20588 5312 20594 5324
rect 20717 5321 20729 5324
rect 20763 5321 20775 5355
rect 20717 5315 20775 5321
rect 20254 5244 20260 5296
rect 20312 5284 20318 5296
rect 20809 5287 20867 5293
rect 20809 5284 20821 5287
rect 20312 5256 20821 5284
rect 20312 5244 20318 5256
rect 20809 5253 20821 5256
rect 20855 5253 20867 5287
rect 20809 5247 20867 5253
rect 21174 5216 21180 5228
rect 19751 5188 20116 5216
rect 20180 5188 21180 5216
rect 19751 5185 19763 5188
rect 19705 5179 19763 5185
rect 17218 5148 17224 5160
rect 15948 5120 17224 5148
rect 15749 5111 15807 5117
rect 11146 5080 11152 5092
rect 9646 5052 11152 5080
rect 11146 5040 11152 5052
rect 11204 5080 11210 5092
rect 14366 5080 14372 5092
rect 11204 5052 14372 5080
rect 11204 5040 11210 5052
rect 14366 5040 14372 5052
rect 14424 5040 14430 5092
rect 15764 5080 15792 5111
rect 17218 5108 17224 5120
rect 17276 5108 17282 5160
rect 17862 5148 17868 5160
rect 17823 5120 17868 5148
rect 17862 5108 17868 5120
rect 17920 5108 17926 5160
rect 18785 5151 18843 5157
rect 18785 5117 18797 5151
rect 18831 5117 18843 5151
rect 18785 5111 18843 5117
rect 16758 5080 16764 5092
rect 15764 5052 16764 5080
rect 16758 5040 16764 5052
rect 16816 5040 16822 5092
rect 16853 5083 16911 5089
rect 16853 5049 16865 5083
rect 16899 5080 16911 5083
rect 18046 5080 18052 5092
rect 16899 5052 18052 5080
rect 16899 5049 16911 5052
rect 16853 5043 16911 5049
rect 18046 5040 18052 5052
rect 18104 5040 18110 5092
rect 18800 5080 18828 5111
rect 18874 5108 18880 5160
rect 18932 5148 18938 5160
rect 18969 5151 19027 5157
rect 18969 5148 18981 5151
rect 18932 5120 18981 5148
rect 18932 5108 18938 5120
rect 18969 5117 18981 5120
rect 19015 5148 19027 5151
rect 19794 5148 19800 5160
rect 19015 5120 19656 5148
rect 19755 5120 19800 5148
rect 19015 5117 19027 5120
rect 18969 5111 19027 5117
rect 19337 5083 19395 5089
rect 19337 5080 19349 5083
rect 18800 5052 19349 5080
rect 19337 5049 19349 5052
rect 19383 5049 19395 5083
rect 19628 5080 19656 5120
rect 19794 5108 19800 5120
rect 19852 5108 19858 5160
rect 19978 5148 19984 5160
rect 19939 5120 19984 5148
rect 19978 5108 19984 5120
rect 20036 5108 20042 5160
rect 20088 5148 20116 5188
rect 21174 5176 21180 5188
rect 21232 5176 21238 5228
rect 20438 5148 20444 5160
rect 20088 5120 20444 5148
rect 20438 5108 20444 5120
rect 20496 5108 20502 5160
rect 20990 5148 20996 5160
rect 20951 5120 20996 5148
rect 20990 5108 20996 5120
rect 21048 5108 21054 5160
rect 21634 5080 21640 5092
rect 19628 5052 21640 5080
rect 19337 5043 19395 5049
rect 21634 5040 21640 5052
rect 21692 5040 21698 5092
rect 2038 4972 2044 5024
rect 2096 5012 2102 5024
rect 5074 5012 5080 5024
rect 2096 4984 5080 5012
rect 2096 4972 2102 4984
rect 5074 4972 5080 4984
rect 5132 4972 5138 5024
rect 8478 5012 8484 5024
rect 8439 4984 8484 5012
rect 8478 4972 8484 4984
rect 8536 5012 8542 5024
rect 8938 5012 8944 5024
rect 8536 4984 8944 5012
rect 8536 4972 8542 4984
rect 8938 4972 8944 4984
rect 8996 4972 9002 5024
rect 13814 4972 13820 5024
rect 13872 5012 13878 5024
rect 14185 5015 14243 5021
rect 14185 5012 14197 5015
rect 13872 4984 14197 5012
rect 13872 4972 13878 4984
rect 14185 4981 14197 4984
rect 14231 5012 14243 5015
rect 14458 5012 14464 5024
rect 14231 4984 14464 5012
rect 14231 4981 14243 4984
rect 14185 4975 14243 4981
rect 14458 4972 14464 4984
rect 14516 4972 14522 5024
rect 15194 4972 15200 5024
rect 15252 5012 15258 5024
rect 15289 5015 15347 5021
rect 15289 5012 15301 5015
rect 15252 4984 15301 5012
rect 15252 4972 15258 4984
rect 15289 4981 15301 4984
rect 15335 4981 15347 5015
rect 15289 4975 15347 4981
rect 16114 4972 16120 5024
rect 16172 5012 16178 5024
rect 17126 5012 17132 5024
rect 16172 4984 17132 5012
rect 16172 4972 16178 4984
rect 17126 4972 17132 4984
rect 17184 4972 17190 5024
rect 17310 5012 17316 5024
rect 17271 4984 17316 5012
rect 17310 4972 17316 4984
rect 17368 4972 17374 5024
rect 20346 5012 20352 5024
rect 20307 4984 20352 5012
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 8481 4811 8539 4817
rect 8481 4808 8493 4811
rect 8260 4780 8493 4808
rect 8260 4768 8266 4780
rect 8481 4777 8493 4780
rect 8527 4777 8539 4811
rect 8481 4771 8539 4777
rect 1394 4700 1400 4752
rect 1452 4740 1458 4752
rect 1452 4712 2774 4740
rect 1452 4700 1458 4712
rect 2746 4536 2774 4712
rect 8496 4672 8524 4771
rect 9122 4768 9128 4820
rect 9180 4808 9186 4820
rect 9493 4811 9551 4817
rect 9493 4808 9505 4811
rect 9180 4780 9505 4808
rect 9180 4768 9186 4780
rect 9493 4777 9505 4780
rect 9539 4777 9551 4811
rect 9493 4771 9551 4777
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 10597 4811 10655 4817
rect 10597 4808 10609 4811
rect 9824 4780 10609 4808
rect 9824 4768 9830 4780
rect 10597 4777 10609 4780
rect 10643 4777 10655 4811
rect 10597 4771 10655 4777
rect 13538 4768 13544 4820
rect 13596 4808 13602 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 13596 4780 14105 4808
rect 13596 4768 13602 4780
rect 14093 4777 14105 4780
rect 14139 4777 14151 4811
rect 14093 4771 14151 4777
rect 15286 4768 15292 4820
rect 15344 4808 15350 4820
rect 16117 4811 16175 4817
rect 16117 4808 16129 4811
rect 15344 4780 16129 4808
rect 15344 4768 15350 4780
rect 16117 4777 16129 4780
rect 16163 4777 16175 4811
rect 16117 4771 16175 4777
rect 17678 4768 17684 4820
rect 17736 4808 17742 4820
rect 17865 4811 17923 4817
rect 17865 4808 17877 4811
rect 17736 4780 17877 4808
rect 17736 4768 17742 4780
rect 17865 4777 17877 4780
rect 17911 4777 17923 4811
rect 17865 4771 17923 4777
rect 19610 4768 19616 4820
rect 19668 4808 19674 4820
rect 19705 4811 19763 4817
rect 19705 4808 19717 4811
rect 19668 4780 19717 4808
rect 19668 4768 19674 4780
rect 19705 4777 19717 4780
rect 19751 4777 19763 4811
rect 20162 4808 20168 4820
rect 20123 4780 20168 4808
rect 19705 4771 19763 4777
rect 20162 4768 20168 4780
rect 20220 4768 20226 4820
rect 21266 4808 21272 4820
rect 21227 4780 21272 4808
rect 21266 4768 21272 4780
rect 21324 4768 21330 4820
rect 13170 4700 13176 4752
rect 13228 4740 13234 4752
rect 13633 4743 13691 4749
rect 13633 4740 13645 4743
rect 13228 4712 13645 4740
rect 13228 4700 13234 4712
rect 13633 4709 13645 4712
rect 13679 4709 13691 4743
rect 13633 4703 13691 4709
rect 17954 4700 17960 4752
rect 18012 4740 18018 4752
rect 21082 4740 21088 4752
rect 18012 4712 21088 4740
rect 18012 4700 18018 4712
rect 21082 4700 21088 4712
rect 21140 4700 21146 4752
rect 10042 4672 10048 4684
rect 8496 4644 9076 4672
rect 10003 4644 10048 4672
rect 7374 4564 7380 4616
rect 7432 4604 7438 4616
rect 8846 4604 8852 4616
rect 7432 4576 8852 4604
rect 7432 4564 7438 4576
rect 8846 4564 8852 4576
rect 8904 4604 8910 4616
rect 8941 4607 8999 4613
rect 8941 4604 8953 4607
rect 8904 4576 8953 4604
rect 8904 4564 8910 4576
rect 8941 4573 8953 4576
rect 8987 4573 8999 4607
rect 9048 4604 9076 4644
rect 10042 4632 10048 4644
rect 10100 4672 10106 4684
rect 10318 4672 10324 4684
rect 10100 4644 10324 4672
rect 10100 4632 10106 4644
rect 10318 4632 10324 4644
rect 10376 4672 10382 4684
rect 11149 4675 11207 4681
rect 11149 4672 11161 4675
rect 10376 4644 11161 4672
rect 10376 4632 10382 4644
rect 11149 4641 11161 4644
rect 11195 4641 11207 4675
rect 12250 4672 12256 4684
rect 12211 4644 12256 4672
rect 11149 4635 11207 4641
rect 12250 4632 12256 4644
rect 12308 4632 12314 4684
rect 13262 4672 13268 4684
rect 13223 4644 13268 4672
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 14734 4672 14740 4684
rect 14695 4644 14740 4672
rect 14734 4632 14740 4644
rect 14792 4632 14798 4684
rect 14918 4632 14924 4684
rect 14976 4672 14982 4684
rect 15102 4672 15108 4684
rect 14976 4644 15108 4672
rect 14976 4632 14982 4644
rect 15102 4632 15108 4644
rect 15160 4632 15166 4684
rect 15654 4672 15660 4684
rect 15615 4644 15660 4672
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 15838 4632 15844 4684
rect 15896 4672 15902 4684
rect 16485 4675 16543 4681
rect 16485 4672 16497 4675
rect 15896 4644 16497 4672
rect 15896 4632 15902 4644
rect 16485 4641 16497 4644
rect 16531 4641 16543 4675
rect 16485 4635 16543 4641
rect 18509 4675 18567 4681
rect 18509 4641 18521 4675
rect 18555 4672 18567 4675
rect 18874 4672 18880 4684
rect 18555 4644 18880 4672
rect 18555 4641 18567 4644
rect 18509 4635 18567 4641
rect 18874 4632 18880 4644
rect 18932 4632 18938 4684
rect 20254 4632 20260 4684
rect 20312 4672 20318 4684
rect 20441 4675 20499 4681
rect 20441 4672 20453 4675
rect 20312 4644 20453 4672
rect 20312 4632 20318 4644
rect 20441 4641 20453 4644
rect 20487 4641 20499 4675
rect 20441 4635 20499 4641
rect 20898 4632 20904 4684
rect 20956 4672 20962 4684
rect 20993 4675 21051 4681
rect 20993 4672 21005 4675
rect 20956 4644 21005 4672
rect 20956 4632 20962 4644
rect 20993 4641 21005 4644
rect 21039 4641 21051 4675
rect 20993 4635 21051 4641
rect 9953 4607 10011 4613
rect 9953 4604 9965 4607
rect 9048 4576 9965 4604
rect 8941 4567 8999 4573
rect 9953 4573 9965 4576
rect 9999 4573 10011 4607
rect 12986 4604 12992 4616
rect 12947 4576 12992 4604
rect 9953 4567 10011 4573
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 17034 4564 17040 4616
rect 17092 4604 17098 4616
rect 17129 4607 17187 4613
rect 17129 4604 17141 4607
rect 17092 4576 17141 4604
rect 17092 4564 17098 4576
rect 17129 4573 17141 4576
rect 17175 4573 17187 4607
rect 17129 4567 17187 4573
rect 17954 4564 17960 4616
rect 18012 4604 18018 4616
rect 18325 4607 18383 4613
rect 18325 4604 18337 4607
rect 18012 4576 18337 4604
rect 18012 4564 18018 4576
rect 18325 4573 18337 4576
rect 18371 4573 18383 4607
rect 18325 4567 18383 4573
rect 9674 4536 9680 4548
rect 2746 4508 9680 4536
rect 9674 4496 9680 4508
rect 9732 4496 9738 4548
rect 9861 4539 9919 4545
rect 9861 4505 9873 4539
rect 9907 4536 9919 4539
rect 10042 4536 10048 4548
rect 9907 4508 10048 4536
rect 9907 4505 9919 4508
rect 9861 4499 9919 4505
rect 10042 4496 10048 4508
rect 10100 4496 10106 4548
rect 10965 4539 11023 4545
rect 10965 4505 10977 4539
rect 11011 4536 11023 4539
rect 11146 4536 11152 4548
rect 11011 4508 11152 4536
rect 11011 4505 11023 4508
rect 10965 4499 11023 4505
rect 11146 4496 11152 4508
rect 11204 4496 11210 4548
rect 11977 4539 12035 4545
rect 11977 4505 11989 4539
rect 12023 4536 12035 4539
rect 13081 4539 13139 4545
rect 12023 4508 12664 4536
rect 12023 4505 12035 4508
rect 11977 4499 12035 4505
rect 9122 4468 9128 4480
rect 9083 4440 9128 4468
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 9692 4468 9720 4496
rect 10686 4468 10692 4480
rect 9692 4440 10692 4468
rect 10686 4428 10692 4440
rect 10744 4468 10750 4480
rect 11057 4471 11115 4477
rect 11057 4468 11069 4471
rect 10744 4440 11069 4468
rect 10744 4428 10750 4440
rect 11057 4437 11069 4440
rect 11103 4437 11115 4471
rect 11057 4431 11115 4437
rect 11609 4471 11667 4477
rect 11609 4437 11621 4471
rect 11655 4468 11667 4471
rect 11882 4468 11888 4480
rect 11655 4440 11888 4468
rect 11655 4437 11667 4440
rect 11609 4431 11667 4437
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 12069 4471 12127 4477
rect 12069 4437 12081 4471
rect 12115 4468 12127 4471
rect 12526 4468 12532 4480
rect 12115 4440 12532 4468
rect 12115 4437 12127 4440
rect 12069 4431 12127 4437
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 12636 4477 12664 4508
rect 13081 4505 13093 4539
rect 13127 4536 13139 4539
rect 13127 4508 15148 4536
rect 13127 4505 13139 4508
rect 13081 4499 13139 4505
rect 12621 4471 12679 4477
rect 12621 4437 12633 4471
rect 12667 4437 12679 4471
rect 12621 4431 12679 4437
rect 14182 4428 14188 4480
rect 14240 4468 14246 4480
rect 14461 4471 14519 4477
rect 14461 4468 14473 4471
rect 14240 4440 14473 4468
rect 14240 4428 14246 4440
rect 14461 4437 14473 4440
rect 14507 4437 14519 4471
rect 14461 4431 14519 4437
rect 14550 4428 14556 4480
rect 14608 4468 14614 4480
rect 15120 4477 15148 4508
rect 15378 4496 15384 4548
rect 15436 4536 15442 4548
rect 15473 4539 15531 4545
rect 15473 4536 15485 4539
rect 15436 4508 15485 4536
rect 15436 4496 15442 4508
rect 15473 4505 15485 4508
rect 15519 4536 15531 4539
rect 16022 4536 16028 4548
rect 15519 4508 16028 4536
rect 15519 4505 15531 4508
rect 15473 4499 15531 4505
rect 16022 4496 16028 4508
rect 16080 4496 16086 4548
rect 17405 4539 17463 4545
rect 17405 4505 17417 4539
rect 17451 4536 17463 4539
rect 17494 4536 17500 4548
rect 17451 4508 17500 4536
rect 17451 4505 17463 4508
rect 17405 4499 17463 4505
rect 17494 4496 17500 4508
rect 17552 4496 17558 4548
rect 18233 4539 18291 4545
rect 18233 4505 18245 4539
rect 18279 4536 18291 4539
rect 19245 4539 19303 4545
rect 19245 4536 19257 4539
rect 18279 4508 19257 4536
rect 18279 4505 18291 4508
rect 18233 4499 18291 4505
rect 19245 4505 19257 4508
rect 19291 4505 19303 4539
rect 19245 4499 19303 4505
rect 15105 4471 15163 4477
rect 14608 4440 14653 4468
rect 14608 4428 14614 4440
rect 15105 4437 15117 4471
rect 15151 4437 15163 4471
rect 15105 4431 15163 4437
rect 15565 4471 15623 4477
rect 15565 4437 15577 4471
rect 15611 4468 15623 4471
rect 15746 4468 15752 4480
rect 15611 4440 15752 4468
rect 15611 4437 15623 4440
rect 15565 4431 15623 4437
rect 15746 4428 15752 4440
rect 15804 4468 15810 4480
rect 20530 4468 20536 4480
rect 15804 4440 20536 4468
rect 15804 4428 15810 4440
rect 20530 4428 20536 4440
rect 20588 4428 20594 4480
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 8846 4264 8852 4276
rect 8807 4236 8852 4264
rect 8846 4224 8852 4236
rect 8904 4224 8910 4276
rect 9674 4264 9680 4276
rect 9635 4236 9680 4264
rect 9674 4224 9680 4236
rect 9732 4224 9738 4276
rect 10318 4264 10324 4276
rect 10279 4236 10324 4264
rect 10318 4224 10324 4236
rect 10376 4264 10382 4276
rect 11057 4267 11115 4273
rect 11057 4264 11069 4267
rect 10376 4236 11069 4264
rect 10376 4224 10382 4236
rect 11057 4233 11069 4236
rect 11103 4233 11115 4267
rect 11885 4267 11943 4273
rect 11885 4264 11897 4267
rect 11057 4227 11115 4233
rect 11164 4236 11897 4264
rect 8864 4196 8892 4224
rect 10689 4199 10747 4205
rect 10689 4196 10701 4199
rect 8864 4168 10701 4196
rect 10689 4165 10701 4168
rect 10735 4196 10747 4199
rect 11164 4196 11192 4236
rect 11885 4233 11897 4236
rect 11931 4233 11943 4267
rect 11885 4227 11943 4233
rect 12158 4224 12164 4276
rect 12216 4264 12222 4276
rect 12253 4267 12311 4273
rect 12253 4264 12265 4267
rect 12216 4236 12265 4264
rect 12216 4224 12222 4236
rect 12253 4233 12265 4236
rect 12299 4233 12311 4267
rect 12253 4227 12311 4233
rect 12526 4224 12532 4276
rect 12584 4264 12590 4276
rect 12989 4267 13047 4273
rect 12989 4264 13001 4267
rect 12584 4236 13001 4264
rect 12584 4224 12590 4236
rect 12989 4233 13001 4236
rect 13035 4233 13047 4267
rect 12989 4227 13047 4233
rect 13357 4267 13415 4273
rect 13357 4233 13369 4267
rect 13403 4264 13415 4267
rect 13722 4264 13728 4276
rect 13403 4236 13728 4264
rect 13403 4233 13415 4236
rect 13357 4227 13415 4233
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 14182 4264 14188 4276
rect 14143 4236 14188 4264
rect 14182 4224 14188 4236
rect 14240 4224 14246 4276
rect 15749 4267 15807 4273
rect 15749 4233 15761 4267
rect 15795 4264 15807 4267
rect 16022 4264 16028 4276
rect 15795 4236 16028 4264
rect 15795 4233 15807 4236
rect 15749 4227 15807 4233
rect 16022 4224 16028 4236
rect 16080 4224 16086 4276
rect 16761 4267 16819 4273
rect 16761 4233 16773 4267
rect 16807 4264 16819 4267
rect 17770 4264 17776 4276
rect 16807 4236 17776 4264
rect 16807 4233 16819 4236
rect 16761 4227 16819 4233
rect 17770 4224 17776 4236
rect 17828 4224 17834 4276
rect 11793 4199 11851 4205
rect 11793 4196 11805 4199
rect 10735 4168 11192 4196
rect 11532 4168 11805 4196
rect 10735 4165 10747 4168
rect 10689 4159 10747 4165
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 5902 4128 5908 4140
rect 3200 4100 5908 4128
rect 3200 4088 3206 4100
rect 5902 4088 5908 4100
rect 5960 4088 5966 4140
rect 10686 4020 10692 4072
rect 10744 4060 10750 4072
rect 11532 4060 11560 4168
rect 11793 4165 11805 4168
rect 11839 4165 11851 4199
rect 12621 4199 12679 4205
rect 12621 4196 12633 4199
rect 11793 4159 11851 4165
rect 12452 4168 12633 4196
rect 12452 4140 12480 4168
rect 12621 4165 12633 4168
rect 12667 4165 12679 4199
rect 12621 4159 12679 4165
rect 15105 4199 15163 4205
rect 15105 4165 15117 4199
rect 15151 4196 15163 4199
rect 16482 4196 16488 4208
rect 15151 4168 16488 4196
rect 15151 4165 15163 4168
rect 15105 4159 15163 4165
rect 16482 4156 16488 4168
rect 16540 4156 16546 4208
rect 17402 4156 17408 4208
rect 17460 4196 17466 4208
rect 19610 4196 19616 4208
rect 17460 4168 19616 4196
rect 17460 4156 17466 4168
rect 19610 4156 19616 4168
rect 19668 4156 19674 4208
rect 12434 4088 12440 4140
rect 12492 4088 12498 4140
rect 12710 4128 12716 4140
rect 12544 4100 12716 4128
rect 10744 4032 11560 4060
rect 11701 4063 11759 4069
rect 10744 4020 10750 4032
rect 11701 4029 11713 4063
rect 11747 4029 11759 4063
rect 12544 4060 12572 4100
rect 12710 4088 12716 4100
rect 12768 4088 12774 4140
rect 13262 4088 13268 4140
rect 13320 4128 13326 4140
rect 13320 4100 13584 4128
rect 13320 4088 13326 4100
rect 13446 4060 13452 4072
rect 11701 4023 11759 4029
rect 11900 4032 12572 4060
rect 13407 4032 13452 4060
rect 11716 3992 11744 4023
rect 11900 3992 11928 4032
rect 13446 4020 13452 4032
rect 13504 4020 13510 4072
rect 13556 4069 13584 4100
rect 14274 4088 14280 4140
rect 14332 4128 14338 4140
rect 17310 4128 17316 4140
rect 14332 4100 15700 4128
rect 17271 4100 17316 4128
rect 14332 4088 14338 4100
rect 13541 4063 13599 4069
rect 13541 4029 13553 4063
rect 13587 4029 13599 4063
rect 13541 4023 13599 4029
rect 14642 4020 14648 4072
rect 14700 4060 14706 4072
rect 15102 4060 15108 4072
rect 14700 4032 15108 4060
rect 14700 4020 14706 4032
rect 15102 4020 15108 4032
rect 15160 4060 15166 4072
rect 15672 4069 15700 4100
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 18693 4131 18751 4137
rect 18693 4097 18705 4131
rect 18739 4128 18751 4131
rect 20346 4128 20352 4140
rect 18739 4100 20352 4128
rect 18739 4097 18751 4100
rect 18693 4091 18751 4097
rect 20346 4088 20352 4100
rect 20404 4088 20410 4140
rect 20530 4128 20536 4140
rect 20491 4100 20536 4128
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 21174 4128 21180 4140
rect 21135 4100 21180 4128
rect 21174 4088 21180 4100
rect 21232 4088 21238 4140
rect 15473 4063 15531 4069
rect 15473 4060 15485 4063
rect 15160 4032 15485 4060
rect 15160 4020 15166 4032
rect 15473 4029 15485 4032
rect 15519 4029 15531 4063
rect 15473 4023 15531 4029
rect 15657 4063 15715 4069
rect 15657 4029 15669 4063
rect 15703 4060 15715 4063
rect 16298 4060 16304 4072
rect 15703 4032 16304 4060
rect 15703 4029 15715 4032
rect 15657 4023 15715 4029
rect 16298 4020 16304 4032
rect 16356 4020 16362 4072
rect 16942 4020 16948 4072
rect 17000 4060 17006 4072
rect 17497 4063 17555 4069
rect 17497 4060 17509 4063
rect 17000 4032 17509 4060
rect 17000 4020 17006 4032
rect 17497 4029 17509 4032
rect 17543 4029 17555 4063
rect 17497 4023 17555 4029
rect 18509 4063 18567 4069
rect 18509 4029 18521 4063
rect 18555 4060 18567 4063
rect 19058 4060 19064 4072
rect 18555 4032 19064 4060
rect 18555 4029 18567 4032
rect 18509 4023 18567 4029
rect 19058 4020 19064 4032
rect 19116 4020 19122 4072
rect 19150 4020 19156 4072
rect 19208 4060 19214 4072
rect 19705 4063 19763 4069
rect 19705 4060 19717 4063
rect 19208 4032 19717 4060
rect 19208 4020 19214 4032
rect 19705 4029 19717 4032
rect 19751 4029 19763 4063
rect 19705 4023 19763 4029
rect 19978 4020 19984 4072
rect 20036 4060 20042 4072
rect 20073 4063 20131 4069
rect 20073 4060 20085 4063
rect 20036 4032 20085 4060
rect 20036 4020 20042 4032
rect 20073 4029 20085 4032
rect 20119 4060 20131 4063
rect 20119 4032 20392 4060
rect 20119 4029 20131 4032
rect 20073 4023 20131 4029
rect 20364 4004 20392 4032
rect 14461 3995 14519 4001
rect 14461 3992 14473 3995
rect 11716 3964 11928 3992
rect 12728 3964 14473 3992
rect 934 3884 940 3936
rect 992 3924 998 3936
rect 8662 3924 8668 3936
rect 992 3896 8668 3924
rect 992 3884 998 3896
rect 8662 3884 8668 3896
rect 8720 3884 8726 3936
rect 10042 3924 10048 3936
rect 10003 3896 10048 3924
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 11698 3884 11704 3936
rect 11756 3924 11762 3936
rect 12728 3924 12756 3964
rect 14461 3961 14473 3964
rect 14507 3992 14519 3995
rect 14550 3992 14556 4004
rect 14507 3964 14556 3992
rect 14507 3961 14519 3964
rect 14461 3955 14519 3961
rect 14550 3952 14556 3964
rect 14608 3952 14614 4004
rect 14660 3964 16252 3992
rect 11756 3896 12756 3924
rect 11756 3884 11762 3896
rect 12802 3884 12808 3936
rect 12860 3924 12866 3936
rect 13630 3924 13636 3936
rect 12860 3896 13636 3924
rect 12860 3884 12866 3896
rect 13630 3884 13636 3896
rect 13688 3924 13694 3936
rect 14660 3924 14688 3964
rect 16114 3924 16120 3936
rect 13688 3896 14688 3924
rect 16075 3896 16120 3924
rect 13688 3884 13694 3896
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 16224 3924 16252 3964
rect 17862 3952 17868 4004
rect 17920 3992 17926 4004
rect 19794 3992 19800 4004
rect 17920 3964 19800 3992
rect 17920 3952 17926 3964
rect 19794 3952 19800 3964
rect 19852 3952 19858 4004
rect 20346 3952 20352 4004
rect 20404 3952 20410 4004
rect 18230 3924 18236 3936
rect 16224 3896 18236 3924
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 18782 3884 18788 3936
rect 18840 3924 18846 3936
rect 18969 3927 19027 3933
rect 18969 3924 18981 3927
rect 18840 3896 18981 3924
rect 18840 3884 18846 3896
rect 18969 3893 18981 3896
rect 19015 3893 19027 3927
rect 18969 3887 19027 3893
rect 19429 3927 19487 3933
rect 19429 3893 19441 3927
rect 19475 3924 19487 3927
rect 19518 3924 19524 3936
rect 19475 3896 19524 3924
rect 19475 3893 19487 3896
rect 19429 3887 19487 3893
rect 19518 3884 19524 3896
rect 19576 3884 19582 3936
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 4614 3680 4620 3732
rect 4672 3720 4678 3732
rect 5902 3720 5908 3732
rect 4672 3692 5908 3720
rect 4672 3680 4678 3692
rect 5902 3680 5908 3692
rect 5960 3680 5966 3732
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 12802 3720 12808 3732
rect 10100 3692 12808 3720
rect 10100 3680 10106 3692
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 12897 3723 12955 3729
rect 12897 3689 12909 3723
rect 12943 3720 12955 3723
rect 14734 3720 14740 3732
rect 12943 3692 14740 3720
rect 12943 3689 12955 3692
rect 12897 3683 12955 3689
rect 14734 3680 14740 3692
rect 14792 3680 14798 3732
rect 14844 3692 17172 3720
rect 9214 3612 9220 3664
rect 9272 3652 9278 3664
rect 11054 3652 11060 3664
rect 9272 3624 11060 3652
rect 9272 3612 9278 3624
rect 11054 3612 11060 3624
rect 11112 3612 11118 3664
rect 5626 3544 5632 3596
rect 5684 3584 5690 3596
rect 10226 3584 10232 3596
rect 5684 3556 10232 3584
rect 5684 3544 5690 3556
rect 10226 3544 10232 3556
rect 10284 3544 10290 3596
rect 10686 3584 10692 3596
rect 10647 3556 10692 3584
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 10870 3544 10876 3596
rect 10928 3584 10934 3596
rect 13814 3584 13820 3596
rect 10928 3556 13820 3584
rect 10928 3544 10934 3556
rect 13814 3544 13820 3556
rect 13872 3544 13878 3596
rect 14844 3593 14872 3692
rect 15470 3612 15476 3664
rect 15528 3652 15534 3664
rect 15528 3624 16804 3652
rect 15528 3612 15534 3624
rect 14829 3587 14887 3593
rect 14829 3553 14841 3587
rect 14875 3553 14887 3587
rect 14829 3547 14887 3553
rect 15102 3544 15108 3596
rect 15160 3584 15166 3596
rect 15749 3587 15807 3593
rect 15749 3584 15761 3587
rect 15160 3556 15761 3584
rect 15160 3544 15166 3556
rect 15749 3553 15761 3556
rect 15795 3553 15807 3587
rect 15749 3547 15807 3553
rect 16114 3544 16120 3596
rect 16172 3584 16178 3596
rect 16776 3593 16804 3624
rect 16669 3587 16727 3593
rect 16669 3584 16681 3587
rect 16172 3556 16681 3584
rect 16172 3544 16178 3556
rect 16669 3553 16681 3556
rect 16715 3553 16727 3587
rect 16669 3547 16727 3553
rect 16761 3587 16819 3593
rect 16761 3553 16773 3587
rect 16807 3553 16819 3587
rect 17144 3584 17172 3692
rect 17218 3680 17224 3732
rect 17276 3720 17282 3732
rect 17589 3723 17647 3729
rect 17589 3720 17601 3723
rect 17276 3692 17601 3720
rect 17276 3680 17282 3692
rect 17589 3689 17601 3692
rect 17635 3689 17647 3723
rect 19610 3720 19616 3732
rect 19571 3692 19616 3720
rect 17589 3683 17647 3689
rect 19610 3680 19616 3692
rect 19668 3680 19674 3732
rect 20806 3680 20812 3732
rect 20864 3720 20870 3732
rect 21269 3723 21327 3729
rect 21269 3720 21281 3723
rect 20864 3692 21281 3720
rect 20864 3680 20870 3692
rect 21269 3689 21281 3692
rect 21315 3689 21327 3723
rect 21269 3683 21327 3689
rect 18325 3655 18383 3661
rect 18325 3621 18337 3655
rect 18371 3652 18383 3655
rect 20254 3652 20260 3664
rect 18371 3624 20260 3652
rect 18371 3621 18383 3624
rect 18325 3615 18383 3621
rect 20254 3612 20260 3624
rect 20312 3612 20318 3664
rect 22094 3652 22100 3664
rect 20364 3624 22100 3652
rect 20364 3593 20392 3624
rect 22094 3612 22100 3624
rect 22152 3612 22158 3664
rect 20349 3587 20407 3593
rect 20349 3584 20361 3587
rect 17144 3556 20361 3584
rect 16761 3547 16819 3553
rect 20349 3553 20361 3556
rect 20395 3553 20407 3587
rect 20349 3547 20407 3553
rect 20809 3587 20867 3593
rect 20809 3553 20821 3587
rect 20855 3584 20867 3587
rect 22370 3584 22376 3596
rect 20855 3556 22376 3584
rect 20855 3553 20867 3556
rect 20809 3547 20867 3553
rect 10962 3516 10968 3528
rect 10923 3488 10968 3516
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 12066 3476 12072 3528
rect 12124 3516 12130 3528
rect 12161 3519 12219 3525
rect 12161 3516 12173 3519
rect 12124 3488 12173 3516
rect 12124 3476 12130 3488
rect 12161 3485 12173 3488
rect 12207 3485 12219 3519
rect 12161 3479 12219 3485
rect 12434 3476 12440 3528
rect 12492 3516 12498 3528
rect 12713 3519 12771 3525
rect 12713 3516 12725 3519
rect 12492 3488 12725 3516
rect 12492 3476 12498 3488
rect 12713 3485 12725 3488
rect 12759 3485 12771 3519
rect 12713 3479 12771 3485
rect 13265 3519 13323 3525
rect 13265 3485 13277 3519
rect 13311 3516 13323 3519
rect 13354 3516 13360 3528
rect 13311 3488 13360 3516
rect 13311 3485 13323 3488
rect 13265 3479 13323 3485
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 15378 3516 15384 3528
rect 13464 3488 15384 3516
rect 9953 3451 10011 3457
rect 9953 3417 9965 3451
rect 9999 3448 10011 3451
rect 11054 3448 11060 3460
rect 9999 3420 11060 3448
rect 9999 3417 10011 3420
rect 9953 3411 10011 3417
rect 11054 3408 11060 3420
rect 11112 3408 11118 3460
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 11241 3451 11299 3457
rect 11241 3448 11253 3451
rect 11204 3420 11253 3448
rect 11204 3408 11210 3420
rect 11241 3417 11253 3420
rect 11287 3417 11299 3451
rect 11241 3411 11299 3417
rect 11885 3451 11943 3457
rect 11885 3417 11897 3451
rect 11931 3448 11943 3451
rect 11974 3448 11980 3460
rect 11931 3420 11980 3448
rect 11931 3417 11943 3420
rect 11885 3411 11943 3417
rect 11974 3408 11980 3420
rect 12032 3408 12038 3460
rect 7006 3340 7012 3392
rect 7064 3380 7070 3392
rect 13078 3380 13084 3392
rect 7064 3352 13084 3380
rect 7064 3340 7070 3352
rect 13078 3340 13084 3352
rect 13136 3340 13142 3392
rect 13464 3389 13492 3488
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 15562 3476 15568 3528
rect 15620 3516 15626 3528
rect 15657 3519 15715 3525
rect 15657 3516 15669 3519
rect 15620 3488 15669 3516
rect 15620 3476 15626 3488
rect 15657 3485 15669 3488
rect 15703 3485 15715 3519
rect 15657 3479 15715 3485
rect 16482 3476 16488 3528
rect 16540 3516 16546 3528
rect 16577 3519 16635 3525
rect 16577 3516 16589 3519
rect 16540 3488 16589 3516
rect 16540 3476 16546 3488
rect 16577 3485 16589 3488
rect 16623 3485 16635 3519
rect 16577 3479 16635 3485
rect 17126 3476 17132 3528
rect 17184 3516 17190 3528
rect 17221 3519 17279 3525
rect 17221 3516 17233 3519
rect 17184 3488 17233 3516
rect 17184 3476 17190 3488
rect 17221 3485 17233 3488
rect 17267 3485 17279 3519
rect 17221 3479 17279 3485
rect 17954 3476 17960 3528
rect 18012 3516 18018 3528
rect 18141 3519 18199 3525
rect 18141 3516 18153 3519
rect 18012 3488 18153 3516
rect 18012 3476 18018 3488
rect 18141 3485 18153 3488
rect 18187 3485 18199 3519
rect 20824 3516 20852 3547
rect 22370 3544 22376 3556
rect 22428 3544 22434 3596
rect 18141 3479 18199 3485
rect 18248 3488 20852 3516
rect 14553 3451 14611 3457
rect 14553 3417 14565 3451
rect 14599 3448 14611 3451
rect 14599 3420 16252 3448
rect 14599 3417 14611 3420
rect 14553 3411 14611 3417
rect 13449 3383 13507 3389
rect 13449 3349 13461 3383
rect 13495 3349 13507 3383
rect 13449 3343 13507 3349
rect 13538 3340 13544 3392
rect 13596 3380 13602 3392
rect 14185 3383 14243 3389
rect 14185 3380 14197 3383
rect 13596 3352 14197 3380
rect 13596 3340 13602 3352
rect 14185 3349 14197 3352
rect 14231 3349 14243 3383
rect 14185 3343 14243 3349
rect 14645 3383 14703 3389
rect 14645 3349 14657 3383
rect 14691 3380 14703 3383
rect 14826 3380 14832 3392
rect 14691 3352 14832 3380
rect 14691 3349 14703 3352
rect 14645 3343 14703 3349
rect 14826 3340 14832 3352
rect 14884 3340 14890 3392
rect 15197 3383 15255 3389
rect 15197 3349 15209 3383
rect 15243 3380 15255 3383
rect 15286 3380 15292 3392
rect 15243 3352 15292 3380
rect 15243 3349 15255 3352
rect 15197 3343 15255 3349
rect 15286 3340 15292 3352
rect 15344 3340 15350 3392
rect 15565 3383 15623 3389
rect 15565 3349 15577 3383
rect 15611 3380 15623 3383
rect 15746 3380 15752 3392
rect 15611 3352 15752 3380
rect 15611 3349 15623 3352
rect 15565 3343 15623 3349
rect 15746 3340 15752 3352
rect 15804 3340 15810 3392
rect 16224 3389 16252 3420
rect 16298 3408 16304 3460
rect 16356 3448 16362 3460
rect 18248 3448 18276 3488
rect 19981 3451 20039 3457
rect 19981 3448 19993 3451
rect 16356 3420 18276 3448
rect 19352 3420 19993 3448
rect 16356 3408 16362 3420
rect 19352 3392 19380 3420
rect 19981 3417 19993 3420
rect 20027 3448 20039 3451
rect 20070 3448 20076 3460
rect 20027 3420 20076 3448
rect 20027 3417 20039 3420
rect 19981 3411 20039 3417
rect 20070 3408 20076 3420
rect 20128 3408 20134 3460
rect 16209 3383 16267 3389
rect 16209 3349 16221 3383
rect 16255 3349 16267 3383
rect 16209 3343 16267 3349
rect 16390 3340 16396 3392
rect 16448 3380 16454 3392
rect 18693 3383 18751 3389
rect 18693 3380 18705 3383
rect 16448 3352 18705 3380
rect 16448 3340 16454 3352
rect 18693 3349 18705 3352
rect 18739 3380 18751 3383
rect 18782 3380 18788 3392
rect 18739 3352 18788 3380
rect 18739 3349 18751 3352
rect 18693 3343 18751 3349
rect 18782 3340 18788 3352
rect 18840 3340 18846 3392
rect 19334 3380 19340 3392
rect 19295 3352 19340 3380
rect 19334 3340 19340 3352
rect 19392 3340 19398 3392
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 8478 3136 8484 3188
rect 8536 3176 8542 3188
rect 9401 3179 9459 3185
rect 9401 3176 9413 3179
rect 8536 3148 9413 3176
rect 8536 3136 8542 3148
rect 9401 3145 9413 3148
rect 9447 3145 9459 3179
rect 9858 3176 9864 3188
rect 9819 3148 9864 3176
rect 9401 3139 9459 3145
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 10134 3176 10140 3188
rect 10095 3148 10140 3176
rect 10134 3136 10140 3148
rect 10192 3136 10198 3188
rect 10594 3176 10600 3188
rect 10555 3148 10600 3176
rect 10594 3136 10600 3148
rect 10652 3136 10658 3188
rect 13446 3136 13452 3188
rect 13504 3176 13510 3188
rect 13817 3179 13875 3185
rect 13817 3176 13829 3179
rect 13504 3148 13829 3176
rect 13504 3136 13510 3148
rect 13817 3145 13829 3148
rect 13863 3145 13875 3179
rect 14182 3176 14188 3188
rect 14095 3148 14188 3176
rect 13817 3139 13875 3145
rect 14182 3136 14188 3148
rect 14240 3176 14246 3188
rect 14826 3176 14832 3188
rect 14240 3148 14688 3176
rect 14787 3148 14832 3176
rect 14240 3136 14246 3148
rect 10152 3108 10180 3136
rect 12066 3108 12072 3120
rect 10152 3080 12072 3108
rect 12066 3068 12072 3080
rect 12124 3068 12130 3120
rect 13354 3108 13360 3120
rect 12406 3080 13360 3108
rect 11146 3040 11152 3052
rect 11107 3012 11152 3040
rect 11146 3000 11152 3012
rect 11204 3000 11210 3052
rect 11882 3040 11888 3052
rect 11843 3012 11888 3040
rect 11882 3000 11888 3012
rect 11940 3000 11946 3052
rect 12406 3040 12434 3080
rect 13354 3068 13360 3080
rect 13412 3108 13418 3120
rect 14277 3111 14335 3117
rect 14277 3108 14289 3111
rect 13412 3080 14289 3108
rect 13412 3068 13418 3080
rect 14277 3077 14289 3080
rect 14323 3077 14335 3111
rect 14660 3108 14688 3148
rect 14826 3136 14832 3148
rect 14884 3136 14890 3188
rect 15286 3176 15292 3188
rect 15247 3148 15292 3176
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 17681 3179 17739 3185
rect 17681 3145 17693 3179
rect 17727 3145 17739 3179
rect 17681 3139 17739 3145
rect 14918 3108 14924 3120
rect 14660 3080 14924 3108
rect 14277 3071 14335 3077
rect 14918 3068 14924 3080
rect 14976 3068 14982 3120
rect 15194 3108 15200 3120
rect 15155 3080 15200 3108
rect 15194 3068 15200 3080
rect 15252 3068 15258 3120
rect 17696 3108 17724 3139
rect 18322 3136 18328 3188
rect 18380 3176 18386 3188
rect 18598 3176 18604 3188
rect 18380 3148 18604 3176
rect 18380 3136 18386 3148
rect 18598 3136 18604 3148
rect 18656 3136 18662 3188
rect 18785 3179 18843 3185
rect 18785 3145 18797 3179
rect 18831 3176 18843 3179
rect 22462 3176 22468 3188
rect 18831 3148 22468 3176
rect 18831 3145 18843 3148
rect 18785 3139 18843 3145
rect 22462 3136 22468 3148
rect 22520 3136 22526 3188
rect 20714 3108 20720 3120
rect 17696 3080 20720 3108
rect 20714 3068 20720 3080
rect 20772 3068 20778 3120
rect 11992 3012 12434 3040
rect 13265 3043 13323 3049
rect 3878 2932 3884 2984
rect 3936 2972 3942 2984
rect 11517 2975 11575 2981
rect 11517 2972 11529 2975
rect 3936 2944 11529 2972
rect 3936 2932 3942 2944
rect 11517 2941 11529 2944
rect 11563 2972 11575 2975
rect 11992 2972 12020 3012
rect 13265 3009 13277 3043
rect 13311 3040 13323 3043
rect 13538 3040 13544 3052
rect 13311 3012 13544 3040
rect 13311 3009 13323 3012
rect 13265 3003 13323 3009
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 15654 3040 15660 3052
rect 14476 3012 15660 3040
rect 12158 2972 12164 2984
rect 11563 2944 12020 2972
rect 12119 2944 12164 2972
rect 11563 2941 11575 2944
rect 11517 2935 11575 2941
rect 12158 2932 12164 2944
rect 12216 2932 12222 2984
rect 13081 2975 13139 2981
rect 13081 2941 13093 2975
rect 13127 2972 13139 2975
rect 13814 2972 13820 2984
rect 13127 2944 13820 2972
rect 13127 2941 13139 2944
rect 13081 2935 13139 2941
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 14476 2981 14504 3012
rect 15654 3000 15660 3012
rect 15712 3000 15718 3052
rect 15838 3000 15844 3052
rect 15896 3040 15902 3052
rect 15933 3043 15991 3049
rect 15933 3040 15945 3043
rect 15896 3012 15945 3040
rect 15896 3000 15902 3012
rect 15933 3009 15945 3012
rect 15979 3009 15991 3043
rect 16942 3040 16948 3052
rect 16903 3012 16948 3040
rect 15933 3003 15991 3009
rect 16942 3000 16948 3012
rect 17000 3000 17006 3052
rect 17494 3040 17500 3052
rect 17455 3012 17500 3040
rect 17494 3000 17500 3012
rect 17552 3000 17558 3052
rect 17862 3000 17868 3052
rect 17920 3040 17926 3052
rect 18325 3043 18383 3049
rect 18325 3040 18337 3043
rect 17920 3012 18337 3040
rect 17920 3000 17926 3012
rect 18325 3009 18337 3012
rect 18371 3009 18383 3043
rect 18325 3003 18383 3009
rect 18601 3043 18659 3049
rect 18601 3009 18613 3043
rect 18647 3009 18659 3043
rect 18601 3003 18659 3009
rect 14461 2975 14519 2981
rect 14461 2941 14473 2975
rect 14507 2941 14519 2975
rect 15470 2972 15476 2984
rect 15431 2944 15476 2972
rect 14461 2935 14519 2941
rect 15470 2932 15476 2944
rect 15528 2932 15534 2984
rect 17218 2932 17224 2984
rect 17276 2972 17282 2984
rect 18616 2972 18644 3003
rect 19058 3000 19064 3052
rect 19116 3040 19122 3052
rect 19153 3043 19211 3049
rect 19153 3040 19165 3043
rect 19116 3012 19165 3040
rect 19116 3000 19122 3012
rect 19153 3009 19165 3012
rect 19199 3009 19211 3043
rect 19153 3003 19211 3009
rect 19334 3000 19340 3052
rect 19392 3040 19398 3052
rect 19705 3043 19763 3049
rect 19705 3040 19717 3043
rect 19392 3012 19717 3040
rect 19392 3000 19398 3012
rect 19705 3009 19717 3012
rect 19751 3009 19763 3043
rect 19705 3003 19763 3009
rect 20438 3000 20444 3052
rect 20496 3040 20502 3052
rect 20809 3043 20867 3049
rect 20809 3040 20821 3043
rect 20496 3012 20821 3040
rect 20496 3000 20502 3012
rect 20809 3009 20821 3012
rect 20855 3009 20867 3043
rect 20809 3003 20867 3009
rect 17276 2944 18644 2972
rect 17276 2932 17282 2944
rect 19518 2932 19524 2984
rect 19576 2972 19582 2984
rect 20257 2975 20315 2981
rect 20257 2972 20269 2975
rect 19576 2944 20269 2972
rect 19576 2932 19582 2944
rect 20257 2941 20269 2944
rect 20303 2941 20315 2975
rect 20257 2935 20315 2941
rect 10965 2907 11023 2913
rect 10965 2873 10977 2907
rect 11011 2904 11023 2907
rect 11882 2904 11888 2916
rect 11011 2876 11888 2904
rect 11011 2873 11023 2876
rect 10965 2867 11023 2873
rect 11882 2864 11888 2876
rect 11940 2864 11946 2916
rect 16117 2907 16175 2913
rect 16117 2873 16129 2907
rect 16163 2904 16175 2907
rect 16163 2876 16896 2904
rect 16163 2873 16175 2876
rect 16117 2867 16175 2873
rect 382 2796 388 2848
rect 440 2836 446 2848
rect 8294 2836 8300 2848
rect 440 2808 8300 2836
rect 440 2796 446 2808
rect 8294 2796 8300 2808
rect 8352 2796 8358 2848
rect 10686 2796 10692 2848
rect 10744 2836 10750 2848
rect 11790 2836 11796 2848
rect 10744 2808 11796 2836
rect 10744 2796 10750 2808
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 16390 2796 16396 2848
rect 16448 2836 16454 2848
rect 16761 2839 16819 2845
rect 16761 2836 16773 2839
rect 16448 2808 16773 2836
rect 16448 2796 16454 2808
rect 16761 2805 16773 2808
rect 16807 2805 16819 2839
rect 16868 2836 16896 2876
rect 16942 2864 16948 2916
rect 17000 2904 17006 2916
rect 18141 2907 18199 2913
rect 18141 2904 18153 2907
rect 17000 2876 18153 2904
rect 17000 2864 17006 2876
rect 18141 2873 18153 2876
rect 18187 2873 18199 2907
rect 18141 2867 18199 2873
rect 18598 2864 18604 2916
rect 18656 2904 18662 2916
rect 19337 2907 19395 2913
rect 19337 2904 19349 2907
rect 18656 2876 19349 2904
rect 18656 2864 18662 2876
rect 19337 2873 19349 2876
rect 19383 2873 19395 2907
rect 19337 2867 19395 2873
rect 19889 2907 19947 2913
rect 19889 2873 19901 2907
rect 19935 2904 19947 2907
rect 21358 2904 21364 2916
rect 19935 2876 21364 2904
rect 19935 2873 19947 2876
rect 19889 2867 19947 2873
rect 21358 2864 21364 2876
rect 21416 2864 21422 2916
rect 17494 2836 17500 2848
rect 16868 2808 17500 2836
rect 16761 2799 16819 2805
rect 17494 2796 17500 2808
rect 17552 2796 17558 2848
rect 20993 2839 21051 2845
rect 20993 2805 21005 2839
rect 21039 2836 21051 2839
rect 21542 2836 21548 2848
rect 21039 2808 21548 2836
rect 21039 2805 21051 2808
rect 20993 2799 21051 2805
rect 21542 2796 21548 2808
rect 21600 2796 21606 2848
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 10226 2592 10232 2644
rect 10284 2632 10290 2644
rect 10689 2635 10747 2641
rect 10689 2632 10701 2635
rect 10284 2604 10701 2632
rect 10284 2592 10290 2604
rect 10689 2601 10701 2604
rect 10735 2601 10747 2635
rect 11146 2632 11152 2644
rect 11107 2604 11152 2632
rect 10689 2595 10747 2601
rect 10413 2567 10471 2573
rect 10413 2533 10425 2567
rect 10459 2564 10471 2567
rect 10502 2564 10508 2576
rect 10459 2536 10508 2564
rect 10459 2533 10471 2536
rect 10413 2527 10471 2533
rect 10502 2524 10508 2536
rect 10560 2524 10566 2576
rect 10704 2496 10732 2595
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 11701 2635 11759 2641
rect 11701 2601 11713 2635
rect 11747 2632 11759 2635
rect 11790 2632 11796 2644
rect 11747 2604 11796 2632
rect 11747 2601 11759 2604
rect 11701 2595 11759 2601
rect 11790 2592 11796 2604
rect 11848 2592 11854 2644
rect 13170 2592 13176 2644
rect 13228 2632 13234 2644
rect 13633 2635 13691 2641
rect 13633 2632 13645 2635
rect 13228 2604 13645 2632
rect 13228 2592 13234 2604
rect 13633 2601 13645 2604
rect 13679 2601 13691 2635
rect 13633 2595 13691 2601
rect 14918 2592 14924 2644
rect 14976 2632 14982 2644
rect 15933 2635 15991 2641
rect 15933 2632 15945 2635
rect 14976 2604 15945 2632
rect 14976 2592 14982 2604
rect 15933 2601 15945 2604
rect 15979 2601 15991 2635
rect 15933 2595 15991 2601
rect 16206 2592 16212 2644
rect 16264 2632 16270 2644
rect 17129 2635 17187 2641
rect 17129 2632 17141 2635
rect 16264 2604 17141 2632
rect 16264 2592 16270 2604
rect 17129 2601 17141 2604
rect 17175 2601 17187 2635
rect 17129 2595 17187 2601
rect 18414 2592 18420 2644
rect 18472 2632 18478 2644
rect 18693 2635 18751 2641
rect 18693 2632 18705 2635
rect 18472 2604 18705 2632
rect 18472 2592 18478 2604
rect 18693 2601 18705 2604
rect 18739 2601 18751 2635
rect 18693 2595 18751 2601
rect 18874 2592 18880 2644
rect 18932 2632 18938 2644
rect 19613 2635 19671 2641
rect 19613 2632 19625 2635
rect 18932 2604 19625 2632
rect 18932 2592 18938 2604
rect 19613 2601 19625 2604
rect 19659 2601 19671 2635
rect 19978 2632 19984 2644
rect 19939 2604 19984 2632
rect 19613 2595 19671 2601
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 20714 2592 20720 2644
rect 20772 2632 20778 2644
rect 21269 2635 21327 2641
rect 21269 2632 21281 2635
rect 20772 2604 21281 2632
rect 20772 2592 20778 2604
rect 21269 2601 21281 2604
rect 21315 2601 21327 2635
rect 21269 2595 21327 2601
rect 15105 2567 15163 2573
rect 13096 2536 14964 2564
rect 13096 2496 13124 2536
rect 10704 2468 13124 2496
rect 14936 2496 14964 2536
rect 15105 2533 15117 2567
rect 15151 2564 15163 2567
rect 15838 2564 15844 2576
rect 15151 2536 15844 2564
rect 15151 2533 15163 2536
rect 15105 2527 15163 2533
rect 15838 2524 15844 2536
rect 15896 2524 15902 2576
rect 16853 2567 16911 2573
rect 16853 2533 16865 2567
rect 16899 2564 16911 2567
rect 17402 2564 17408 2576
rect 16899 2536 17408 2564
rect 16899 2533 16911 2536
rect 16853 2527 16911 2533
rect 17402 2524 17408 2536
rect 17460 2524 17466 2576
rect 18325 2567 18383 2573
rect 18325 2533 18337 2567
rect 18371 2564 18383 2567
rect 19702 2564 19708 2576
rect 18371 2536 19708 2564
rect 18371 2533 18383 2536
rect 18325 2527 18383 2533
rect 19702 2524 19708 2536
rect 19760 2524 19766 2576
rect 15562 2496 15568 2508
rect 14936 2468 15568 2496
rect 11974 2428 11980 2440
rect 11935 2400 11980 2428
rect 11974 2388 11980 2400
rect 12032 2388 12038 2440
rect 12158 2388 12164 2440
rect 12216 2428 12222 2440
rect 12529 2431 12587 2437
rect 12529 2428 12541 2431
rect 12216 2400 12541 2428
rect 12216 2388 12222 2400
rect 12529 2397 12541 2400
rect 12575 2397 12587 2431
rect 12529 2391 12587 2397
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 10045 2363 10103 2369
rect 10045 2329 10057 2363
rect 10091 2360 10103 2363
rect 11054 2360 11060 2372
rect 10091 2332 11060 2360
rect 10091 2329 10103 2332
rect 10045 2323 10103 2329
rect 11054 2320 11060 2332
rect 11112 2320 11118 2372
rect 11790 2320 11796 2372
rect 11848 2360 11854 2372
rect 13096 2360 13124 2391
rect 13814 2388 13820 2440
rect 13872 2428 13878 2440
rect 14936 2437 14964 2468
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 16022 2456 16028 2508
rect 16080 2496 16086 2508
rect 16209 2499 16267 2505
rect 16209 2496 16221 2499
rect 16080 2468 16221 2496
rect 16080 2456 16086 2468
rect 16209 2465 16221 2468
rect 16255 2496 16267 2499
rect 17497 2499 17555 2505
rect 17497 2496 17509 2499
rect 16255 2468 17509 2496
rect 16255 2465 16267 2468
rect 16209 2459 16267 2465
rect 17497 2465 17509 2468
rect 17543 2465 17555 2499
rect 17497 2459 17555 2465
rect 17770 2456 17776 2508
rect 17828 2496 17834 2508
rect 19245 2499 19303 2505
rect 19245 2496 19257 2499
rect 17828 2468 19257 2496
rect 17828 2456 17834 2468
rect 19245 2465 19257 2468
rect 19291 2465 19303 2499
rect 19245 2459 19303 2465
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 13872 2400 14105 2428
rect 13872 2388 13878 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 14921 2431 14979 2437
rect 14921 2397 14933 2431
rect 14967 2397 14979 2431
rect 14921 2391 14979 2397
rect 15930 2388 15936 2440
rect 15988 2428 15994 2440
rect 18141 2431 18199 2437
rect 18141 2428 18153 2431
rect 15988 2400 18153 2428
rect 15988 2388 15994 2400
rect 18141 2397 18153 2400
rect 18187 2397 18199 2431
rect 18141 2391 18199 2397
rect 18506 2388 18512 2440
rect 18564 2428 18570 2440
rect 20717 2431 20775 2437
rect 20717 2428 20729 2431
rect 18564 2400 20729 2428
rect 18564 2388 18570 2400
rect 20717 2397 20729 2400
rect 20763 2397 20775 2431
rect 20717 2391 20775 2397
rect 11848 2332 13124 2360
rect 11848 2320 11854 2332
rect 15746 2320 15752 2372
rect 15804 2360 15810 2372
rect 19150 2360 19156 2372
rect 15804 2332 19156 2360
rect 15804 2320 15810 2332
rect 19150 2320 19156 2332
rect 19208 2320 19214 2372
rect 12161 2295 12219 2301
rect 12161 2261 12173 2295
rect 12207 2292 12219 2295
rect 12526 2292 12532 2304
rect 12207 2264 12532 2292
rect 12207 2261 12219 2264
rect 12161 2255 12219 2261
rect 12526 2252 12532 2264
rect 12584 2252 12590 2304
rect 12713 2295 12771 2301
rect 12713 2261 12725 2295
rect 12759 2292 12771 2295
rect 13078 2292 13084 2304
rect 12759 2264 13084 2292
rect 12759 2261 12771 2264
rect 12713 2255 12771 2261
rect 13078 2252 13084 2264
rect 13136 2252 13142 2304
rect 13265 2295 13323 2301
rect 13265 2261 13277 2295
rect 13311 2292 13323 2295
rect 13538 2292 13544 2304
rect 13311 2264 13544 2292
rect 13311 2261 13323 2264
rect 13265 2255 13323 2261
rect 13538 2252 13544 2264
rect 13596 2252 13602 2304
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 14240 2264 14289 2292
rect 14240 2252 14246 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 15470 2292 15476 2304
rect 15431 2264 15476 2292
rect 14277 2255 14335 2261
rect 15470 2252 15476 2264
rect 15528 2252 15534 2304
rect 15562 2252 15568 2304
rect 15620 2292 15626 2304
rect 17034 2292 17040 2304
rect 15620 2264 17040 2292
rect 15620 2252 15626 2264
rect 17034 2252 17040 2264
rect 17092 2252 17098 2304
rect 18690 2252 18696 2304
rect 18748 2292 18754 2304
rect 20349 2295 20407 2301
rect 20349 2292 20361 2295
rect 18748 2264 20361 2292
rect 18748 2252 18754 2264
rect 20349 2261 20361 2264
rect 20395 2261 20407 2295
rect 20349 2255 20407 2261
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
rect 11054 2048 11060 2100
rect 11112 2088 11118 2100
rect 12250 2088 12256 2100
rect 11112 2060 12256 2088
rect 11112 2048 11118 2060
rect 12250 2048 12256 2060
rect 12308 2088 12314 2100
rect 15930 2088 15936 2100
rect 12308 2060 15936 2088
rect 12308 2048 12314 2060
rect 15930 2048 15936 2060
rect 15988 2048 15994 2100
rect 14642 1980 14648 2032
rect 14700 2020 14706 2032
rect 15746 2020 15752 2032
rect 14700 1992 15752 2020
rect 14700 1980 14706 1992
rect 15746 1980 15752 1992
rect 15804 1980 15810 2032
rect 10502 1912 10508 1964
rect 10560 1952 10566 1964
rect 15470 1952 15476 1964
rect 10560 1924 15476 1952
rect 10560 1912 10566 1924
rect 15470 1912 15476 1924
rect 15528 1912 15534 1964
<< via1 >>
rect 10232 21020 10284 21072
rect 11980 21020 12032 21072
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 6552 20476 6604 20528
rect 6736 20408 6788 20460
rect 7748 20451 7800 20460
rect 7748 20417 7757 20451
rect 7757 20417 7791 20451
rect 7791 20417 7800 20451
rect 7748 20408 7800 20417
rect 11704 20544 11756 20596
rect 18604 20544 18656 20596
rect 18696 20587 18748 20596
rect 18696 20553 18705 20587
rect 18705 20553 18739 20587
rect 18739 20553 18748 20587
rect 18696 20544 18748 20553
rect 21364 20544 21416 20596
rect 10232 20408 10284 20460
rect 10508 20451 10560 20460
rect 10508 20417 10517 20451
rect 10517 20417 10551 20451
rect 10551 20417 10560 20451
rect 10508 20408 10560 20417
rect 12624 20408 12676 20460
rect 7380 20340 7432 20392
rect 7564 20340 7616 20392
rect 14648 20408 14700 20460
rect 15660 20451 15712 20460
rect 15660 20417 15669 20451
rect 15669 20417 15703 20451
rect 15703 20417 15712 20451
rect 15660 20408 15712 20417
rect 5632 20247 5684 20256
rect 5632 20213 5641 20247
rect 5641 20213 5675 20247
rect 5675 20213 5684 20247
rect 5632 20204 5684 20213
rect 6552 20204 6604 20256
rect 7288 20204 7340 20256
rect 8392 20204 8444 20256
rect 8576 20204 8628 20256
rect 10324 20204 10376 20256
rect 17592 20476 17644 20528
rect 18144 20408 18196 20460
rect 18420 20408 18472 20460
rect 13728 20315 13780 20324
rect 13728 20281 13737 20315
rect 13737 20281 13771 20315
rect 13771 20281 13780 20315
rect 13728 20272 13780 20281
rect 10968 20204 11020 20256
rect 12164 20247 12216 20256
rect 12164 20213 12173 20247
rect 12173 20213 12207 20247
rect 12207 20213 12216 20247
rect 12164 20204 12216 20213
rect 12716 20204 12768 20256
rect 16764 20340 16816 20392
rect 20260 20476 20312 20528
rect 18880 20408 18932 20460
rect 16304 20272 16356 20324
rect 20812 20408 20864 20460
rect 21088 20451 21140 20460
rect 21088 20417 21106 20451
rect 21106 20417 21140 20451
rect 21088 20408 21140 20417
rect 21364 20383 21416 20392
rect 21364 20349 21373 20383
rect 21373 20349 21407 20383
rect 21407 20349 21416 20383
rect 21364 20340 21416 20349
rect 14648 20247 14700 20256
rect 14648 20213 14657 20247
rect 14657 20213 14691 20247
rect 14691 20213 14700 20247
rect 14648 20204 14700 20213
rect 15936 20204 15988 20256
rect 16212 20247 16264 20256
rect 16212 20213 16221 20247
rect 16221 20213 16255 20247
rect 16255 20213 16264 20247
rect 16212 20204 16264 20213
rect 17960 20204 18012 20256
rect 18144 20204 18196 20256
rect 20168 20272 20220 20324
rect 19984 20247 20036 20256
rect 19984 20213 19993 20247
rect 19993 20213 20027 20247
rect 20027 20213 20036 20247
rect 19984 20204 20036 20213
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 13084 20000 13136 20052
rect 5724 19932 5776 19984
rect 6736 19907 6788 19916
rect 6736 19873 6745 19907
rect 6745 19873 6779 19907
rect 6779 19873 6788 19907
rect 6736 19864 6788 19873
rect 4620 19703 4672 19712
rect 4620 19669 4629 19703
rect 4629 19669 4663 19703
rect 4663 19669 4672 19703
rect 4620 19660 4672 19669
rect 7012 19839 7064 19848
rect 7012 19805 7021 19839
rect 7021 19805 7055 19839
rect 7055 19805 7064 19839
rect 7012 19796 7064 19805
rect 7196 19796 7248 19848
rect 11980 19864 12032 19916
rect 10968 19796 11020 19848
rect 7104 19728 7156 19780
rect 5172 19660 5224 19712
rect 5724 19703 5776 19712
rect 5724 19669 5733 19703
rect 5733 19669 5767 19703
rect 5767 19669 5776 19703
rect 5724 19660 5776 19669
rect 6920 19660 6972 19712
rect 7380 19703 7432 19712
rect 7380 19669 7389 19703
rect 7389 19669 7423 19703
rect 7423 19669 7432 19703
rect 7380 19660 7432 19669
rect 9312 19660 9364 19712
rect 10324 19771 10376 19780
rect 10324 19737 10342 19771
rect 10342 19737 10376 19771
rect 10324 19728 10376 19737
rect 10692 19728 10744 19780
rect 15476 19839 15528 19848
rect 11060 19660 11112 19712
rect 11520 19728 11572 19780
rect 13636 19728 13688 19780
rect 11428 19660 11480 19712
rect 12256 19703 12308 19712
rect 12256 19669 12265 19703
rect 12265 19669 12299 19703
rect 12299 19669 12308 19703
rect 12256 19660 12308 19669
rect 12532 19703 12584 19712
rect 12532 19669 12541 19703
rect 12541 19669 12575 19703
rect 12575 19669 12584 19703
rect 12532 19660 12584 19669
rect 13820 19660 13872 19712
rect 14648 19728 14700 19780
rect 15476 19805 15485 19839
rect 15485 19805 15519 19839
rect 15519 19805 15528 19839
rect 15476 19796 15528 19805
rect 15568 19796 15620 19848
rect 17592 19932 17644 19984
rect 18052 20000 18104 20052
rect 18696 20000 18748 20052
rect 21088 20000 21140 20052
rect 17040 19796 17092 19848
rect 17316 19796 17368 19848
rect 18236 19839 18288 19848
rect 18236 19805 18245 19839
rect 18245 19805 18279 19839
rect 18279 19805 18288 19839
rect 18236 19796 18288 19805
rect 16948 19728 17000 19780
rect 16396 19660 16448 19712
rect 18420 19864 18472 19916
rect 21364 19907 21416 19916
rect 21364 19873 21373 19907
rect 21373 19873 21407 19907
rect 21407 19873 21416 19907
rect 21364 19864 21416 19873
rect 18788 19839 18840 19848
rect 18788 19805 18797 19839
rect 18797 19805 18831 19839
rect 18831 19805 18840 19839
rect 18788 19796 18840 19805
rect 18420 19728 18472 19780
rect 19708 19728 19760 19780
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 5356 19456 5408 19508
rect 6828 19456 6880 19508
rect 4988 19388 5040 19440
rect 7748 19388 7800 19440
rect 5632 19363 5684 19372
rect 5632 19329 5641 19363
rect 5641 19329 5675 19363
rect 5675 19329 5684 19363
rect 5632 19320 5684 19329
rect 7840 19363 7892 19372
rect 4804 19252 4856 19304
rect 7840 19329 7849 19363
rect 7849 19329 7883 19363
rect 7883 19329 7892 19363
rect 7840 19320 7892 19329
rect 12072 19456 12124 19508
rect 8208 19388 8260 19440
rect 10324 19388 10376 19440
rect 14648 19499 14700 19508
rect 14648 19465 14657 19499
rect 14657 19465 14691 19499
rect 14691 19465 14700 19499
rect 14648 19456 14700 19465
rect 16948 19456 17000 19508
rect 18972 19456 19024 19508
rect 20536 19456 20588 19508
rect 12532 19388 12584 19440
rect 13728 19388 13780 19440
rect 6000 19252 6052 19304
rect 8208 19252 8260 19304
rect 9680 19252 9732 19304
rect 11244 19320 11296 19372
rect 15384 19388 15436 19440
rect 15476 19320 15528 19372
rect 18328 19320 18380 19372
rect 18696 19320 18748 19372
rect 19800 19363 19852 19372
rect 19800 19329 19818 19363
rect 19818 19329 19852 19363
rect 19800 19320 19852 19329
rect 11704 19252 11756 19304
rect 16028 19295 16080 19304
rect 16028 19261 16037 19295
rect 16037 19261 16071 19295
rect 16071 19261 16080 19295
rect 16028 19252 16080 19261
rect 8024 19184 8076 19236
rect 10968 19184 11020 19236
rect 5264 19159 5316 19168
rect 5264 19125 5273 19159
rect 5273 19125 5307 19159
rect 5307 19125 5316 19159
rect 5264 19116 5316 19125
rect 7288 19116 7340 19168
rect 12440 19184 12492 19236
rect 11888 19159 11940 19168
rect 11888 19125 11897 19159
rect 11897 19125 11931 19159
rect 11931 19125 11940 19159
rect 11888 19116 11940 19125
rect 12624 19116 12676 19168
rect 15844 19116 15896 19168
rect 20628 19388 20680 19440
rect 21364 19388 21416 19440
rect 20536 19363 20588 19372
rect 20536 19329 20545 19363
rect 20545 19329 20579 19363
rect 20579 19329 20588 19363
rect 20536 19320 20588 19329
rect 20260 19252 20312 19304
rect 17040 19116 17092 19168
rect 19064 19184 19116 19236
rect 20352 19116 20404 19168
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 8392 18912 8444 18964
rect 14740 18912 14792 18964
rect 15936 18912 15988 18964
rect 18696 18955 18748 18964
rect 1492 18844 1544 18896
rect 3332 18844 3384 18896
rect 7196 18776 7248 18828
rect 940 18708 992 18760
rect 4436 18708 4488 18760
rect 6828 18708 6880 18760
rect 10600 18844 10652 18896
rect 18696 18921 18705 18955
rect 18705 18921 18739 18955
rect 18739 18921 18748 18955
rect 18696 18912 18748 18921
rect 9680 18708 9732 18760
rect 10324 18751 10376 18760
rect 10324 18717 10333 18751
rect 10333 18717 10367 18751
rect 10367 18717 10376 18751
rect 10324 18708 10376 18717
rect 8116 18640 8168 18692
rect 5632 18572 5684 18624
rect 6000 18572 6052 18624
rect 7380 18572 7432 18624
rect 9864 18640 9916 18692
rect 10600 18640 10652 18692
rect 14188 18751 14240 18760
rect 14188 18717 14197 18751
rect 14197 18717 14231 18751
rect 14231 18717 14240 18751
rect 14188 18708 14240 18717
rect 16028 18708 16080 18760
rect 16304 18751 16356 18760
rect 16304 18717 16313 18751
rect 16313 18717 16347 18751
rect 16347 18717 16356 18751
rect 16304 18708 16356 18717
rect 19524 18844 19576 18896
rect 22468 18912 22520 18964
rect 20628 18819 20680 18828
rect 20628 18785 20637 18819
rect 20637 18785 20671 18819
rect 20671 18785 20680 18819
rect 20628 18776 20680 18785
rect 18696 18708 18748 18760
rect 18880 18751 18932 18760
rect 18880 18717 18889 18751
rect 18889 18717 18923 18751
rect 18923 18717 18932 18751
rect 18880 18708 18932 18717
rect 20352 18751 20404 18760
rect 20352 18717 20370 18751
rect 20370 18717 20404 18751
rect 20352 18708 20404 18717
rect 20720 18708 20772 18760
rect 12072 18640 12124 18692
rect 13268 18640 13320 18692
rect 9036 18572 9088 18624
rect 10508 18572 10560 18624
rect 10692 18615 10744 18624
rect 10692 18581 10701 18615
rect 10701 18581 10735 18615
rect 10735 18581 10744 18615
rect 10968 18615 11020 18624
rect 10692 18572 10744 18581
rect 10968 18581 10977 18615
rect 10977 18581 11011 18615
rect 11011 18581 11020 18615
rect 10968 18572 11020 18581
rect 11060 18572 11112 18624
rect 12716 18572 12768 18624
rect 12808 18572 12860 18624
rect 14464 18572 14516 18624
rect 16488 18640 16540 18692
rect 16672 18640 16724 18692
rect 19984 18640 20036 18692
rect 21180 18683 21232 18692
rect 21180 18649 21189 18683
rect 21189 18649 21223 18683
rect 21223 18649 21232 18683
rect 21180 18640 21232 18649
rect 15844 18615 15896 18624
rect 15844 18581 15853 18615
rect 15853 18581 15887 18615
rect 15887 18581 15896 18615
rect 15844 18572 15896 18581
rect 17132 18572 17184 18624
rect 17684 18572 17736 18624
rect 19800 18572 19852 18624
rect 20076 18572 20128 18624
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 6736 18411 6788 18420
rect 6736 18377 6745 18411
rect 6745 18377 6779 18411
rect 6779 18377 6788 18411
rect 6736 18368 6788 18377
rect 9220 18368 9272 18420
rect 6920 18300 6972 18352
rect 14280 18368 14332 18420
rect 16028 18411 16080 18420
rect 16028 18377 16037 18411
rect 16037 18377 16071 18411
rect 16071 18377 16080 18411
rect 16028 18368 16080 18377
rect 6644 18232 6696 18284
rect 2596 18096 2648 18148
rect 4896 18096 4948 18148
rect 3148 18028 3200 18080
rect 5448 18028 5500 18080
rect 7472 18071 7524 18080
rect 7472 18037 7481 18071
rect 7481 18037 7515 18071
rect 7515 18037 7524 18071
rect 7472 18028 7524 18037
rect 8116 18207 8168 18216
rect 8116 18173 8125 18207
rect 8125 18173 8159 18207
rect 8159 18173 8168 18207
rect 8116 18164 8168 18173
rect 8024 18096 8076 18148
rect 11152 18300 11204 18352
rect 12256 18300 12308 18352
rect 13820 18300 13872 18352
rect 18788 18368 18840 18420
rect 19708 18411 19760 18420
rect 19708 18377 19717 18411
rect 19717 18377 19751 18411
rect 19751 18377 19760 18411
rect 19708 18368 19760 18377
rect 9680 18232 9732 18284
rect 9864 18232 9916 18284
rect 10140 18275 10192 18284
rect 10140 18241 10158 18275
rect 10158 18241 10192 18275
rect 10140 18232 10192 18241
rect 10324 18232 10376 18284
rect 11336 18232 11388 18284
rect 11888 18232 11940 18284
rect 12624 18164 12676 18216
rect 14188 18232 14240 18284
rect 15844 18232 15896 18284
rect 18696 18300 18748 18352
rect 20628 18300 20680 18352
rect 16028 18164 16080 18216
rect 16488 18164 16540 18216
rect 18144 18164 18196 18216
rect 11704 18096 11756 18148
rect 10692 18071 10744 18080
rect 10692 18037 10701 18071
rect 10701 18037 10735 18071
rect 10735 18037 10744 18071
rect 10692 18028 10744 18037
rect 13544 18028 13596 18080
rect 16304 18096 16356 18148
rect 17684 18096 17736 18148
rect 17040 18028 17092 18080
rect 18052 18071 18104 18080
rect 18052 18037 18061 18071
rect 18061 18037 18095 18071
rect 18095 18037 18104 18071
rect 18052 18028 18104 18037
rect 21456 18028 21508 18080
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 9772 17824 9824 17876
rect 7104 17688 7156 17740
rect 7380 17688 7432 17740
rect 7656 17620 7708 17672
rect 9128 17620 9180 17672
rect 11704 17688 11756 17740
rect 4068 17552 4120 17604
rect 6736 17484 6788 17536
rect 10968 17484 11020 17536
rect 11152 17527 11204 17536
rect 11152 17493 11161 17527
rect 11161 17493 11195 17527
rect 11195 17493 11204 17527
rect 11152 17484 11204 17493
rect 11244 17484 11296 17536
rect 11888 17552 11940 17604
rect 16028 17824 16080 17876
rect 18144 17824 18196 17876
rect 19616 17799 19668 17808
rect 19616 17765 19625 17799
rect 19625 17765 19659 17799
rect 19659 17765 19668 17799
rect 19616 17756 19668 17765
rect 16488 17620 16540 17672
rect 19524 17620 19576 17672
rect 20628 17620 20680 17672
rect 18052 17552 18104 17604
rect 18604 17552 18656 17604
rect 15108 17484 15160 17536
rect 18788 17527 18840 17536
rect 18788 17493 18797 17527
rect 18797 17493 18831 17527
rect 18831 17493 18840 17527
rect 18788 17484 18840 17493
rect 21456 17552 21508 17604
rect 21548 17484 21600 17536
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 4252 17280 4304 17332
rect 4896 17323 4948 17332
rect 4896 17289 4905 17323
rect 4905 17289 4939 17323
rect 4939 17289 4948 17323
rect 4896 17280 4948 17289
rect 7656 17323 7708 17332
rect 7656 17289 7665 17323
rect 7665 17289 7699 17323
rect 7699 17289 7708 17323
rect 7656 17280 7708 17289
rect 8208 17280 8260 17332
rect 10048 17280 10100 17332
rect 10876 17280 10928 17332
rect 18972 17280 19024 17332
rect 6000 17212 6052 17264
rect 5540 17076 5592 17128
rect 9864 17144 9916 17196
rect 12348 17212 12400 17264
rect 12900 17144 12952 17196
rect 19708 17212 19760 17264
rect 14832 17187 14884 17196
rect 14832 17153 14850 17187
rect 14850 17153 14884 17187
rect 14832 17144 14884 17153
rect 8668 17008 8720 17060
rect 9128 17008 9180 17060
rect 12716 17008 12768 17060
rect 6644 16940 6696 16992
rect 10508 16940 10560 16992
rect 10692 16983 10744 16992
rect 10692 16949 10701 16983
rect 10701 16949 10735 16983
rect 10735 16949 10744 16983
rect 10692 16940 10744 16949
rect 11244 16940 11296 16992
rect 12348 16940 12400 16992
rect 13452 16983 13504 16992
rect 13452 16949 13461 16983
rect 13461 16949 13495 16983
rect 13495 16949 13504 16983
rect 13452 16940 13504 16949
rect 15752 17076 15804 17128
rect 18788 17144 18840 17196
rect 19984 17187 20036 17196
rect 19984 17153 20002 17187
rect 20002 17153 20036 17187
rect 19984 17144 20036 17153
rect 20168 17144 20220 17196
rect 20536 17144 20588 17196
rect 16028 16940 16080 16992
rect 18604 17008 18656 17060
rect 18696 16940 18748 16992
rect 18972 16940 19024 16992
rect 21180 16940 21232 16992
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 8668 16736 8720 16788
rect 11704 16736 11756 16788
rect 12992 16736 13044 16788
rect 13452 16736 13504 16788
rect 19524 16736 19576 16788
rect 9128 16532 9180 16584
rect 10692 16575 10744 16584
rect 10692 16541 10701 16575
rect 10701 16541 10735 16575
rect 10735 16541 10744 16575
rect 10692 16532 10744 16541
rect 12256 16600 12308 16652
rect 5540 16464 5592 16516
rect 4160 16396 4212 16448
rect 5908 16396 5960 16448
rect 7564 16464 7616 16516
rect 9956 16464 10008 16516
rect 12072 16532 12124 16584
rect 13268 16532 13320 16584
rect 12716 16464 12768 16516
rect 9588 16396 9640 16448
rect 10600 16396 10652 16448
rect 11244 16396 11296 16448
rect 12072 16439 12124 16448
rect 12072 16405 12081 16439
rect 12081 16405 12115 16439
rect 12115 16405 12124 16439
rect 12072 16396 12124 16405
rect 13268 16396 13320 16448
rect 15752 16575 15804 16584
rect 15752 16541 15761 16575
rect 15761 16541 15795 16575
rect 15795 16541 15804 16575
rect 15752 16532 15804 16541
rect 16028 16575 16080 16584
rect 16028 16541 16062 16575
rect 16062 16541 16080 16575
rect 16028 16532 16080 16541
rect 13452 16464 13504 16516
rect 15936 16464 15988 16516
rect 18328 16532 18380 16584
rect 20812 16532 20864 16584
rect 18236 16464 18288 16516
rect 18972 16464 19024 16516
rect 14740 16396 14792 16448
rect 18696 16396 18748 16448
rect 19708 16464 19760 16516
rect 19984 16464 20036 16516
rect 19156 16396 19208 16448
rect 20076 16396 20128 16448
rect 20168 16396 20220 16448
rect 21088 16439 21140 16448
rect 21088 16405 21097 16439
rect 21097 16405 21131 16439
rect 21131 16405 21140 16439
rect 21088 16396 21140 16405
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 4160 16235 4212 16244
rect 4160 16201 4169 16235
rect 4169 16201 4203 16235
rect 4203 16201 4212 16235
rect 4160 16192 4212 16201
rect 5356 16192 5408 16244
rect 7472 16192 7524 16244
rect 4620 15988 4672 16040
rect 4528 15895 4580 15904
rect 4528 15861 4537 15895
rect 4537 15861 4571 15895
rect 4571 15861 4580 15895
rect 4528 15852 4580 15861
rect 4804 15895 4856 15904
rect 4804 15861 4813 15895
rect 4813 15861 4847 15895
rect 4847 15861 4856 15895
rect 4804 15852 4856 15861
rect 7656 16056 7708 16108
rect 7748 16056 7800 16108
rect 12808 16192 12860 16244
rect 6920 15988 6972 16040
rect 7380 15988 7432 16040
rect 9128 15988 9180 16040
rect 17040 16124 17092 16176
rect 17132 16124 17184 16176
rect 20444 16192 20496 16244
rect 20904 16235 20956 16244
rect 20904 16201 20913 16235
rect 20913 16201 20947 16235
rect 20947 16201 20956 16235
rect 20904 16192 20956 16201
rect 10508 16056 10560 16108
rect 12256 16056 12308 16108
rect 14280 16056 14332 16108
rect 20720 16099 20772 16108
rect 10692 15988 10744 16040
rect 13268 16031 13320 16040
rect 5816 15895 5868 15904
rect 5816 15861 5825 15895
rect 5825 15861 5859 15895
rect 5859 15861 5868 15895
rect 5816 15852 5868 15861
rect 7104 15895 7156 15904
rect 7104 15861 7113 15895
rect 7113 15861 7147 15895
rect 7147 15861 7156 15895
rect 7104 15852 7156 15861
rect 7472 15852 7524 15904
rect 9404 15852 9456 15904
rect 13268 15997 13277 16031
rect 13277 15997 13311 16031
rect 13311 15997 13320 16031
rect 13268 15988 13320 15997
rect 15476 15920 15528 15972
rect 11060 15852 11112 15904
rect 12164 15852 12216 15904
rect 14648 15852 14700 15904
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15200 15852 15252 15861
rect 15752 15852 15804 15904
rect 18512 16031 18564 16040
rect 18512 15997 18521 16031
rect 18521 15997 18555 16031
rect 18555 15997 18564 16031
rect 18512 15988 18564 15997
rect 20720 16065 20729 16099
rect 20729 16065 20763 16099
rect 20763 16065 20772 16099
rect 20720 16056 20772 16065
rect 20996 15988 21048 16040
rect 20076 15852 20128 15904
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 21272 15852 21324 15861
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 6920 15580 6972 15632
rect 5908 15487 5960 15496
rect 5908 15453 5917 15487
rect 5917 15453 5951 15487
rect 5951 15453 5960 15487
rect 5908 15444 5960 15453
rect 7104 15512 7156 15564
rect 11152 15648 11204 15700
rect 11704 15648 11756 15700
rect 14372 15648 14424 15700
rect 7932 15580 7984 15632
rect 10140 15580 10192 15632
rect 10324 15444 10376 15496
rect 6092 15376 6144 15428
rect 4620 15351 4672 15360
rect 4620 15317 4629 15351
rect 4629 15317 4663 15351
rect 4663 15317 4672 15351
rect 4620 15308 4672 15317
rect 7564 15376 7616 15428
rect 9588 15376 9640 15428
rect 7288 15351 7340 15360
rect 7288 15317 7297 15351
rect 7297 15317 7331 15351
rect 7331 15317 7340 15351
rect 7288 15308 7340 15317
rect 7656 15351 7708 15360
rect 7656 15317 7665 15351
rect 7665 15317 7699 15351
rect 7699 15317 7708 15351
rect 7656 15308 7708 15317
rect 9128 15351 9180 15360
rect 9128 15317 9137 15351
rect 9137 15317 9171 15351
rect 9171 15317 9180 15351
rect 9128 15308 9180 15317
rect 11060 15308 11112 15360
rect 13268 15444 13320 15496
rect 16396 15444 16448 15496
rect 18512 15444 18564 15496
rect 21272 15444 21324 15496
rect 15200 15376 15252 15428
rect 15292 15419 15344 15428
rect 15292 15385 15310 15419
rect 15310 15385 15344 15419
rect 15292 15376 15344 15385
rect 15476 15376 15528 15428
rect 21088 15419 21140 15428
rect 21088 15385 21106 15419
rect 21106 15385 21140 15419
rect 21088 15376 21140 15385
rect 11704 15308 11756 15360
rect 13728 15351 13780 15360
rect 13728 15317 13737 15351
rect 13737 15317 13771 15351
rect 13771 15317 13780 15351
rect 13728 15308 13780 15317
rect 14280 15308 14332 15360
rect 15108 15308 15160 15360
rect 18052 15308 18104 15360
rect 18512 15308 18564 15360
rect 18696 15308 18748 15360
rect 19708 15351 19760 15360
rect 19708 15317 19717 15351
rect 19717 15317 19751 15351
rect 19751 15317 19760 15351
rect 19708 15308 19760 15317
rect 19892 15308 19944 15360
rect 20260 15308 20312 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 4528 15104 4580 15156
rect 6828 15147 6880 15156
rect 6828 15113 6837 15147
rect 6837 15113 6871 15147
rect 6871 15113 6880 15147
rect 6828 15104 6880 15113
rect 8024 15104 8076 15156
rect 12072 15104 12124 15156
rect 12348 15104 12400 15156
rect 15292 15104 15344 15156
rect 6184 15036 6236 15088
rect 6736 15036 6788 15088
rect 4804 14968 4856 15020
rect 7564 14968 7616 15020
rect 9404 14968 9456 15020
rect 20076 15036 20128 15088
rect 12900 14968 12952 15020
rect 13636 14968 13688 15020
rect 16396 14968 16448 15020
rect 17316 14968 17368 15020
rect 6736 14900 6788 14952
rect 8024 14900 8076 14952
rect 9128 14900 9180 14952
rect 19708 14943 19760 14952
rect 9680 14832 9732 14884
rect 5080 14764 5132 14816
rect 5356 14764 5408 14816
rect 19708 14909 19717 14943
rect 19717 14909 19751 14943
rect 19751 14909 19760 14943
rect 19708 14900 19760 14909
rect 11060 14832 11112 14884
rect 11152 14807 11204 14816
rect 11152 14773 11161 14807
rect 11161 14773 11195 14807
rect 11195 14773 11204 14807
rect 11152 14764 11204 14773
rect 12256 14764 12308 14816
rect 13728 14764 13780 14816
rect 15200 14764 15252 14816
rect 18052 14764 18104 14816
rect 21548 14832 21600 14884
rect 21088 14807 21140 14816
rect 21088 14773 21097 14807
rect 21097 14773 21131 14807
rect 21131 14773 21140 14807
rect 21088 14764 21140 14773
rect 22192 14764 22244 14816
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 3332 14603 3384 14612
rect 3332 14569 3341 14603
rect 3341 14569 3375 14603
rect 3375 14569 3384 14603
rect 3332 14560 3384 14569
rect 4528 14560 4580 14612
rect 6184 14603 6236 14612
rect 6184 14569 6193 14603
rect 6193 14569 6227 14603
rect 6227 14569 6236 14603
rect 6184 14560 6236 14569
rect 7840 14560 7892 14612
rect 9864 14560 9916 14612
rect 11704 14560 11756 14612
rect 13268 14560 13320 14612
rect 4804 14424 4856 14476
rect 4436 14356 4488 14408
rect 5448 14356 5500 14408
rect 9772 14356 9824 14408
rect 7104 14288 7156 14340
rect 10324 14331 10376 14340
rect 10324 14297 10342 14331
rect 10342 14297 10376 14331
rect 14556 14424 14608 14476
rect 11060 14356 11112 14408
rect 10324 14288 10376 14297
rect 3884 14220 3936 14272
rect 4712 14263 4764 14272
rect 4712 14229 4721 14263
rect 4721 14229 4755 14263
rect 4755 14229 4764 14263
rect 4712 14220 4764 14229
rect 5816 14220 5868 14272
rect 6920 14220 6972 14272
rect 7288 14263 7340 14272
rect 7288 14229 7297 14263
rect 7297 14229 7331 14263
rect 7331 14229 7340 14263
rect 9220 14263 9272 14272
rect 7288 14220 7340 14229
rect 9220 14229 9229 14263
rect 9229 14229 9263 14263
rect 9263 14229 9272 14263
rect 9220 14220 9272 14229
rect 11060 14220 11112 14272
rect 13452 14220 13504 14272
rect 13728 14220 13780 14272
rect 14924 14288 14976 14340
rect 19524 14424 19576 14476
rect 20076 14424 20128 14476
rect 16396 14356 16448 14408
rect 19708 14399 19760 14408
rect 19708 14365 19717 14399
rect 19717 14365 19751 14399
rect 19751 14365 19760 14399
rect 19708 14356 19760 14365
rect 21272 14356 21324 14408
rect 20168 14288 20220 14340
rect 21088 14331 21140 14340
rect 21088 14297 21106 14331
rect 21106 14297 21140 14331
rect 21088 14288 21140 14297
rect 17592 14220 17644 14272
rect 19340 14263 19392 14272
rect 19340 14229 19349 14263
rect 19349 14229 19383 14263
rect 19383 14229 19392 14263
rect 19340 14220 19392 14229
rect 19892 14220 19944 14272
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 3884 14016 3936 14068
rect 4436 14016 4488 14068
rect 5448 14016 5500 14068
rect 9680 14016 9732 14068
rect 7104 13948 7156 14000
rect 10140 13948 10192 14000
rect 10324 13991 10376 14000
rect 10324 13957 10342 13991
rect 10342 13957 10376 13991
rect 13176 14016 13228 14068
rect 13636 14016 13688 14068
rect 19340 14016 19392 14068
rect 10324 13948 10376 13957
rect 15292 13948 15344 14000
rect 17592 13948 17644 14000
rect 6092 13880 6144 13932
rect 6736 13880 6788 13932
rect 9956 13880 10008 13932
rect 12532 13880 12584 13932
rect 8300 13676 8352 13728
rect 8392 13676 8444 13728
rect 8668 13676 8720 13728
rect 11060 13812 11112 13864
rect 15660 13855 15712 13864
rect 15660 13821 15669 13855
rect 15669 13821 15703 13855
rect 15703 13821 15712 13855
rect 15660 13812 15712 13821
rect 19064 13948 19116 14000
rect 21640 14016 21692 14068
rect 19432 13923 19484 13932
rect 19432 13889 19450 13923
rect 19450 13889 19484 13923
rect 19432 13880 19484 13889
rect 20168 13880 20220 13932
rect 21272 13880 21324 13932
rect 13544 13676 13596 13728
rect 15016 13676 15068 13728
rect 16856 13676 16908 13728
rect 17040 13676 17092 13728
rect 17776 13676 17828 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 6736 13472 6788 13524
rect 8668 13472 8720 13524
rect 6092 13404 6144 13456
rect 10232 13472 10284 13524
rect 11704 13472 11756 13524
rect 11888 13472 11940 13524
rect 12256 13472 12308 13524
rect 13544 13472 13596 13524
rect 5264 13379 5316 13388
rect 5264 13345 5273 13379
rect 5273 13345 5307 13379
rect 5307 13345 5316 13379
rect 5264 13336 5316 13345
rect 8300 13336 8352 13388
rect 5448 13268 5500 13320
rect 6460 13268 6512 13320
rect 6552 13268 6604 13320
rect 9128 13268 9180 13320
rect 12072 13311 12124 13320
rect 12072 13277 12081 13311
rect 12081 13277 12115 13311
rect 12115 13277 12124 13311
rect 13728 13311 13780 13320
rect 12072 13268 12124 13277
rect 13728 13277 13737 13311
rect 13737 13277 13771 13311
rect 13771 13277 13780 13311
rect 13728 13268 13780 13277
rect 17868 13472 17920 13524
rect 20628 13472 20680 13524
rect 18236 13447 18288 13456
rect 18236 13413 18245 13447
rect 18245 13413 18279 13447
rect 18279 13413 18288 13447
rect 18236 13404 18288 13413
rect 18788 13447 18840 13456
rect 18788 13413 18797 13447
rect 18797 13413 18831 13447
rect 18831 13413 18840 13447
rect 18788 13404 18840 13413
rect 17500 13336 17552 13388
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 15660 13268 15712 13320
rect 16304 13268 16356 13320
rect 21272 13336 21324 13388
rect 20904 13311 20956 13320
rect 20904 13277 20913 13311
rect 20913 13277 20947 13311
rect 20947 13277 20956 13311
rect 20904 13268 20956 13277
rect 5724 13175 5776 13184
rect 5724 13141 5733 13175
rect 5733 13141 5767 13175
rect 5767 13141 5776 13175
rect 5724 13132 5776 13141
rect 8392 13200 8444 13252
rect 13084 13200 13136 13252
rect 15016 13200 15068 13252
rect 6828 13132 6880 13184
rect 7840 13132 7892 13184
rect 9680 13132 9732 13184
rect 10416 13175 10468 13184
rect 10416 13141 10425 13175
rect 10425 13141 10459 13175
rect 10459 13141 10468 13175
rect 10416 13132 10468 13141
rect 14004 13132 14056 13184
rect 14280 13132 14332 13184
rect 16028 13200 16080 13252
rect 17040 13200 17092 13252
rect 15844 13132 15896 13184
rect 22008 13132 22060 13184
rect 22560 13132 22612 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 5724 12928 5776 12980
rect 7840 12971 7892 12980
rect 7840 12937 7849 12971
rect 7849 12937 7883 12971
rect 7883 12937 7892 12971
rect 7840 12928 7892 12937
rect 8484 12928 8536 12980
rect 17224 12928 17276 12980
rect 5356 12903 5408 12912
rect 5356 12869 5365 12903
rect 5365 12869 5399 12903
rect 5399 12869 5408 12903
rect 5356 12860 5408 12869
rect 8300 12860 8352 12912
rect 5724 12792 5776 12844
rect 5908 12792 5960 12844
rect 6552 12792 6604 12844
rect 6736 12835 6788 12844
rect 6736 12801 6770 12835
rect 6770 12801 6788 12835
rect 6736 12792 6788 12801
rect 8116 12835 8168 12844
rect 8116 12801 8125 12835
rect 8125 12801 8159 12835
rect 8159 12801 8168 12835
rect 8116 12792 8168 12801
rect 9312 12792 9364 12844
rect 11060 12860 11112 12912
rect 12072 12860 12124 12912
rect 12716 12860 12768 12912
rect 4988 12724 5040 12776
rect 11980 12792 12032 12844
rect 12256 12792 12308 12844
rect 14004 12835 14056 12844
rect 15476 12860 15528 12912
rect 14004 12801 14022 12835
rect 14022 12801 14056 12835
rect 14004 12792 14056 12801
rect 14648 12792 14700 12844
rect 14832 12792 14884 12844
rect 18696 12860 18748 12912
rect 20168 12860 20220 12912
rect 21640 12860 21692 12912
rect 16120 12792 16172 12844
rect 19708 12792 19760 12844
rect 21272 12792 21324 12844
rect 10876 12724 10928 12776
rect 18052 12767 18104 12776
rect 18052 12733 18061 12767
rect 18061 12733 18095 12767
rect 18095 12733 18104 12767
rect 18052 12724 18104 12733
rect 16028 12656 16080 12708
rect 8484 12588 8536 12640
rect 9036 12588 9088 12640
rect 9220 12588 9272 12640
rect 11152 12631 11204 12640
rect 11152 12597 11161 12631
rect 11161 12597 11195 12631
rect 11195 12597 11204 12631
rect 11152 12588 11204 12597
rect 11796 12588 11848 12640
rect 14280 12588 14332 12640
rect 14556 12631 14608 12640
rect 14556 12597 14565 12631
rect 14565 12597 14599 12631
rect 14599 12597 14608 12631
rect 14556 12588 14608 12597
rect 18696 12588 18748 12640
rect 19892 12588 19944 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 6736 12248 6788 12300
rect 10416 12384 10468 12436
rect 12716 12384 12768 12436
rect 5632 12180 5684 12232
rect 6000 12180 6052 12232
rect 6552 12180 6604 12232
rect 7932 12180 7984 12232
rect 9036 12316 9088 12368
rect 13820 12316 13872 12368
rect 16028 12384 16080 12436
rect 16120 12316 16172 12368
rect 9036 12180 9088 12232
rect 10600 12248 10652 12300
rect 11152 12248 11204 12300
rect 15476 12291 15528 12300
rect 9864 12180 9916 12232
rect 10876 12180 10928 12232
rect 11060 12180 11112 12232
rect 15476 12257 15485 12291
rect 15485 12257 15519 12291
rect 15519 12257 15528 12291
rect 15476 12248 15528 12257
rect 17592 12248 17644 12300
rect 17776 12248 17828 12300
rect 17040 12180 17092 12232
rect 18052 12180 18104 12232
rect 19064 12180 19116 12232
rect 20444 12384 20496 12436
rect 21272 12180 21324 12232
rect 4988 12087 5040 12096
rect 4988 12053 4997 12087
rect 4997 12053 5031 12087
rect 5031 12053 5040 12087
rect 4988 12044 5040 12053
rect 5908 12087 5960 12096
rect 5908 12053 5917 12087
rect 5917 12053 5951 12087
rect 5951 12053 5960 12087
rect 5908 12044 5960 12053
rect 6000 12044 6052 12096
rect 6736 12044 6788 12096
rect 7196 12044 7248 12096
rect 7656 12044 7708 12096
rect 9680 12112 9732 12164
rect 10324 12112 10376 12164
rect 9128 12044 9180 12096
rect 9496 12044 9548 12096
rect 12992 12112 13044 12164
rect 15568 12112 15620 12164
rect 11152 12044 11204 12096
rect 12532 12044 12584 12096
rect 12716 12044 12768 12096
rect 14924 12044 14976 12096
rect 16948 12112 17000 12164
rect 17592 12112 17644 12164
rect 17960 12112 18012 12164
rect 18144 12112 18196 12164
rect 21548 12112 21600 12164
rect 22100 12112 22152 12164
rect 18788 12044 18840 12096
rect 19064 12044 19116 12096
rect 19524 12044 19576 12096
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 6460 11840 6512 11892
rect 6828 11840 6880 11892
rect 7012 11883 7064 11892
rect 7012 11849 7021 11883
rect 7021 11849 7055 11883
rect 7055 11849 7064 11883
rect 7012 11840 7064 11849
rect 8024 11840 8076 11892
rect 8208 11840 8260 11892
rect 9128 11840 9180 11892
rect 12900 11883 12952 11892
rect 5172 11704 5224 11756
rect 6092 11704 6144 11756
rect 6828 11704 6880 11756
rect 7104 11704 7156 11756
rect 7840 11704 7892 11756
rect 8392 11636 8444 11688
rect 8576 11679 8628 11688
rect 8576 11645 8585 11679
rect 8585 11645 8619 11679
rect 8619 11645 8628 11679
rect 8576 11636 8628 11645
rect 11060 11772 11112 11824
rect 11244 11772 11296 11824
rect 12900 11849 12909 11883
rect 12909 11849 12943 11883
rect 12943 11849 12952 11883
rect 12900 11840 12952 11849
rect 14372 11883 14424 11892
rect 14372 11849 14381 11883
rect 14381 11849 14415 11883
rect 14415 11849 14424 11883
rect 14372 11840 14424 11849
rect 14740 11840 14792 11892
rect 14924 11840 14976 11892
rect 15476 11840 15528 11892
rect 16120 11840 16172 11892
rect 16948 11840 17000 11892
rect 17868 11840 17920 11892
rect 15752 11772 15804 11824
rect 17040 11772 17092 11824
rect 11796 11704 11848 11756
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 14372 11704 14424 11756
rect 15200 11704 15252 11756
rect 17224 11747 17276 11756
rect 17224 11713 17233 11747
rect 17233 11713 17267 11747
rect 17267 11713 17276 11747
rect 17224 11704 17276 11713
rect 18052 11772 18104 11824
rect 18696 11840 18748 11892
rect 20904 11840 20956 11892
rect 21272 11772 21324 11824
rect 5172 11500 5224 11552
rect 7104 11500 7156 11552
rect 8484 11500 8536 11552
rect 8760 11500 8812 11552
rect 9312 11500 9364 11552
rect 10876 11500 10928 11552
rect 11336 11636 11388 11688
rect 12164 11636 12216 11688
rect 14832 11679 14884 11688
rect 11060 11568 11112 11620
rect 11152 11500 11204 11552
rect 11704 11500 11756 11552
rect 12624 11568 12676 11620
rect 14832 11645 14841 11679
rect 14841 11645 14875 11679
rect 14875 11645 14884 11679
rect 14832 11636 14884 11645
rect 16948 11679 17000 11688
rect 13636 11500 13688 11552
rect 16948 11645 16957 11679
rect 16957 11645 16991 11679
rect 16991 11645 17000 11679
rect 16948 11636 17000 11645
rect 19892 11636 19944 11688
rect 18144 11500 18196 11552
rect 19708 11500 19760 11552
rect 21548 11568 21600 11620
rect 21088 11500 21140 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 6092 11296 6144 11348
rect 7288 11296 7340 11348
rect 7564 11339 7616 11348
rect 7564 11305 7573 11339
rect 7573 11305 7607 11339
rect 7607 11305 7616 11339
rect 7564 11296 7616 11305
rect 7840 11339 7892 11348
rect 7840 11305 7849 11339
rect 7849 11305 7883 11339
rect 7883 11305 7892 11339
rect 7840 11296 7892 11305
rect 6000 11160 6052 11212
rect 9496 11271 9548 11280
rect 9496 11237 9505 11271
rect 9505 11237 9539 11271
rect 9539 11237 9548 11271
rect 9496 11228 9548 11237
rect 10876 11228 10928 11280
rect 12164 11271 12216 11280
rect 8208 11160 8260 11212
rect 7104 11135 7156 11144
rect 5908 11024 5960 11076
rect 7104 11101 7113 11135
rect 7113 11101 7147 11135
rect 7147 11101 7156 11135
rect 7104 11092 7156 11101
rect 11060 11160 11112 11212
rect 11428 11160 11480 11212
rect 12164 11237 12173 11271
rect 12173 11237 12207 11271
rect 12207 11237 12216 11271
rect 12164 11228 12216 11237
rect 13452 11296 13504 11348
rect 14556 11296 14608 11348
rect 14832 11296 14884 11348
rect 15200 11339 15252 11348
rect 15200 11305 15209 11339
rect 15209 11305 15243 11339
rect 15243 11305 15252 11339
rect 15200 11296 15252 11305
rect 17040 11339 17092 11348
rect 17040 11305 17049 11339
rect 17049 11305 17083 11339
rect 17083 11305 17092 11339
rect 17040 11296 17092 11305
rect 18420 11296 18472 11348
rect 12624 11228 12676 11280
rect 12532 11160 12584 11212
rect 11152 11092 11204 11144
rect 11244 11092 11296 11144
rect 12624 11092 12676 11144
rect 6460 10956 6512 11008
rect 7012 10956 7064 11008
rect 7196 10999 7248 11008
rect 7196 10965 7205 10999
rect 7205 10965 7239 10999
rect 7239 10965 7248 10999
rect 7196 10956 7248 10965
rect 8392 10956 8444 11008
rect 10416 10956 10468 11008
rect 11336 11024 11388 11076
rect 12164 10956 12216 11008
rect 12440 10999 12492 11008
rect 12440 10965 12449 10999
rect 12449 10965 12483 10999
rect 12483 10965 12492 10999
rect 12900 11228 12952 11280
rect 13084 11203 13136 11212
rect 13084 11169 13093 11203
rect 13093 11169 13127 11203
rect 13127 11169 13136 11203
rect 13084 11160 13136 11169
rect 15752 11203 15804 11212
rect 15752 11169 15761 11203
rect 15761 11169 15795 11203
rect 15795 11169 15804 11203
rect 15752 11160 15804 11169
rect 16948 11228 17000 11280
rect 14096 11092 14148 11144
rect 14556 11092 14608 11144
rect 14648 11092 14700 11144
rect 14832 11092 14884 11144
rect 16120 11092 16172 11144
rect 16212 11092 16264 11144
rect 18696 11160 18748 11212
rect 18420 11135 18472 11144
rect 18420 11101 18429 11135
rect 18429 11101 18463 11135
rect 18463 11101 18472 11135
rect 18420 11092 18472 11101
rect 19800 11203 19852 11212
rect 19800 11169 19809 11203
rect 19809 11169 19843 11203
rect 19843 11169 19852 11203
rect 19800 11160 19852 11169
rect 20352 11160 20404 11212
rect 12900 11067 12952 11076
rect 12900 11033 12909 11067
rect 12909 11033 12943 11067
rect 12943 11033 12952 11067
rect 15660 11067 15712 11076
rect 12900 11024 12952 11033
rect 15660 11033 15669 11067
rect 15669 11033 15703 11067
rect 15703 11033 15712 11067
rect 15660 11024 15712 11033
rect 17040 11024 17092 11076
rect 12440 10956 12492 10965
rect 13084 10956 13136 11008
rect 14188 10956 14240 11008
rect 14648 10956 14700 11008
rect 15016 10956 15068 11008
rect 17316 10999 17368 11008
rect 17316 10965 17325 10999
rect 17325 10965 17359 10999
rect 17359 10965 17368 10999
rect 17316 10956 17368 10965
rect 17960 11024 18012 11076
rect 19708 11067 19760 11076
rect 19708 11033 19717 11067
rect 19717 11033 19751 11067
rect 19751 11033 19760 11067
rect 19708 11024 19760 11033
rect 20168 11024 20220 11076
rect 20536 11024 20588 11076
rect 21272 11067 21324 11076
rect 21272 11033 21281 11067
rect 21281 11033 21315 11067
rect 21315 11033 21324 11067
rect 21272 11024 21324 11033
rect 22008 11024 22060 11076
rect 22376 11024 22428 11076
rect 18880 10956 18932 11008
rect 19340 10956 19392 11008
rect 19800 10956 19852 11008
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 5724 10752 5776 10804
rect 5908 10752 5960 10804
rect 6736 10752 6788 10804
rect 7196 10752 7248 10804
rect 7932 10795 7984 10804
rect 7932 10761 7941 10795
rect 7941 10761 7975 10795
rect 7975 10761 7984 10795
rect 7932 10752 7984 10761
rect 8576 10752 8628 10804
rect 10140 10795 10192 10804
rect 10140 10761 10149 10795
rect 10149 10761 10183 10795
rect 10183 10761 10192 10795
rect 10140 10752 10192 10761
rect 10416 10752 10468 10804
rect 10692 10752 10744 10804
rect 12164 10752 12216 10804
rect 12440 10752 12492 10804
rect 13636 10752 13688 10804
rect 13912 10752 13964 10804
rect 14372 10795 14424 10804
rect 14372 10761 14381 10795
rect 14381 10761 14415 10795
rect 14415 10761 14424 10795
rect 14372 10752 14424 10761
rect 8392 10684 8444 10736
rect 11612 10684 11664 10736
rect 17316 10752 17368 10804
rect 17684 10752 17736 10804
rect 18144 10752 18196 10804
rect 18420 10752 18472 10804
rect 19340 10752 19392 10804
rect 20628 10752 20680 10804
rect 6736 10659 6788 10668
rect 6736 10625 6745 10659
rect 6745 10625 6779 10659
rect 6779 10625 6788 10659
rect 6736 10616 6788 10625
rect 7932 10616 7984 10668
rect 8852 10616 8904 10668
rect 6552 10548 6604 10600
rect 6920 10548 6972 10600
rect 7472 10480 7524 10532
rect 5724 10412 5776 10464
rect 7104 10455 7156 10464
rect 7104 10421 7113 10455
rect 7113 10421 7147 10455
rect 7147 10421 7156 10455
rect 7104 10412 7156 10421
rect 9128 10548 9180 10600
rect 9864 10616 9916 10668
rect 11152 10616 11204 10668
rect 11244 10616 11296 10668
rect 13728 10659 13780 10668
rect 13728 10625 13737 10659
rect 13737 10625 13771 10659
rect 13771 10625 13780 10659
rect 13728 10616 13780 10625
rect 13820 10616 13872 10668
rect 10324 10548 10376 10600
rect 10600 10591 10652 10600
rect 10600 10557 10609 10591
rect 10609 10557 10643 10591
rect 10643 10557 10652 10591
rect 10600 10548 10652 10557
rect 11060 10548 11112 10600
rect 12256 10548 12308 10600
rect 13636 10591 13688 10600
rect 10968 10480 11020 10532
rect 13636 10557 13645 10591
rect 13645 10557 13679 10591
rect 13679 10557 13688 10591
rect 13636 10548 13688 10557
rect 14924 10591 14976 10600
rect 14924 10557 14933 10591
rect 14933 10557 14967 10591
rect 14967 10557 14976 10591
rect 14924 10548 14976 10557
rect 15200 10616 15252 10668
rect 16304 10684 16356 10736
rect 19800 10684 19852 10736
rect 16672 10659 16724 10668
rect 16672 10625 16681 10659
rect 16681 10625 16715 10659
rect 16715 10625 16724 10659
rect 16672 10616 16724 10625
rect 17500 10616 17552 10668
rect 17960 10616 18012 10668
rect 18696 10616 18748 10668
rect 20076 10616 20128 10668
rect 20628 10659 20680 10668
rect 20628 10625 20637 10659
rect 20637 10625 20671 10659
rect 20671 10625 20680 10659
rect 20628 10616 20680 10625
rect 22008 10616 22060 10668
rect 22284 10616 22336 10668
rect 16212 10548 16264 10600
rect 16580 10548 16632 10600
rect 18144 10591 18196 10600
rect 18144 10557 18153 10591
rect 18153 10557 18187 10591
rect 18187 10557 18196 10591
rect 18144 10548 18196 10557
rect 18972 10548 19024 10600
rect 19524 10480 19576 10532
rect 12440 10412 12492 10464
rect 12808 10412 12860 10464
rect 13820 10412 13872 10464
rect 13912 10412 13964 10464
rect 14188 10412 14240 10464
rect 15752 10412 15804 10464
rect 17500 10412 17552 10464
rect 18052 10412 18104 10464
rect 18972 10412 19024 10464
rect 20444 10548 20496 10600
rect 20352 10480 20404 10532
rect 20168 10412 20220 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 7288 10208 7340 10260
rect 8208 10208 8260 10260
rect 12808 10208 12860 10260
rect 14556 10251 14608 10260
rect 14556 10217 14565 10251
rect 14565 10217 14599 10251
rect 14599 10217 14608 10251
rect 14556 10208 14608 10217
rect 17408 10208 17460 10260
rect 21180 10251 21232 10260
rect 21180 10217 21189 10251
rect 21189 10217 21223 10251
rect 21223 10217 21232 10251
rect 21180 10208 21232 10217
rect 5540 10140 5592 10192
rect 7104 10140 7156 10192
rect 16672 10140 16724 10192
rect 5264 10072 5316 10124
rect 5448 10115 5500 10124
rect 5448 10081 5457 10115
rect 5457 10081 5491 10115
rect 5491 10081 5500 10115
rect 5448 10072 5500 10081
rect 5908 10072 5960 10124
rect 4988 10004 5040 10056
rect 6828 10072 6880 10124
rect 9220 10115 9272 10124
rect 9220 10081 9229 10115
rect 9229 10081 9263 10115
rect 9263 10081 9272 10115
rect 9220 10072 9272 10081
rect 9312 10072 9364 10124
rect 11152 10115 11204 10124
rect 11152 10081 11161 10115
rect 11161 10081 11195 10115
rect 11195 10081 11204 10115
rect 11152 10072 11204 10081
rect 11612 10115 11664 10124
rect 11612 10081 11621 10115
rect 11621 10081 11655 10115
rect 11655 10081 11664 10115
rect 11612 10072 11664 10081
rect 13544 10072 13596 10124
rect 13728 10072 13780 10124
rect 15936 10072 15988 10124
rect 7288 10004 7340 10056
rect 7932 10004 7984 10056
rect 10508 10004 10560 10056
rect 12256 10004 12308 10056
rect 15200 10004 15252 10056
rect 17960 10072 18012 10124
rect 18328 10115 18380 10124
rect 18328 10081 18337 10115
rect 18337 10081 18371 10115
rect 18371 10081 18380 10115
rect 18328 10072 18380 10081
rect 18696 10115 18748 10124
rect 18696 10081 18705 10115
rect 18705 10081 18739 10115
rect 18739 10081 18748 10115
rect 18696 10072 18748 10081
rect 16948 10047 17000 10056
rect 5356 9936 5408 9988
rect 8392 9936 8444 9988
rect 9956 9936 10008 9988
rect 16948 10013 16957 10047
rect 16957 10013 16991 10047
rect 16991 10013 17000 10047
rect 16948 10004 17000 10013
rect 19524 10047 19576 10056
rect 19524 10013 19533 10047
rect 19533 10013 19567 10047
rect 19567 10013 19576 10047
rect 20260 10047 20312 10056
rect 19524 10004 19576 10013
rect 20260 10013 20269 10047
rect 20269 10013 20303 10047
rect 20303 10013 20312 10047
rect 20260 10004 20312 10013
rect 15936 9936 15988 9988
rect 16580 9936 16632 9988
rect 17408 9936 17460 9988
rect 5724 9911 5776 9920
rect 5724 9877 5733 9911
rect 5733 9877 5767 9911
rect 5767 9877 5776 9911
rect 5724 9868 5776 9877
rect 6000 9868 6052 9920
rect 7012 9868 7064 9920
rect 7472 9868 7524 9920
rect 7932 9868 7984 9920
rect 8576 9911 8628 9920
rect 8576 9877 8585 9911
rect 8585 9877 8619 9911
rect 8619 9877 8628 9911
rect 8576 9868 8628 9877
rect 9680 9868 9732 9920
rect 9864 9911 9916 9920
rect 9864 9877 9873 9911
rect 9873 9877 9907 9911
rect 9907 9877 9916 9911
rect 9864 9868 9916 9877
rect 10416 9911 10468 9920
rect 10416 9877 10425 9911
rect 10425 9877 10459 9911
rect 10459 9877 10468 9911
rect 10416 9868 10468 9877
rect 10508 9911 10560 9920
rect 10508 9877 10517 9911
rect 10517 9877 10551 9911
rect 10551 9877 10560 9911
rect 10508 9868 10560 9877
rect 11244 9868 11296 9920
rect 12624 9911 12676 9920
rect 12624 9877 12633 9911
rect 12633 9877 12667 9911
rect 12667 9877 12676 9911
rect 12624 9868 12676 9877
rect 13360 9868 13412 9920
rect 13728 9868 13780 9920
rect 15108 9911 15160 9920
rect 15108 9877 15117 9911
rect 15117 9877 15151 9911
rect 15151 9877 15160 9911
rect 15108 9868 15160 9877
rect 15200 9868 15252 9920
rect 17040 9868 17092 9920
rect 18052 9911 18104 9920
rect 18052 9877 18061 9911
rect 18061 9877 18095 9911
rect 18095 9877 18104 9911
rect 18052 9868 18104 9877
rect 18144 9911 18196 9920
rect 18144 9877 18153 9911
rect 18153 9877 18187 9911
rect 18187 9877 18196 9911
rect 19892 9936 19944 9988
rect 18144 9868 18196 9877
rect 20812 9868 20864 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 6000 9664 6052 9716
rect 9864 9664 9916 9716
rect 10508 9664 10560 9716
rect 11244 9664 11296 9716
rect 6644 9639 6696 9648
rect 6644 9605 6653 9639
rect 6653 9605 6687 9639
rect 6687 9605 6696 9639
rect 6644 9596 6696 9605
rect 8668 9639 8720 9648
rect 5724 9528 5776 9580
rect 7748 9571 7800 9580
rect 7748 9537 7757 9571
rect 7757 9537 7791 9571
rect 7791 9537 7800 9571
rect 7748 9528 7800 9537
rect 8668 9605 8677 9639
rect 8677 9605 8711 9639
rect 8711 9605 8720 9639
rect 8668 9596 8720 9605
rect 11704 9596 11756 9648
rect 15108 9664 15160 9716
rect 17040 9707 17092 9716
rect 17040 9673 17049 9707
rect 17049 9673 17083 9707
rect 17083 9673 17092 9707
rect 17040 9664 17092 9673
rect 18144 9664 18196 9716
rect 20536 9664 20588 9716
rect 8760 9571 8812 9580
rect 8760 9537 8769 9571
rect 8769 9537 8803 9571
rect 8803 9537 8812 9571
rect 8760 9528 8812 9537
rect 9312 9528 9364 9580
rect 4804 9460 4856 9512
rect 5724 9392 5776 9444
rect 5908 9460 5960 9512
rect 6276 9460 6328 9512
rect 6644 9460 6696 9512
rect 7564 9503 7616 9512
rect 7564 9469 7573 9503
rect 7573 9469 7607 9503
rect 7607 9469 7616 9503
rect 7564 9460 7616 9469
rect 9220 9460 9272 9512
rect 11980 9528 12032 9580
rect 8116 9435 8168 9444
rect 8116 9401 8125 9435
rect 8125 9401 8159 9435
rect 8159 9401 8168 9435
rect 8116 9392 8168 9401
rect 12164 9435 12216 9444
rect 7196 9324 7248 9376
rect 7288 9324 7340 9376
rect 11888 9324 11940 9376
rect 12164 9401 12173 9435
rect 12173 9401 12207 9435
rect 12207 9401 12216 9435
rect 12164 9392 12216 9401
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 13268 9528 13320 9580
rect 14924 9528 14976 9580
rect 15660 9571 15712 9580
rect 15660 9537 15669 9571
rect 15669 9537 15703 9571
rect 15703 9537 15712 9571
rect 15660 9528 15712 9537
rect 13728 9460 13780 9512
rect 14556 9460 14608 9512
rect 15108 9460 15160 9512
rect 15752 9460 15804 9512
rect 16396 9460 16448 9512
rect 16580 9460 16632 9512
rect 17132 9528 17184 9580
rect 17684 9528 17736 9580
rect 20260 9596 20312 9648
rect 19892 9571 19944 9580
rect 19892 9537 19901 9571
rect 19901 9537 19935 9571
rect 19935 9537 19944 9571
rect 19892 9528 19944 9537
rect 16948 9503 17000 9512
rect 16948 9469 16957 9503
rect 16957 9469 16991 9503
rect 16991 9469 17000 9503
rect 16948 9460 17000 9469
rect 17132 9392 17184 9444
rect 18144 9460 18196 9512
rect 18880 9503 18932 9512
rect 18880 9469 18889 9503
rect 18889 9469 18923 9503
rect 18923 9469 18932 9503
rect 18880 9460 18932 9469
rect 19340 9460 19392 9512
rect 14556 9324 14608 9376
rect 16304 9324 16356 9376
rect 16948 9324 17000 9376
rect 17040 9324 17092 9376
rect 18052 9392 18104 9444
rect 20352 9392 20404 9444
rect 19340 9324 19392 9376
rect 19984 9324 20036 9376
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 6552 9120 6604 9172
rect 6644 9120 6696 9172
rect 9588 9120 9640 9172
rect 9956 9163 10008 9172
rect 9956 9129 9965 9163
rect 9965 9129 9999 9163
rect 9999 9129 10008 9163
rect 9956 9120 10008 9129
rect 10416 9120 10468 9172
rect 11980 9120 12032 9172
rect 14004 9120 14056 9172
rect 14188 9163 14240 9172
rect 14188 9129 14197 9163
rect 14197 9129 14231 9163
rect 14231 9129 14240 9163
rect 14188 9120 14240 9129
rect 14924 9120 14976 9172
rect 15108 9163 15160 9172
rect 15108 9129 15117 9163
rect 15117 9129 15151 9163
rect 15151 9129 15160 9163
rect 15108 9120 15160 9129
rect 15752 9120 15804 9172
rect 16212 9120 16264 9172
rect 17684 9163 17736 9172
rect 17684 9129 17693 9163
rect 17693 9129 17727 9163
rect 17727 9129 17736 9163
rect 17684 9120 17736 9129
rect 6000 8984 6052 9036
rect 7840 9052 7892 9104
rect 10876 9052 10928 9104
rect 15660 9052 15712 9104
rect 17960 9052 18012 9104
rect 9404 9027 9456 9036
rect 9404 8993 9413 9027
rect 9413 8993 9447 9027
rect 9447 8993 9456 9027
rect 9404 8984 9456 8993
rect 9680 8984 9732 9036
rect 12532 9027 12584 9036
rect 12532 8993 12541 9027
rect 12541 8993 12575 9027
rect 12575 8993 12584 9027
rect 12532 8984 12584 8993
rect 13268 9027 13320 9036
rect 13268 8993 13277 9027
rect 13277 8993 13311 9027
rect 13311 8993 13320 9027
rect 13268 8984 13320 8993
rect 16580 8984 16632 9036
rect 18788 9120 18840 9172
rect 19432 9120 19484 9172
rect 19708 9120 19760 9172
rect 18236 9052 18288 9104
rect 18512 8984 18564 9036
rect 18972 8984 19024 9036
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 7196 8959 7248 8968
rect 7196 8925 7205 8959
rect 7205 8925 7239 8959
rect 7239 8925 7248 8959
rect 7196 8916 7248 8925
rect 10140 8916 10192 8968
rect 11152 8916 11204 8968
rect 14004 8916 14056 8968
rect 18052 8959 18104 8968
rect 18052 8925 18061 8959
rect 18061 8925 18095 8959
rect 18095 8925 18104 8959
rect 18052 8916 18104 8925
rect 18236 8916 18288 8968
rect 4712 8848 4764 8900
rect 5816 8848 5868 8900
rect 6276 8823 6328 8832
rect 6276 8789 6285 8823
rect 6285 8789 6319 8823
rect 6319 8789 6328 8823
rect 6276 8780 6328 8789
rect 7288 8780 7340 8832
rect 7656 8780 7708 8832
rect 7840 8823 7892 8832
rect 7840 8789 7849 8823
rect 7849 8789 7883 8823
rect 7883 8789 7892 8823
rect 7840 8780 7892 8789
rect 8668 8780 8720 8832
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 11152 8780 11204 8832
rect 16396 8848 16448 8900
rect 13820 8780 13872 8832
rect 15200 8780 15252 8832
rect 15384 8780 15436 8832
rect 15568 8780 15620 8832
rect 16304 8780 16356 8832
rect 16948 8780 17000 8832
rect 20812 8916 20864 8968
rect 19524 8891 19576 8900
rect 19524 8857 19533 8891
rect 19533 8857 19567 8891
rect 19567 8857 19576 8891
rect 19524 8848 19576 8857
rect 18880 8780 18932 8832
rect 22284 8848 22336 8900
rect 20904 8823 20956 8832
rect 20904 8789 20913 8823
rect 20913 8789 20947 8823
rect 20947 8789 20956 8823
rect 20904 8780 20956 8789
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 9404 8576 9456 8628
rect 10140 8619 10192 8628
rect 10140 8585 10149 8619
rect 10149 8585 10183 8619
rect 10183 8585 10192 8619
rect 10140 8576 10192 8585
rect 12808 8576 12860 8628
rect 13544 8576 13596 8628
rect 15200 8619 15252 8628
rect 15200 8585 15209 8619
rect 15209 8585 15243 8619
rect 15243 8585 15252 8619
rect 15200 8576 15252 8585
rect 15936 8576 15988 8628
rect 16948 8619 17000 8628
rect 16948 8585 16957 8619
rect 16957 8585 16991 8619
rect 16991 8585 17000 8619
rect 16948 8576 17000 8585
rect 17040 8619 17092 8628
rect 17040 8585 17049 8619
rect 17049 8585 17083 8619
rect 17083 8585 17092 8619
rect 17040 8576 17092 8585
rect 4988 8508 5040 8560
rect 5356 8415 5408 8424
rect 5356 8381 5365 8415
rect 5365 8381 5399 8415
rect 5399 8381 5408 8415
rect 5356 8372 5408 8381
rect 5540 8372 5592 8424
rect 8668 8508 8720 8560
rect 9772 8508 9824 8560
rect 11980 8440 12032 8492
rect 9680 8372 9732 8424
rect 10600 8415 10652 8424
rect 5264 8304 5316 8356
rect 6920 8279 6972 8288
rect 6920 8245 6929 8279
rect 6929 8245 6963 8279
rect 6963 8245 6972 8279
rect 6920 8236 6972 8245
rect 9128 8279 9180 8288
rect 9128 8245 9137 8279
rect 9137 8245 9171 8279
rect 9171 8245 9180 8279
rect 9128 8236 9180 8245
rect 10600 8381 10609 8415
rect 10609 8381 10643 8415
rect 10643 8381 10652 8415
rect 10600 8372 10652 8381
rect 10876 8372 10928 8424
rect 10968 8372 11020 8424
rect 13268 8372 13320 8424
rect 11888 8304 11940 8356
rect 11244 8236 11296 8288
rect 12532 8236 12584 8288
rect 14280 8508 14332 8560
rect 16028 8551 16080 8560
rect 16028 8517 16037 8551
rect 16037 8517 16071 8551
rect 16071 8517 16080 8551
rect 16028 8508 16080 8517
rect 16856 8508 16908 8560
rect 17960 8576 18012 8628
rect 18144 8619 18196 8628
rect 18144 8585 18153 8619
rect 18153 8585 18187 8619
rect 18187 8585 18196 8619
rect 18144 8576 18196 8585
rect 18420 8576 18472 8628
rect 19616 8576 19668 8628
rect 20260 8619 20312 8628
rect 20260 8585 20269 8619
rect 20269 8585 20303 8619
rect 20303 8585 20312 8619
rect 20260 8576 20312 8585
rect 20904 8576 20956 8628
rect 20996 8576 21048 8628
rect 21180 8576 21232 8628
rect 18236 8508 18288 8560
rect 18696 8508 18748 8560
rect 18328 8440 18380 8492
rect 18788 8440 18840 8492
rect 19524 8483 19576 8492
rect 19524 8449 19533 8483
rect 19533 8449 19567 8483
rect 19567 8449 19576 8483
rect 19524 8440 19576 8449
rect 19984 8440 20036 8492
rect 20904 8440 20956 8492
rect 13912 8372 13964 8424
rect 15200 8372 15252 8424
rect 17224 8372 17276 8424
rect 13544 8236 13596 8288
rect 14832 8347 14884 8356
rect 14832 8313 14841 8347
rect 14841 8313 14875 8347
rect 14875 8313 14884 8347
rect 14832 8304 14884 8313
rect 15384 8304 15436 8356
rect 14280 8236 14332 8288
rect 18512 8304 18564 8356
rect 21180 8372 21232 8424
rect 21456 8372 21508 8424
rect 18328 8236 18380 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 6736 8032 6788 8084
rect 7748 8032 7800 8084
rect 10140 8075 10192 8084
rect 10140 8041 10149 8075
rect 10149 8041 10183 8075
rect 10183 8041 10192 8075
rect 10140 8032 10192 8041
rect 10324 8032 10376 8084
rect 12624 8032 12676 8084
rect 13728 8075 13780 8084
rect 13728 8041 13737 8075
rect 13737 8041 13771 8075
rect 13771 8041 13780 8075
rect 13728 8032 13780 8041
rect 14556 8032 14608 8084
rect 15384 8032 15436 8084
rect 16856 8032 16908 8084
rect 21364 8032 21416 8084
rect 8668 7964 8720 8016
rect 10416 7964 10468 8016
rect 10968 7964 11020 8016
rect 5264 7939 5316 7948
rect 5264 7905 5273 7939
rect 5273 7905 5307 7939
rect 5307 7905 5316 7939
rect 5264 7896 5316 7905
rect 6000 7896 6052 7948
rect 6920 7896 6972 7948
rect 9128 7896 9180 7948
rect 9588 7939 9640 7948
rect 9588 7905 9597 7939
rect 9597 7905 9631 7939
rect 9631 7905 9640 7939
rect 9588 7896 9640 7905
rect 12440 7964 12492 8016
rect 16212 7964 16264 8016
rect 17960 7964 18012 8016
rect 22192 7964 22244 8016
rect 12164 7896 12216 7948
rect 12716 7896 12768 7948
rect 14372 7896 14424 7948
rect 5540 7828 5592 7880
rect 12532 7871 12584 7880
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 17500 7896 17552 7948
rect 18696 7939 18748 7948
rect 18696 7905 18705 7939
rect 18705 7905 18739 7939
rect 18739 7905 18748 7939
rect 18696 7896 18748 7905
rect 20720 7896 20772 7948
rect 4252 7692 4304 7744
rect 5448 7692 5500 7744
rect 10692 7760 10744 7812
rect 12440 7803 12492 7812
rect 12440 7769 12449 7803
rect 12449 7769 12483 7803
rect 12483 7769 12492 7803
rect 12440 7760 12492 7769
rect 12624 7760 12676 7812
rect 14924 7828 14976 7880
rect 20168 7871 20220 7880
rect 20168 7837 20177 7871
rect 20177 7837 20211 7871
rect 20211 7837 20220 7871
rect 20168 7828 20220 7837
rect 20812 7828 20864 7880
rect 13728 7760 13780 7812
rect 17132 7760 17184 7812
rect 19524 7803 19576 7812
rect 19524 7769 19533 7803
rect 19533 7769 19567 7803
rect 19567 7769 19576 7803
rect 19524 7760 19576 7769
rect 5908 7692 5960 7744
rect 8668 7692 8720 7744
rect 11980 7692 12032 7744
rect 12164 7692 12216 7744
rect 13084 7692 13136 7744
rect 13452 7692 13504 7744
rect 14556 7692 14608 7744
rect 15936 7692 15988 7744
rect 16304 7735 16356 7744
rect 16304 7701 16313 7735
rect 16313 7701 16347 7735
rect 16347 7701 16356 7735
rect 16304 7692 16356 7701
rect 16396 7692 16448 7744
rect 17776 7735 17828 7744
rect 17776 7701 17785 7735
rect 17785 7701 17819 7735
rect 17819 7701 17828 7735
rect 17776 7692 17828 7701
rect 18420 7735 18472 7744
rect 18420 7701 18429 7735
rect 18429 7701 18463 7735
rect 18463 7701 18472 7735
rect 18420 7692 18472 7701
rect 18512 7735 18564 7744
rect 18512 7701 18521 7735
rect 18521 7701 18555 7735
rect 18555 7701 18564 7735
rect 18512 7692 18564 7701
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 5356 7488 5408 7540
rect 5908 7488 5960 7540
rect 9588 7488 9640 7540
rect 10600 7488 10652 7540
rect 11060 7488 11112 7540
rect 11980 7531 12032 7540
rect 11980 7497 11989 7531
rect 11989 7497 12023 7531
rect 12023 7497 12032 7531
rect 11980 7488 12032 7497
rect 9404 7463 9456 7472
rect 4988 7327 5040 7336
rect 4988 7293 4997 7327
rect 4997 7293 5031 7327
rect 5031 7293 5040 7327
rect 4988 7284 5040 7293
rect 5172 7327 5224 7336
rect 5172 7293 5181 7327
rect 5181 7293 5215 7327
rect 5215 7293 5224 7327
rect 5172 7284 5224 7293
rect 5724 7284 5776 7336
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 6644 7327 6696 7336
rect 6644 7293 6653 7327
rect 6653 7293 6687 7327
rect 6687 7293 6696 7327
rect 6644 7284 6696 7293
rect 9404 7429 9413 7463
rect 9413 7429 9447 7463
rect 9447 7429 9456 7463
rect 10140 7463 10192 7472
rect 9404 7420 9456 7429
rect 10140 7429 10149 7463
rect 10149 7429 10183 7463
rect 10183 7429 10192 7463
rect 10140 7420 10192 7429
rect 8208 7352 8260 7404
rect 10692 7420 10744 7472
rect 12164 7420 12216 7472
rect 13636 7488 13688 7540
rect 14556 7531 14608 7540
rect 14556 7497 14565 7531
rect 14565 7497 14599 7531
rect 14599 7497 14608 7531
rect 14556 7488 14608 7497
rect 14924 7531 14976 7540
rect 14924 7497 14933 7531
rect 14933 7497 14967 7531
rect 14967 7497 14976 7531
rect 14924 7488 14976 7497
rect 16304 7488 16356 7540
rect 17776 7488 17828 7540
rect 18420 7488 18472 7540
rect 2596 7216 2648 7268
rect 13084 7352 13136 7404
rect 14280 7420 14332 7472
rect 16396 7420 16448 7472
rect 21088 7420 21140 7472
rect 14832 7352 14884 7404
rect 15568 7395 15620 7404
rect 15568 7361 15577 7395
rect 15577 7361 15611 7395
rect 15611 7361 15620 7395
rect 15568 7352 15620 7361
rect 12072 7327 12124 7336
rect 12072 7293 12081 7327
rect 12081 7293 12115 7327
rect 12115 7293 12124 7327
rect 12072 7284 12124 7293
rect 13820 7284 13872 7336
rect 14464 7284 14516 7336
rect 15844 7327 15896 7336
rect 15844 7293 15853 7327
rect 15853 7293 15887 7327
rect 15887 7293 15896 7327
rect 15844 7284 15896 7293
rect 17316 7352 17368 7404
rect 17776 7352 17828 7404
rect 18328 7352 18380 7404
rect 16948 7327 17000 7336
rect 16948 7293 16957 7327
rect 16957 7293 16991 7327
rect 16991 7293 17000 7327
rect 16948 7284 17000 7293
rect 17960 7327 18012 7336
rect 17960 7293 17969 7327
rect 17969 7293 18003 7327
rect 18003 7293 18012 7327
rect 17960 7284 18012 7293
rect 18144 7327 18196 7336
rect 18144 7293 18153 7327
rect 18153 7293 18187 7327
rect 18187 7293 18196 7327
rect 18144 7284 18196 7293
rect 4160 7148 4212 7200
rect 5172 7148 5224 7200
rect 5908 7191 5960 7200
rect 5908 7157 5917 7191
rect 5917 7157 5951 7191
rect 5951 7157 5960 7191
rect 5908 7148 5960 7157
rect 6644 7148 6696 7200
rect 12072 7148 12124 7200
rect 19524 7352 19576 7404
rect 20720 7395 20772 7404
rect 20720 7361 20729 7395
rect 20729 7361 20763 7395
rect 20763 7361 20772 7395
rect 20720 7352 20772 7361
rect 19616 7327 19668 7336
rect 19616 7293 19625 7327
rect 19625 7293 19659 7327
rect 19659 7293 19668 7327
rect 19616 7284 19668 7293
rect 20812 7284 20864 7336
rect 13820 7148 13872 7200
rect 15660 7148 15712 7200
rect 16212 7148 16264 7200
rect 18328 7148 18380 7200
rect 18604 7148 18656 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 8392 6944 8444 6996
rect 15568 6987 15620 6996
rect 6644 6876 6696 6928
rect 10876 6876 10928 6928
rect 13084 6876 13136 6928
rect 15568 6953 15577 6987
rect 15577 6953 15611 6987
rect 15611 6953 15620 6987
rect 15568 6944 15620 6953
rect 16948 6944 17000 6996
rect 18512 6944 18564 6996
rect 15936 6876 15988 6928
rect 6736 6808 6788 6860
rect 9864 6808 9916 6860
rect 10692 6851 10744 6860
rect 10692 6817 10701 6851
rect 10701 6817 10735 6851
rect 10735 6817 10744 6851
rect 10692 6808 10744 6817
rect 11152 6851 11204 6860
rect 11152 6817 11161 6851
rect 11161 6817 11195 6851
rect 11195 6817 11204 6851
rect 11152 6808 11204 6817
rect 11980 6851 12032 6860
rect 11980 6817 11989 6851
rect 11989 6817 12023 6851
rect 12023 6817 12032 6851
rect 11980 6808 12032 6817
rect 12532 6808 12584 6860
rect 13544 6808 13596 6860
rect 15016 6808 15068 6860
rect 16120 6808 16172 6860
rect 17500 6876 17552 6928
rect 17684 6808 17736 6860
rect 17960 6851 18012 6860
rect 17960 6817 17969 6851
rect 17969 6817 18003 6851
rect 18003 6817 18012 6851
rect 17960 6808 18012 6817
rect 19340 6851 19392 6860
rect 19340 6817 19349 6851
rect 19349 6817 19383 6851
rect 19383 6817 19392 6851
rect 19340 6808 19392 6817
rect 19524 6808 19576 6860
rect 20444 6851 20496 6860
rect 20444 6817 20453 6851
rect 20453 6817 20487 6851
rect 20487 6817 20496 6851
rect 20444 6808 20496 6817
rect 10600 6740 10652 6792
rect 11244 6740 11296 6792
rect 12716 6672 12768 6724
rect 9680 6604 9732 6656
rect 10600 6604 10652 6656
rect 10876 6604 10928 6656
rect 12532 6647 12584 6656
rect 12532 6613 12541 6647
rect 12541 6613 12575 6647
rect 12575 6613 12584 6647
rect 18052 6740 18104 6792
rect 20076 6740 20128 6792
rect 20812 6783 20864 6792
rect 20812 6749 20821 6783
rect 20821 6749 20855 6783
rect 20855 6749 20864 6783
rect 20812 6740 20864 6749
rect 14280 6672 14332 6724
rect 14924 6672 14976 6724
rect 15384 6672 15436 6724
rect 16304 6672 16356 6724
rect 12532 6604 12584 6613
rect 13820 6604 13872 6656
rect 15016 6604 15068 6656
rect 16948 6647 17000 6656
rect 16948 6613 16957 6647
rect 16957 6613 16991 6647
rect 16991 6613 17000 6647
rect 16948 6604 17000 6613
rect 18604 6604 18656 6656
rect 20352 6604 20404 6656
rect 22560 6604 22612 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 10508 6443 10560 6452
rect 10508 6409 10517 6443
rect 10517 6409 10551 6443
rect 10551 6409 10560 6443
rect 10508 6400 10560 6409
rect 11152 6400 11204 6452
rect 12440 6400 12492 6452
rect 12624 6400 12676 6452
rect 13176 6443 13228 6452
rect 13176 6409 13185 6443
rect 13185 6409 13219 6443
rect 13219 6409 13228 6443
rect 13176 6400 13228 6409
rect 17500 6400 17552 6452
rect 18788 6400 18840 6452
rect 18972 6400 19024 6452
rect 19248 6400 19300 6452
rect 12716 6332 12768 6384
rect 12900 6332 12952 6384
rect 13544 6332 13596 6384
rect 14924 6332 14976 6384
rect 9128 6307 9180 6316
rect 9128 6273 9137 6307
rect 9137 6273 9171 6307
rect 9171 6273 9180 6307
rect 9128 6264 9180 6273
rect 10140 6307 10192 6316
rect 10140 6273 10149 6307
rect 10149 6273 10183 6307
rect 10183 6273 10192 6307
rect 10140 6264 10192 6273
rect 12164 6307 12216 6316
rect 12164 6273 12173 6307
rect 12173 6273 12207 6307
rect 12207 6273 12216 6307
rect 12164 6264 12216 6273
rect 12992 6264 13044 6316
rect 9772 6196 9824 6248
rect 10232 6196 10284 6248
rect 10692 6196 10744 6248
rect 12900 6196 12952 6248
rect 13728 6264 13780 6316
rect 14464 6307 14516 6316
rect 14464 6273 14473 6307
rect 14473 6273 14507 6307
rect 14507 6273 14516 6307
rect 14464 6264 14516 6273
rect 15936 6264 15988 6316
rect 16120 6264 16172 6316
rect 17040 6264 17092 6316
rect 18236 6332 18288 6384
rect 19524 6332 19576 6384
rect 19984 6375 20036 6384
rect 19984 6341 19993 6375
rect 19993 6341 20027 6375
rect 20027 6341 20036 6375
rect 19984 6332 20036 6341
rect 20904 6332 20956 6384
rect 19708 6307 19760 6316
rect 14740 6239 14792 6248
rect 14740 6205 14749 6239
rect 14749 6205 14783 6239
rect 14783 6205 14792 6239
rect 14740 6196 14792 6205
rect 15292 6239 15344 6248
rect 15292 6205 15301 6239
rect 15301 6205 15335 6239
rect 15335 6205 15344 6239
rect 15292 6196 15344 6205
rect 16948 6196 17000 6248
rect 17224 6196 17276 6248
rect 17592 6196 17644 6248
rect 17776 6196 17828 6248
rect 19708 6273 19717 6307
rect 19717 6273 19751 6307
rect 19751 6273 19760 6307
rect 19708 6264 19760 6273
rect 19616 6196 19668 6248
rect 19892 6196 19944 6248
rect 21088 6239 21140 6248
rect 21088 6205 21097 6239
rect 21097 6205 21131 6239
rect 21131 6205 21140 6239
rect 21088 6196 21140 6205
rect 21180 6239 21232 6248
rect 21180 6205 21189 6239
rect 21189 6205 21223 6239
rect 21223 6205 21232 6239
rect 21180 6196 21232 6205
rect 21548 6196 21600 6248
rect 9496 6128 9548 6180
rect 11152 6128 11204 6180
rect 16764 6128 16816 6180
rect 8024 6060 8076 6112
rect 11888 6060 11940 6112
rect 13452 6060 13504 6112
rect 15016 6060 15068 6112
rect 17960 6128 18012 6180
rect 18052 6128 18104 6180
rect 17132 6060 17184 6112
rect 18144 6060 18196 6112
rect 19340 6060 19392 6112
rect 19892 6060 19944 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 3516 5856 3568 5908
rect 8300 5856 8352 5908
rect 9220 5856 9272 5908
rect 10140 5856 10192 5908
rect 10416 5899 10468 5908
rect 10416 5865 10425 5899
rect 10425 5865 10459 5899
rect 10459 5865 10468 5899
rect 10416 5856 10468 5865
rect 11888 5899 11940 5908
rect 11888 5865 11897 5899
rect 11897 5865 11931 5899
rect 11931 5865 11940 5899
rect 11888 5856 11940 5865
rect 12900 5899 12952 5908
rect 12900 5865 12909 5899
rect 12909 5865 12943 5899
rect 12943 5865 12952 5899
rect 12900 5856 12952 5865
rect 8484 5788 8536 5840
rect 9496 5763 9548 5772
rect 9496 5729 9505 5763
rect 9505 5729 9539 5763
rect 9539 5729 9548 5763
rect 9496 5720 9548 5729
rect 9956 5788 10008 5840
rect 12348 5720 12400 5772
rect 9680 5695 9732 5704
rect 9680 5661 9689 5695
rect 9689 5661 9723 5695
rect 9723 5661 9732 5695
rect 9680 5652 9732 5661
rect 11152 5652 11204 5704
rect 12532 5652 12584 5704
rect 8300 5584 8352 5636
rect 9588 5559 9640 5568
rect 9588 5525 9597 5559
rect 9597 5525 9631 5559
rect 9631 5525 9640 5559
rect 9588 5516 9640 5525
rect 10968 5516 11020 5568
rect 11152 5559 11204 5568
rect 11152 5525 11161 5559
rect 11161 5525 11195 5559
rect 11195 5525 11204 5559
rect 13820 5856 13872 5908
rect 15200 5856 15252 5908
rect 15936 5899 15988 5908
rect 13728 5788 13780 5840
rect 15384 5788 15436 5840
rect 15936 5865 15945 5899
rect 15945 5865 15979 5899
rect 15979 5865 15988 5899
rect 15936 5856 15988 5865
rect 16948 5899 17000 5908
rect 16948 5865 16957 5899
rect 16957 5865 16991 5899
rect 16991 5865 17000 5899
rect 16948 5856 17000 5865
rect 17040 5856 17092 5908
rect 18144 5856 18196 5908
rect 13544 5763 13596 5772
rect 13544 5729 13553 5763
rect 13553 5729 13587 5763
rect 13587 5729 13596 5763
rect 13544 5720 13596 5729
rect 17316 5788 17368 5840
rect 17776 5788 17828 5840
rect 15660 5720 15712 5772
rect 16028 5720 16080 5772
rect 16212 5720 16264 5772
rect 17500 5763 17552 5772
rect 17500 5729 17509 5763
rect 17509 5729 17543 5763
rect 17543 5729 17552 5763
rect 17500 5720 17552 5729
rect 17592 5720 17644 5772
rect 18144 5720 18196 5772
rect 19064 5788 19116 5840
rect 19984 5788 20036 5840
rect 18420 5763 18472 5772
rect 18420 5729 18429 5763
rect 18429 5729 18463 5763
rect 18463 5729 18472 5763
rect 18420 5720 18472 5729
rect 19800 5720 19852 5772
rect 13176 5652 13228 5704
rect 13820 5652 13872 5704
rect 15200 5652 15252 5704
rect 17408 5695 17460 5704
rect 17408 5661 17417 5695
rect 17417 5661 17451 5695
rect 17451 5661 17460 5695
rect 17408 5652 17460 5661
rect 18512 5695 18564 5704
rect 18512 5661 18521 5695
rect 18521 5661 18555 5695
rect 18555 5661 18564 5695
rect 18512 5652 18564 5661
rect 18880 5652 18932 5704
rect 19892 5695 19944 5704
rect 19892 5661 19901 5695
rect 19901 5661 19935 5695
rect 19935 5661 19944 5695
rect 19892 5652 19944 5661
rect 20904 5652 20956 5704
rect 22284 5652 22336 5704
rect 16488 5584 16540 5636
rect 11152 5516 11204 5525
rect 15200 5516 15252 5568
rect 16120 5516 16172 5568
rect 16764 5516 16816 5568
rect 17040 5516 17092 5568
rect 17500 5516 17552 5568
rect 17684 5516 17736 5568
rect 18880 5559 18932 5568
rect 18880 5525 18889 5559
rect 18889 5525 18923 5559
rect 18923 5525 18932 5559
rect 18880 5516 18932 5525
rect 20260 5559 20312 5568
rect 20260 5525 20269 5559
rect 20269 5525 20303 5559
rect 20303 5525 20312 5559
rect 20260 5516 20312 5525
rect 20536 5559 20588 5568
rect 20536 5525 20545 5559
rect 20545 5525 20579 5559
rect 20579 5525 20588 5559
rect 20536 5516 20588 5525
rect 20904 5559 20956 5568
rect 20904 5525 20913 5559
rect 20913 5525 20947 5559
rect 20947 5525 20956 5559
rect 20904 5516 20956 5525
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 8116 5312 8168 5364
rect 8576 5312 8628 5364
rect 8760 5312 8812 5364
rect 5080 5244 5132 5296
rect 6828 5176 6880 5228
rect 8760 5219 8812 5228
rect 8760 5185 8769 5219
rect 8769 5185 8803 5219
rect 8803 5185 8812 5219
rect 8760 5176 8812 5185
rect 8944 5244 8996 5296
rect 9312 5244 9364 5296
rect 9588 5312 9640 5364
rect 9956 5355 10008 5364
rect 9956 5321 9965 5355
rect 9965 5321 9999 5355
rect 9999 5321 10008 5355
rect 9956 5312 10008 5321
rect 10140 5244 10192 5296
rect 7840 5108 7892 5160
rect 10048 5108 10100 5160
rect 10784 5312 10836 5364
rect 11152 5312 11204 5364
rect 13452 5355 13504 5364
rect 13452 5321 13461 5355
rect 13461 5321 13495 5355
rect 13495 5321 13504 5355
rect 13452 5312 13504 5321
rect 13912 5355 13964 5364
rect 13912 5321 13921 5355
rect 13921 5321 13955 5355
rect 13955 5321 13964 5355
rect 13912 5312 13964 5321
rect 14924 5355 14976 5364
rect 14924 5321 14933 5355
rect 14933 5321 14967 5355
rect 14967 5321 14976 5355
rect 14924 5312 14976 5321
rect 15200 5312 15252 5364
rect 15384 5312 15436 5364
rect 15844 5355 15896 5364
rect 15844 5321 15853 5355
rect 15853 5321 15887 5355
rect 15887 5321 15896 5355
rect 15844 5312 15896 5321
rect 16396 5312 16448 5364
rect 16764 5312 16816 5364
rect 17132 5244 17184 5296
rect 18880 5312 18932 5364
rect 13544 5219 13596 5228
rect 13544 5185 13553 5219
rect 13553 5185 13587 5219
rect 13587 5185 13596 5219
rect 13544 5176 13596 5185
rect 15016 5176 15068 5228
rect 12164 5151 12216 5160
rect 12164 5117 12173 5151
rect 12173 5117 12207 5151
rect 12207 5117 12216 5151
rect 12164 5108 12216 5117
rect 12808 5108 12860 5160
rect 12992 5108 13044 5160
rect 13360 5151 13412 5160
rect 13360 5117 13369 5151
rect 13369 5117 13403 5151
rect 13403 5117 13412 5151
rect 13360 5108 13412 5117
rect 14648 5151 14700 5160
rect 14648 5117 14657 5151
rect 14657 5117 14691 5151
rect 14691 5117 14700 5151
rect 14648 5108 14700 5117
rect 17408 5176 17460 5228
rect 17684 5219 17736 5228
rect 17684 5185 17693 5219
rect 17693 5185 17727 5219
rect 17727 5185 17736 5219
rect 17684 5176 17736 5185
rect 20536 5312 20588 5364
rect 20260 5244 20312 5296
rect 11152 5083 11204 5092
rect 11152 5049 11161 5083
rect 11161 5049 11195 5083
rect 11195 5049 11204 5083
rect 11152 5040 11204 5049
rect 14372 5040 14424 5092
rect 17224 5108 17276 5160
rect 17868 5151 17920 5160
rect 17868 5117 17877 5151
rect 17877 5117 17911 5151
rect 17911 5117 17920 5151
rect 17868 5108 17920 5117
rect 16764 5040 16816 5092
rect 18052 5040 18104 5092
rect 18880 5108 18932 5160
rect 19800 5151 19852 5160
rect 19800 5117 19809 5151
rect 19809 5117 19843 5151
rect 19843 5117 19852 5151
rect 19800 5108 19852 5117
rect 19984 5151 20036 5160
rect 19984 5117 19993 5151
rect 19993 5117 20027 5151
rect 20027 5117 20036 5151
rect 19984 5108 20036 5117
rect 21180 5176 21232 5228
rect 20444 5108 20496 5160
rect 20996 5151 21048 5160
rect 20996 5117 21005 5151
rect 21005 5117 21039 5151
rect 21039 5117 21048 5151
rect 20996 5108 21048 5117
rect 21640 5040 21692 5092
rect 2044 4972 2096 5024
rect 5080 4972 5132 5024
rect 8484 5015 8536 5024
rect 8484 4981 8493 5015
rect 8493 4981 8527 5015
rect 8527 4981 8536 5015
rect 8484 4972 8536 4981
rect 8944 4972 8996 5024
rect 13820 4972 13872 5024
rect 14464 4972 14516 5024
rect 15200 4972 15252 5024
rect 16120 4972 16172 5024
rect 17132 4972 17184 5024
rect 17316 5015 17368 5024
rect 17316 4981 17325 5015
rect 17325 4981 17359 5015
rect 17359 4981 17368 5015
rect 17316 4972 17368 4981
rect 20352 5015 20404 5024
rect 20352 4981 20361 5015
rect 20361 4981 20395 5015
rect 20395 4981 20404 5015
rect 20352 4972 20404 4981
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 8208 4768 8260 4820
rect 1400 4700 1452 4752
rect 9128 4768 9180 4820
rect 9772 4768 9824 4820
rect 13544 4768 13596 4820
rect 15292 4768 15344 4820
rect 17684 4768 17736 4820
rect 19616 4768 19668 4820
rect 20168 4811 20220 4820
rect 20168 4777 20177 4811
rect 20177 4777 20211 4811
rect 20211 4777 20220 4811
rect 20168 4768 20220 4777
rect 21272 4811 21324 4820
rect 21272 4777 21281 4811
rect 21281 4777 21315 4811
rect 21315 4777 21324 4811
rect 21272 4768 21324 4777
rect 13176 4700 13228 4752
rect 17960 4700 18012 4752
rect 21088 4700 21140 4752
rect 10048 4675 10100 4684
rect 7380 4564 7432 4616
rect 8852 4564 8904 4616
rect 10048 4641 10057 4675
rect 10057 4641 10091 4675
rect 10091 4641 10100 4675
rect 10048 4632 10100 4641
rect 10324 4632 10376 4684
rect 12256 4675 12308 4684
rect 12256 4641 12265 4675
rect 12265 4641 12299 4675
rect 12299 4641 12308 4675
rect 12256 4632 12308 4641
rect 13268 4675 13320 4684
rect 13268 4641 13277 4675
rect 13277 4641 13311 4675
rect 13311 4641 13320 4675
rect 13268 4632 13320 4641
rect 14740 4675 14792 4684
rect 14740 4641 14749 4675
rect 14749 4641 14783 4675
rect 14783 4641 14792 4675
rect 14740 4632 14792 4641
rect 14924 4632 14976 4684
rect 15108 4632 15160 4684
rect 15660 4675 15712 4684
rect 15660 4641 15669 4675
rect 15669 4641 15703 4675
rect 15703 4641 15712 4675
rect 15660 4632 15712 4641
rect 15844 4632 15896 4684
rect 18880 4632 18932 4684
rect 20260 4632 20312 4684
rect 20904 4632 20956 4684
rect 12992 4607 13044 4616
rect 12992 4573 13001 4607
rect 13001 4573 13035 4607
rect 13035 4573 13044 4607
rect 12992 4564 13044 4573
rect 17040 4564 17092 4616
rect 17960 4564 18012 4616
rect 9680 4496 9732 4548
rect 10048 4496 10100 4548
rect 11152 4496 11204 4548
rect 9128 4471 9180 4480
rect 9128 4437 9137 4471
rect 9137 4437 9171 4471
rect 9171 4437 9180 4471
rect 9128 4428 9180 4437
rect 10692 4428 10744 4480
rect 11888 4428 11940 4480
rect 12532 4428 12584 4480
rect 14188 4428 14240 4480
rect 14556 4471 14608 4480
rect 14556 4437 14565 4471
rect 14565 4437 14599 4471
rect 14599 4437 14608 4471
rect 15384 4496 15436 4548
rect 16028 4496 16080 4548
rect 17500 4496 17552 4548
rect 14556 4428 14608 4437
rect 15752 4428 15804 4480
rect 20536 4428 20588 4480
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 8852 4267 8904 4276
rect 8852 4233 8861 4267
rect 8861 4233 8895 4267
rect 8895 4233 8904 4267
rect 8852 4224 8904 4233
rect 9680 4267 9732 4276
rect 9680 4233 9689 4267
rect 9689 4233 9723 4267
rect 9723 4233 9732 4267
rect 9680 4224 9732 4233
rect 10324 4267 10376 4276
rect 10324 4233 10333 4267
rect 10333 4233 10367 4267
rect 10367 4233 10376 4267
rect 10324 4224 10376 4233
rect 12164 4224 12216 4276
rect 12532 4224 12584 4276
rect 13728 4224 13780 4276
rect 14188 4267 14240 4276
rect 14188 4233 14197 4267
rect 14197 4233 14231 4267
rect 14231 4233 14240 4267
rect 14188 4224 14240 4233
rect 16028 4224 16080 4276
rect 17776 4224 17828 4276
rect 3148 4088 3200 4140
rect 5908 4088 5960 4140
rect 10692 4020 10744 4072
rect 16488 4156 16540 4208
rect 17408 4156 17460 4208
rect 19616 4156 19668 4208
rect 12440 4088 12492 4140
rect 12716 4088 12768 4140
rect 13268 4088 13320 4140
rect 13452 4063 13504 4072
rect 13452 4029 13461 4063
rect 13461 4029 13495 4063
rect 13495 4029 13504 4063
rect 13452 4020 13504 4029
rect 14280 4088 14332 4140
rect 17316 4131 17368 4140
rect 14648 4020 14700 4072
rect 15108 4020 15160 4072
rect 17316 4097 17325 4131
rect 17325 4097 17359 4131
rect 17359 4097 17368 4131
rect 17316 4088 17368 4097
rect 20352 4088 20404 4140
rect 20536 4131 20588 4140
rect 20536 4097 20545 4131
rect 20545 4097 20579 4131
rect 20579 4097 20588 4131
rect 20536 4088 20588 4097
rect 21180 4131 21232 4140
rect 21180 4097 21189 4131
rect 21189 4097 21223 4131
rect 21223 4097 21232 4131
rect 21180 4088 21232 4097
rect 16304 4020 16356 4072
rect 16948 4020 17000 4072
rect 19064 4020 19116 4072
rect 19156 4020 19208 4072
rect 19984 4020 20036 4072
rect 940 3884 992 3936
rect 8668 3884 8720 3936
rect 10048 3927 10100 3936
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 11704 3884 11756 3936
rect 14556 3952 14608 4004
rect 12808 3884 12860 3936
rect 13636 3884 13688 3936
rect 16120 3927 16172 3936
rect 16120 3893 16129 3927
rect 16129 3893 16163 3927
rect 16163 3893 16172 3927
rect 16120 3884 16172 3893
rect 17868 3952 17920 4004
rect 19800 3952 19852 4004
rect 20352 3952 20404 4004
rect 18236 3884 18288 3936
rect 18788 3884 18840 3936
rect 19524 3884 19576 3936
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 4620 3680 4672 3732
rect 5908 3680 5960 3732
rect 10048 3680 10100 3732
rect 12808 3680 12860 3732
rect 14740 3680 14792 3732
rect 9220 3612 9272 3664
rect 11060 3612 11112 3664
rect 5632 3544 5684 3596
rect 10232 3587 10284 3596
rect 10232 3553 10241 3587
rect 10241 3553 10275 3587
rect 10275 3553 10284 3587
rect 10232 3544 10284 3553
rect 10692 3587 10744 3596
rect 10692 3553 10701 3587
rect 10701 3553 10735 3587
rect 10735 3553 10744 3587
rect 10692 3544 10744 3553
rect 10876 3544 10928 3596
rect 13820 3544 13872 3596
rect 15476 3612 15528 3664
rect 15108 3544 15160 3596
rect 16120 3544 16172 3596
rect 17224 3680 17276 3732
rect 19616 3723 19668 3732
rect 19616 3689 19625 3723
rect 19625 3689 19659 3723
rect 19659 3689 19668 3723
rect 19616 3680 19668 3689
rect 20812 3680 20864 3732
rect 20260 3612 20312 3664
rect 22100 3612 22152 3664
rect 10968 3519 11020 3528
rect 10968 3485 10977 3519
rect 10977 3485 11011 3519
rect 11011 3485 11020 3519
rect 10968 3476 11020 3485
rect 12072 3476 12124 3528
rect 12440 3476 12492 3528
rect 13360 3476 13412 3528
rect 11060 3408 11112 3460
rect 11152 3408 11204 3460
rect 11980 3408 12032 3460
rect 7012 3340 7064 3392
rect 13084 3340 13136 3392
rect 15384 3476 15436 3528
rect 15568 3476 15620 3528
rect 16488 3476 16540 3528
rect 17132 3476 17184 3528
rect 17960 3476 18012 3528
rect 22376 3544 22428 3596
rect 13544 3340 13596 3392
rect 14832 3340 14884 3392
rect 15292 3340 15344 3392
rect 15752 3340 15804 3392
rect 16304 3408 16356 3460
rect 20076 3408 20128 3460
rect 16396 3340 16448 3392
rect 18788 3340 18840 3392
rect 19340 3383 19392 3392
rect 19340 3349 19349 3383
rect 19349 3349 19383 3383
rect 19383 3349 19392 3383
rect 19340 3340 19392 3349
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 8484 3136 8536 3188
rect 9864 3179 9916 3188
rect 9864 3145 9873 3179
rect 9873 3145 9907 3179
rect 9907 3145 9916 3179
rect 9864 3136 9916 3145
rect 10140 3179 10192 3188
rect 10140 3145 10149 3179
rect 10149 3145 10183 3179
rect 10183 3145 10192 3179
rect 10140 3136 10192 3145
rect 10600 3179 10652 3188
rect 10600 3145 10609 3179
rect 10609 3145 10643 3179
rect 10643 3145 10652 3179
rect 10600 3136 10652 3145
rect 13452 3136 13504 3188
rect 14188 3179 14240 3188
rect 14188 3145 14197 3179
rect 14197 3145 14231 3179
rect 14231 3145 14240 3179
rect 14832 3179 14884 3188
rect 14188 3136 14240 3145
rect 12072 3068 12124 3120
rect 11152 3043 11204 3052
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 11888 3043 11940 3052
rect 11888 3009 11897 3043
rect 11897 3009 11931 3043
rect 11931 3009 11940 3043
rect 11888 3000 11940 3009
rect 13360 3068 13412 3120
rect 14832 3145 14841 3179
rect 14841 3145 14875 3179
rect 14875 3145 14884 3179
rect 14832 3136 14884 3145
rect 15292 3179 15344 3188
rect 15292 3145 15301 3179
rect 15301 3145 15335 3179
rect 15335 3145 15344 3179
rect 15292 3136 15344 3145
rect 14924 3068 14976 3120
rect 15200 3111 15252 3120
rect 15200 3077 15209 3111
rect 15209 3077 15243 3111
rect 15243 3077 15252 3111
rect 15200 3068 15252 3077
rect 18328 3136 18380 3188
rect 18604 3136 18656 3188
rect 22468 3136 22520 3188
rect 20720 3068 20772 3120
rect 3884 2932 3936 2984
rect 13544 3000 13596 3052
rect 12164 2975 12216 2984
rect 12164 2941 12173 2975
rect 12173 2941 12207 2975
rect 12207 2941 12216 2975
rect 12164 2932 12216 2941
rect 13820 2932 13872 2984
rect 15660 3000 15712 3052
rect 15844 3000 15896 3052
rect 16948 3043 17000 3052
rect 16948 3009 16957 3043
rect 16957 3009 16991 3043
rect 16991 3009 17000 3043
rect 16948 3000 17000 3009
rect 17500 3043 17552 3052
rect 17500 3009 17509 3043
rect 17509 3009 17543 3043
rect 17543 3009 17552 3043
rect 17500 3000 17552 3009
rect 17868 3000 17920 3052
rect 15476 2975 15528 2984
rect 15476 2941 15485 2975
rect 15485 2941 15519 2975
rect 15519 2941 15528 2975
rect 15476 2932 15528 2941
rect 17224 2932 17276 2984
rect 19064 3000 19116 3052
rect 19340 3000 19392 3052
rect 20444 3000 20496 3052
rect 19524 2932 19576 2984
rect 11888 2864 11940 2916
rect 388 2796 440 2848
rect 8300 2796 8352 2848
rect 10692 2796 10744 2848
rect 11796 2796 11848 2848
rect 16396 2796 16448 2848
rect 16948 2864 17000 2916
rect 18604 2864 18656 2916
rect 21364 2864 21416 2916
rect 17500 2796 17552 2848
rect 21548 2796 21600 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 10232 2592 10284 2644
rect 11152 2635 11204 2644
rect 10508 2524 10560 2576
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 11796 2592 11848 2644
rect 13176 2592 13228 2644
rect 14924 2592 14976 2644
rect 16212 2592 16264 2644
rect 18420 2592 18472 2644
rect 18880 2592 18932 2644
rect 19984 2635 20036 2644
rect 19984 2601 19993 2635
rect 19993 2601 20027 2635
rect 20027 2601 20036 2635
rect 19984 2592 20036 2601
rect 20720 2592 20772 2644
rect 15844 2524 15896 2576
rect 17408 2524 17460 2576
rect 19708 2524 19760 2576
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 12164 2388 12216 2440
rect 11060 2320 11112 2372
rect 11796 2320 11848 2372
rect 13820 2388 13872 2440
rect 15568 2456 15620 2508
rect 16028 2456 16080 2508
rect 17776 2456 17828 2508
rect 15936 2388 15988 2440
rect 18512 2388 18564 2440
rect 15752 2320 15804 2372
rect 19156 2320 19208 2372
rect 12532 2252 12584 2304
rect 13084 2252 13136 2304
rect 13544 2252 13596 2304
rect 14188 2252 14240 2304
rect 15476 2295 15528 2304
rect 15476 2261 15485 2295
rect 15485 2261 15519 2295
rect 15519 2261 15528 2295
rect 15476 2252 15528 2261
rect 15568 2252 15620 2304
rect 17040 2252 17092 2304
rect 18696 2252 18748 2304
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
rect 11060 2048 11112 2100
rect 12256 2048 12308 2100
rect 15936 2048 15988 2100
rect 14648 1980 14700 2032
rect 15752 1980 15804 2032
rect 10508 1912 10560 1964
rect 15476 1912 15528 1964
<< metal2 >>
rect 386 22200 442 23000
rect 938 22200 994 23000
rect 1490 22200 1546 23000
rect 1688 22222 1992 22250
rect 400 18737 428 22200
rect 952 18766 980 22200
rect 1504 18902 1532 22200
rect 1492 18896 1544 18902
rect 1492 18838 1544 18844
rect 940 18760 992 18766
rect 386 18728 442 18737
rect 940 18702 992 18708
rect 386 18663 442 18672
rect 1688 6914 1716 22222
rect 1964 22114 1992 22222
rect 2042 22200 2098 23000
rect 2594 22200 2650 23000
rect 3146 22200 3202 23000
rect 3698 22200 3754 23000
rect 4250 22200 4306 23000
rect 4802 22200 4858 23000
rect 5354 22200 5410 23000
rect 5906 22200 5962 23000
rect 6458 22200 6514 23000
rect 7010 22200 7066 23000
rect 7562 22200 7618 23000
rect 8114 22200 8170 23000
rect 8666 22200 8722 23000
rect 9218 22200 9274 23000
rect 9770 22200 9826 23000
rect 10322 22200 10378 23000
rect 10428 22222 10824 22250
rect 2056 22114 2084 22200
rect 1964 22086 2084 22114
rect 2608 18154 2636 22200
rect 2596 18148 2648 18154
rect 2596 18090 2648 18096
rect 3160 18086 3188 22200
rect 3712 20346 3740 22200
rect 3712 20318 3924 20346
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3332 18896 3384 18902
rect 3332 18838 3384 18844
rect 3148 18080 3200 18086
rect 3148 18022 3200 18028
rect 3344 14618 3372 18838
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3896 14278 3924 20318
rect 4068 17604 4120 17610
rect 4068 17546 4120 17552
rect 4080 17241 4108 17546
rect 4264 17338 4292 22200
rect 4620 19712 4672 19718
rect 4620 19654 4672 19660
rect 4632 18873 4660 19654
rect 4816 19310 4844 22200
rect 5172 19712 5224 19718
rect 5172 19654 5224 19660
rect 5368 19666 5396 22200
rect 5632 20256 5684 20262
rect 5630 20224 5632 20233
rect 5684 20224 5686 20233
rect 5630 20159 5686 20168
rect 5724 19984 5776 19990
rect 5724 19926 5776 19932
rect 5736 19718 5764 19926
rect 5724 19712 5776 19718
rect 4988 19440 5040 19446
rect 4988 19382 5040 19388
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4618 18864 4674 18873
rect 4618 18799 4674 18808
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 4066 17232 4122 17241
rect 4066 17167 4122 17176
rect 4160 16448 4212 16454
rect 4160 16390 4212 16396
rect 4172 16250 4200 16390
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4448 14414 4476 18702
rect 4896 18148 4948 18154
rect 4896 18090 4948 18096
rect 4908 17338 4936 18090
rect 4896 17332 4948 17338
rect 4896 17274 4948 17280
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4540 15162 4568 15846
rect 4632 15366 4660 15982
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3896 14074 3924 14214
rect 4448 14074 4476 14350
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 2596 7268 2648 7274
rect 2596 7210 2648 7216
rect 1412 6886 1716 6914
rect 1412 4758 1440 6886
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 1400 4752 1452 4758
rect 1400 4694 1452 4700
rect 940 3936 992 3942
rect 940 3878 992 3884
rect 388 2848 440 2854
rect 388 2790 440 2796
rect 400 800 428 2790
rect 952 800 980 3878
rect 1490 3088 1546 3097
rect 1490 3023 1546 3032
rect 1504 800 1532 3023
rect 2056 800 2084 4966
rect 2608 800 2636 7210
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3528 5817 3556 5850
rect 3514 5808 3570 5817
rect 3514 5743 3570 5752
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3160 800 3188 4082
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 3896 2990 3924 14010
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 3884 2984 3936 2990
rect 3884 2926 3936 2932
rect 4172 2774 4200 7142
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 4080 2746 4200 2774
rect 3712 870 3832 898
rect 3712 800 3740 870
rect 386 0 442 800
rect 938 0 994 800
rect 1490 0 1546 800
rect 2042 0 2098 800
rect 2594 0 2650 800
rect 3146 0 3202 800
rect 3698 0 3754 800
rect 3804 762 3832 870
rect 4080 762 4108 2746
rect 4264 800 4292 7686
rect 4540 6905 4568 14554
rect 4632 9081 4660 15302
rect 4816 15026 4844 15846
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 4804 14476 4856 14482
rect 4804 14418 4856 14424
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4618 9072 4674 9081
rect 4618 9007 4674 9016
rect 4526 6896 4582 6905
rect 4526 6831 4582 6840
rect 4632 3738 4660 9007
rect 4724 8906 4752 14214
rect 4816 9518 4844 14418
rect 5000 12782 5028 19382
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 5000 10146 5028 12038
rect 5092 11257 5120 14758
rect 5184 11762 5212 19654
rect 5368 19638 5488 19666
rect 5724 19654 5776 19660
rect 5356 19508 5408 19514
rect 5356 19450 5408 19456
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5276 13394 5304 19110
rect 5368 16250 5396 19450
rect 5460 19394 5488 19638
rect 5460 19378 5672 19394
rect 5460 19372 5684 19378
rect 5460 19366 5632 19372
rect 5632 19314 5684 19320
rect 5644 18630 5672 19314
rect 5632 18624 5684 18630
rect 5632 18566 5684 18572
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5368 12918 5396 14758
rect 5460 14414 5488 18022
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5552 16522 5580 17070
rect 5540 16516 5592 16522
rect 5540 16458 5592 16464
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5460 14074 5488 14350
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5460 13433 5488 14010
rect 5446 13424 5502 13433
rect 5446 13359 5502 13368
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5356 12912 5408 12918
rect 5356 12854 5408 12860
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 5184 11558 5212 11698
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5078 11248 5134 11257
rect 5078 11183 5134 11192
rect 5000 10118 5120 10146
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 5000 8566 5028 9998
rect 4988 8560 5040 8566
rect 4988 8502 5040 8508
rect 5000 7342 5028 8502
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 5092 5302 5120 10118
rect 5184 7342 5212 11494
rect 5460 10418 5488 13262
rect 5368 10390 5488 10418
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5276 8362 5304 10066
rect 5368 9994 5396 10390
rect 5552 10282 5580 16458
rect 5644 12345 5672 18566
rect 5736 13297 5764 19654
rect 5920 19394 5948 22200
rect 6472 20890 6500 22200
rect 6472 20862 6684 20890
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 6552 20528 6604 20534
rect 6552 20470 6604 20476
rect 6564 20262 6592 20470
rect 6552 20256 6604 20262
rect 6552 20198 6604 20204
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 5920 19366 6040 19394
rect 6012 19310 6040 19366
rect 6000 19304 6052 19310
rect 6000 19246 6052 19252
rect 6012 18630 6040 19246
rect 6000 18624 6052 18630
rect 6000 18566 6052 18572
rect 6012 17377 6040 18566
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 5998 17368 6054 17377
rect 6148 17371 6456 17380
rect 5998 17303 6054 17312
rect 6000 17264 6052 17270
rect 6000 17206 6052 17212
rect 5908 16448 5960 16454
rect 5908 16390 5960 16396
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 5828 14940 5856 15846
rect 5920 15502 5948 16390
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 5828 14912 5948 14940
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5722 13288 5778 13297
rect 5722 13223 5778 13232
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 5736 12986 5764 13126
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5630 12336 5686 12345
rect 5630 12271 5686 12280
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5460 10254 5580 10282
rect 5460 10130 5488 10254
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 5368 9674 5396 9930
rect 5368 9646 5488 9674
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 5276 7954 5304 8298
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5368 7546 5396 8366
rect 5460 7750 5488 9646
rect 5552 8974 5580 10134
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5552 7886 5580 8366
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5184 7206 5212 7278
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5354 6896 5410 6905
rect 5354 6831 5410 6840
rect 5080 5296 5132 5302
rect 5080 5238 5132 5244
rect 5092 5030 5120 5238
rect 5080 5024 5132 5030
rect 5080 4966 5132 4972
rect 4802 4040 4858 4049
rect 4802 3975 4858 3984
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4816 800 4844 3975
rect 5368 800 5396 6831
rect 5644 3602 5672 12174
rect 5736 10810 5764 12786
rect 5828 12594 5856 14214
rect 5920 12850 5948 14912
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5828 12566 5948 12594
rect 5920 12186 5948 12566
rect 6012 12238 6040 17206
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6090 15464 6146 15473
rect 6090 15399 6092 15408
rect 6144 15399 6146 15408
rect 6092 15370 6144 15376
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6184 15088 6236 15094
rect 6184 15030 6236 15036
rect 6196 14618 6224 15030
rect 6184 14612 6236 14618
rect 6184 14554 6236 14560
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6092 13932 6144 13938
rect 6092 13874 6144 13880
rect 6104 13462 6132 13874
rect 6092 13456 6144 13462
rect 6564 13410 6592 20198
rect 6656 18290 6684 20862
rect 6736 20460 6788 20466
rect 6736 20402 6788 20408
rect 6748 19922 6776 20402
rect 7024 19938 7052 22200
rect 7576 20398 7604 22200
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 7564 20392 7616 20398
rect 7564 20334 7616 20340
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 6736 19916 6788 19922
rect 6736 19858 6788 19864
rect 6840 19910 7052 19938
rect 6840 19514 6868 19910
rect 7012 19848 7064 19854
rect 7012 19790 7064 19796
rect 7196 19848 7248 19854
rect 7196 19790 7248 19796
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 6840 19224 6868 19450
rect 6748 19196 6868 19224
rect 6748 18426 6776 19196
rect 6828 18760 6880 18766
rect 6828 18702 6880 18708
rect 6736 18420 6788 18426
rect 6736 18362 6788 18368
rect 6644 18284 6696 18290
rect 6644 18226 6696 18232
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6092 13398 6144 13404
rect 6472 13382 6592 13410
rect 6472 13326 6500 13382
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 6564 12850 6592 13262
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6550 12744 6606 12753
rect 6550 12679 6606 12688
rect 6564 12238 6592 12679
rect 5828 12158 5948 12186
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 9926 5764 10406
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5736 9586 5764 9862
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5724 9444 5776 9450
rect 5724 9386 5776 9392
rect 5736 7342 5764 9386
rect 5828 8906 5856 12158
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 5920 11082 5948 12038
rect 6012 11218 6040 12038
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6182 11792 6238 11801
rect 6092 11756 6144 11762
rect 6182 11727 6238 11736
rect 6092 11698 6144 11704
rect 6104 11354 6132 11698
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6104 11121 6132 11290
rect 6090 11112 6146 11121
rect 5908 11076 5960 11082
rect 6090 11047 6146 11056
rect 5908 11018 5960 11024
rect 6196 10996 6224 11727
rect 6472 11014 6500 11834
rect 6012 10968 6224 10996
rect 6460 11008 6512 11014
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 5920 10130 5948 10746
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5920 9518 5948 10066
rect 6012 10033 6040 10968
rect 6460 10950 6512 10956
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 5998 10024 6054 10033
rect 5998 9959 6054 9968
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 6012 9722 6040 9862
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 5816 8900 5868 8906
rect 5816 8842 5868 8848
rect 6012 7954 6040 8978
rect 6288 8838 6316 9454
rect 6564 9178 6592 10542
rect 6656 9654 6684 16934
rect 6748 15094 6776 17478
rect 6840 15162 6868 18702
rect 6932 18358 6960 19654
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6932 15638 6960 15982
rect 6920 15632 6972 15638
rect 6920 15574 6972 15580
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6736 15088 6788 15094
rect 6736 15030 6788 15036
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6748 13938 6776 14894
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6748 12850 6776 13466
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6748 12102 6776 12242
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6748 10810 6776 12038
rect 6840 11898 6868 13126
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 6828 11756 6880 11762
rect 6828 11698 6880 11704
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6656 9178 6684 9454
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6748 8090 6776 10610
rect 6840 10130 6868 11698
rect 6932 10606 6960 14214
rect 7024 11898 7052 19790
rect 7104 19780 7156 19786
rect 7104 19722 7156 19728
rect 7116 17746 7144 19722
rect 7208 18834 7236 19790
rect 7300 19174 7328 20198
rect 7392 19718 7420 20334
rect 7380 19712 7432 19718
rect 7380 19654 7432 19660
rect 7288 19168 7340 19174
rect 7288 19110 7340 19116
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7392 18714 7420 19654
rect 7760 19446 7788 20402
rect 7748 19440 7800 19446
rect 7748 19382 7800 19388
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 7300 18686 7420 18714
rect 7104 17740 7156 17746
rect 7104 17682 7156 17688
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7300 15858 7328 18686
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7392 17746 7420 18566
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7392 16046 7420 17682
rect 7484 16250 7512 18022
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7668 17338 7696 17614
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7564 16516 7616 16522
rect 7564 16458 7616 16464
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7576 16130 7604 16458
rect 7484 16102 7604 16130
rect 7656 16108 7708 16114
rect 7380 16040 7432 16046
rect 7380 15982 7432 15988
rect 7484 15910 7512 16102
rect 7656 16050 7708 16056
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 7562 16008 7618 16017
rect 7562 15943 7618 15952
rect 7472 15904 7524 15910
rect 7116 15570 7144 15846
rect 7300 15830 7420 15858
rect 7472 15846 7524 15852
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7300 14929 7328 15302
rect 7286 14920 7342 14929
rect 7286 14855 7342 14864
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 7116 14006 7144 14282
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 7116 11762 7144 13942
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7116 11150 7144 11494
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 7208 11098 7236 12038
rect 7300 11354 7328 14214
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7208 11070 7328 11098
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6826 10024 6882 10033
rect 6826 9959 6882 9968
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5920 7546 5948 7686
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 5724 7336 5776 7342
rect 6644 7336 6696 7342
rect 5724 7278 5776 7284
rect 5906 7304 5962 7313
rect 6644 7278 6696 7284
rect 5906 7239 5962 7248
rect 5920 7206 5948 7239
rect 6656 7206 6684 7278
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 5920 4146 5948 7142
rect 6656 6934 6684 7142
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 6748 6866 6776 7346
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 6840 5234 6868 9959
rect 7024 9926 7052 10950
rect 7208 10810 7236 10950
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7116 10198 7144 10406
rect 7300 10266 7328 11070
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7300 10062 7328 10202
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7208 8974 7236 9318
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7300 8838 7328 9318
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6932 7954 6960 8230
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 7392 4622 7420 15830
rect 7484 10538 7512 15846
rect 7576 15473 7604 15943
rect 7562 15464 7618 15473
rect 7562 15399 7564 15408
rect 7616 15399 7618 15408
rect 7564 15370 7616 15376
rect 7668 15366 7696 16050
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7576 11354 7604 14962
rect 7668 12102 7696 15302
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7654 11928 7710 11937
rect 7654 11863 7710 11872
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7484 8820 7512 9862
rect 7564 9512 7616 9518
rect 7668 9500 7696 11863
rect 7760 9674 7788 16050
rect 7852 14618 7880 19314
rect 8024 19236 8076 19242
rect 8024 19178 8076 19184
rect 8036 18154 8064 19178
rect 8128 18850 8156 22200
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8208 19440 8260 19446
rect 8208 19382 8260 19388
rect 8220 19310 8248 19382
rect 8208 19304 8260 19310
rect 8208 19246 8260 19252
rect 8404 18970 8432 20198
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8128 18822 8248 18850
rect 8116 18692 8168 18698
rect 8116 18634 8168 18640
rect 8128 18222 8156 18634
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8024 18148 8076 18154
rect 8024 18090 8076 18096
rect 8220 17649 8248 18822
rect 8206 17640 8262 17649
rect 8206 17575 8262 17584
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7852 12986 7880 13126
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7852 12889 7880 12922
rect 7838 12880 7894 12889
rect 7838 12815 7894 12824
rect 7944 12434 7972 15574
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 8036 14958 8064 15098
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 7852 12406 7972 12434
rect 7852 11937 7880 12406
rect 8128 12322 8156 12786
rect 7944 12294 8156 12322
rect 7944 12238 7972 12294
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 7838 11928 7894 11937
rect 7838 11863 7894 11872
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7852 11354 7880 11698
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 7944 10810 7972 12174
rect 8220 11898 8248 17274
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8312 13394 8340 13670
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8312 12918 8340 13330
rect 8404 13258 8432 13670
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8404 12434 8432 13194
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8496 12646 8524 12922
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8312 12406 8432 12434
rect 8482 12472 8538 12481
rect 8482 12407 8538 12416
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 7944 10062 7972 10610
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7944 9926 7972 9998
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7760 9646 7880 9674
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7616 9472 7696 9500
rect 7564 9454 7616 9460
rect 7656 8832 7708 8838
rect 7484 8792 7656 8820
rect 7656 8774 7708 8780
rect 7760 8090 7788 9522
rect 7852 9110 7880 9646
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7852 5166 7880 8774
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 6550 3904 6606 3913
rect 6550 3839 6606 3848
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5920 800 5948 3674
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 6564 1986 6592 3839
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 6472 1958 6592 1986
rect 6472 800 6500 1958
rect 7024 800 7052 3334
rect 7944 2774 7972 9862
rect 8036 6118 8064 11834
rect 8206 11792 8262 11801
rect 8206 11727 8262 11736
rect 8220 11218 8248 11727
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8114 10160 8170 10169
rect 8114 10095 8170 10104
rect 8128 9450 8156 10095
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 8220 7410 8248 10202
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 7944 2746 8064 2774
rect 7576 870 7696 898
rect 7576 800 7604 870
rect 3804 734 4108 762
rect 4250 0 4306 800
rect 4802 0 4858 800
rect 5354 0 5410 800
rect 5906 0 5962 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7562 0 7618 800
rect 7668 762 7696 870
rect 8036 762 8064 2746
rect 8128 800 8156 5306
rect 8220 4826 8248 7346
rect 8312 5914 8340 12406
rect 8496 11778 8524 12407
rect 8404 11750 8524 11778
rect 8588 11778 8616 20198
rect 8680 17218 8708 22200
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 9034 18728 9090 18737
rect 9034 18663 9090 18672
rect 9048 18630 9076 18663
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 9232 18426 9260 22200
rect 9310 19816 9366 19825
rect 9310 19751 9366 19760
rect 9324 19718 9352 19751
rect 9312 19712 9364 19718
rect 9312 19654 9364 19660
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 8680 17190 8800 17218
rect 8772 17105 8800 17190
rect 8758 17096 8814 17105
rect 8668 17060 8720 17066
rect 9140 17066 9168 17614
rect 8758 17031 8814 17040
rect 9128 17060 9180 17066
rect 8668 17002 8720 17008
rect 9128 17002 9180 17008
rect 8680 16794 8708 17002
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 9140 16590 9168 17002
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9140 16046 9168 16526
rect 9128 16040 9180 16046
rect 9128 15982 9180 15988
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 9140 15366 9168 15982
rect 9128 15360 9180 15366
rect 9128 15302 9180 15308
rect 9140 14958 9168 15302
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 9324 14804 9352 19654
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9692 18766 9720 19246
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9416 15026 9444 15846
rect 9600 15434 9628 16390
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 9140 14776 9352 14804
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8680 13530 8708 13670
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8680 12434 8708 13466
rect 9140 13410 9168 14776
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9048 13382 9168 13410
rect 9048 12646 9076 13382
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 8680 12406 8800 12434
rect 8588 11750 8708 11778
rect 8404 11694 8432 11750
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8404 10849 8432 10950
rect 8390 10840 8446 10849
rect 8390 10775 8446 10784
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 8404 9994 8432 10678
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8390 7032 8446 7041
rect 8390 6967 8392 6976
rect 8444 6967 8446 6976
rect 8392 6938 8444 6944
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8312 2854 8340 5578
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 7668 734 8064 762
rect 8114 0 8170 800
rect 8404 762 8432 6938
rect 8496 5846 8524 11494
rect 8588 10810 8616 11630
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8574 10704 8630 10713
rect 8574 10639 8630 10648
rect 8588 10033 8616 10639
rect 8574 10024 8630 10033
rect 8574 9959 8630 9968
rect 8588 9926 8616 9959
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8588 5370 8616 9862
rect 8680 9654 8708 11750
rect 8772 11558 8800 12406
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 9048 12238 9076 12310
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 9140 12102 9168 13262
rect 9232 12753 9260 14214
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9218 12744 9274 12753
rect 9218 12679 9274 12688
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 8760 11552 8812 11558
rect 8760 11494 8812 11500
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 9034 10976 9090 10985
rect 9034 10911 9090 10920
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 8864 10577 8892 10610
rect 8850 10568 8906 10577
rect 8850 10503 8906 10512
rect 9048 10452 9076 10911
rect 9140 10606 9168 11834
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9048 10424 9168 10452
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 8772 9466 8800 9522
rect 8680 9438 8800 9466
rect 8680 8838 8708 9438
rect 9140 9330 9168 10424
rect 9232 10130 9260 12582
rect 9324 11558 9352 12786
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9324 10130 9352 11494
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9232 9518 9260 10066
rect 9310 9616 9366 9625
rect 9310 9551 9312 9560
rect 9364 9551 9366 9560
rect 9312 9522 9364 9528
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9140 9302 9352 9330
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8680 8022 8708 8502
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 9140 7954 9168 8230
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8496 3194 8524 4966
rect 8680 3942 8708 7686
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 9218 6352 9274 6361
rect 9128 6316 9180 6322
rect 9218 6287 9274 6296
rect 9128 6258 9180 6264
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8772 5234 8800 5306
rect 8944 5296 8996 5302
rect 8944 5238 8996 5244
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8956 5030 8984 5238
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 9140 4826 9168 6258
rect 9232 5914 9260 6287
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9324 5302 9352 9302
rect 9416 9042 9444 14962
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9508 11286 9536 12038
rect 9496 11280 9548 11286
rect 9496 11222 9548 11228
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9416 7478 9444 8570
rect 9404 7472 9456 7478
rect 9404 7414 9456 7420
rect 9508 6186 9536 11222
rect 9600 9178 9628 15370
rect 9692 14890 9720 18226
rect 9784 18057 9812 22200
rect 10336 22114 10364 22200
rect 10428 22114 10456 22222
rect 10336 22086 10456 22114
rect 10232 21072 10284 21078
rect 10232 21014 10284 21020
rect 10244 20466 10272 21014
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 10324 20256 10376 20262
rect 10324 20198 10376 20204
rect 10336 19786 10364 20198
rect 10520 19961 10548 20402
rect 10506 19952 10562 19961
rect 10506 19887 10562 19896
rect 10324 19780 10376 19786
rect 10324 19722 10376 19728
rect 10692 19780 10744 19786
rect 10692 19722 10744 19728
rect 10336 19446 10364 19722
rect 10324 19440 10376 19446
rect 10324 19382 10376 19388
rect 10704 18986 10732 19722
rect 10428 18958 10732 18986
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9876 18290 9904 18634
rect 10336 18290 10364 18702
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 10140 18284 10192 18290
rect 10140 18226 10192 18232
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 9770 18048 9826 18057
rect 9770 17983 9826 17992
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 9784 14414 9812 17818
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9876 14618 9904 17138
rect 9956 16516 10008 16522
rect 9956 16458 10008 16464
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9692 13190 9720 14010
rect 9968 13938 9996 16458
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9692 10441 9720 12106
rect 9876 10674 9904 12174
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 9678 10432 9734 10441
rect 9678 10367 9734 10376
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9600 8922 9628 9114
rect 9692 9042 9720 9862
rect 9876 9722 9904 9862
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9862 9480 9918 9489
rect 9862 9415 9918 9424
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9600 8894 9720 8922
rect 9692 8514 9720 8894
rect 9600 8486 9720 8514
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9600 7954 9628 8486
rect 9680 8424 9732 8430
rect 9678 8392 9680 8401
rect 9732 8392 9734 8401
rect 9678 8327 9734 8336
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9784 7834 9812 8502
rect 9600 7806 9812 7834
rect 9600 7546 9628 7806
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9876 6866 9904 9415
rect 9968 9178 9996 9930
rect 9956 9172 10008 9178
rect 9956 9114 10008 9120
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9496 6180 9548 6186
rect 9496 6122 9548 6128
rect 9508 5778 9536 6122
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9692 5710 9720 6598
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9600 5370 9628 5510
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 9784 4826 9812 6190
rect 9956 5840 10008 5846
rect 9956 5782 10008 5788
rect 10060 5794 10088 17274
rect 10152 15638 10180 18226
rect 10428 15722 10456 18958
rect 10600 18896 10652 18902
rect 10600 18838 10652 18844
rect 10612 18698 10640 18838
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10520 17082 10548 18566
rect 10704 18086 10732 18566
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10520 17054 10640 17082
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 10520 16114 10548 16934
rect 10612 16454 10640 17054
rect 10704 16998 10732 18022
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10704 16590 10732 16934
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10600 16448 10652 16454
rect 10600 16390 10652 16396
rect 10508 16108 10560 16114
rect 10508 16050 10560 16056
rect 10520 15858 10548 16050
rect 10704 16046 10732 16526
rect 10692 16040 10744 16046
rect 10692 15982 10744 15988
rect 10520 15830 10732 15858
rect 10428 15694 10640 15722
rect 10140 15632 10192 15638
rect 10140 15574 10192 15580
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10336 14498 10364 15438
rect 10244 14470 10364 14498
rect 10138 14240 10194 14249
rect 10138 14175 10194 14184
rect 10152 14006 10180 14175
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10244 13530 10272 14470
rect 10324 14340 10376 14346
rect 10324 14282 10376 14288
rect 10336 14113 10364 14282
rect 10322 14104 10378 14113
rect 10322 14039 10378 14048
rect 10324 14000 10376 14006
rect 10324 13942 10376 13948
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10138 10840 10194 10849
rect 10138 10775 10140 10784
rect 10192 10775 10194 10784
rect 10140 10746 10192 10752
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10152 8634 10180 8910
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10138 8256 10194 8265
rect 10138 8191 10194 8200
rect 10152 8090 10180 8191
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10152 7478 10180 8026
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10152 5914 10180 6258
rect 10244 6254 10272 13466
rect 10336 12170 10364 13942
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10428 12442 10456 13126
rect 10416 12436 10468 12442
rect 10612 12434 10640 15694
rect 10416 12378 10468 12384
rect 10520 12406 10640 12434
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10428 10810 10456 10950
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10336 8090 10364 10542
rect 10520 10062 10548 12406
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10612 10606 10640 12242
rect 10704 11132 10732 15830
rect 10796 11642 10824 22222
rect 10874 22200 10930 23000
rect 11426 22200 11482 23000
rect 11532 22222 11744 22250
rect 10888 17338 10916 22200
rect 11440 22114 11468 22200
rect 11532 22114 11560 22222
rect 11440 22086 11560 22114
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 11716 20602 11744 22222
rect 11978 22200 12034 23000
rect 12530 22200 12586 23000
rect 13082 22200 13138 23000
rect 13634 22200 13690 23000
rect 14186 22200 14242 23000
rect 14738 22200 14794 23000
rect 15290 22200 15346 23000
rect 15842 22200 15898 23000
rect 16394 22200 16450 23000
rect 16946 22200 17002 23000
rect 17498 22200 17554 23000
rect 18050 22200 18106 23000
rect 18602 22200 18658 23000
rect 19154 22200 19210 23000
rect 19706 22200 19762 23000
rect 20258 22200 20314 23000
rect 20810 22200 20866 23000
rect 21362 22200 21418 23000
rect 21560 22222 21864 22250
rect 11992 21078 12020 22200
rect 11980 21072 12032 21078
rect 11980 21014 12032 21020
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 12162 20360 12218 20369
rect 12162 20295 12218 20304
rect 12176 20262 12204 20295
rect 10968 20256 11020 20262
rect 10968 20198 11020 20204
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 10980 19854 11008 20198
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 10980 19242 11008 19790
rect 11072 19786 11560 19802
rect 11072 19780 11572 19786
rect 11072 19774 11520 19780
rect 11072 19718 11100 19774
rect 11520 19722 11572 19728
rect 11060 19712 11112 19718
rect 11428 19712 11480 19718
rect 11060 19654 11112 19660
rect 11164 19672 11428 19700
rect 10968 19236 11020 19242
rect 10968 19178 11020 19184
rect 10980 18630 11008 19178
rect 10968 18624 11020 18630
rect 10968 18566 11020 18572
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 11072 18408 11100 18566
rect 10980 18380 11100 18408
rect 10980 17542 11008 18380
rect 11164 18358 11192 19672
rect 11428 19654 11480 19660
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11244 19372 11296 19378
rect 11244 19314 11296 19320
rect 11152 18352 11204 18358
rect 11152 18294 11204 18300
rect 11256 18136 11284 19314
rect 11704 19304 11756 19310
rect 11704 19246 11756 19252
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11348 18193 11376 18226
rect 11164 18108 11284 18136
rect 11334 18184 11390 18193
rect 11716 18154 11744 19246
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11900 18290 11928 19110
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11334 18119 11390 18128
rect 11704 18148 11756 18154
rect 11164 17542 11192 18108
rect 11704 18090 11756 18096
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 11072 15366 11100 15846
rect 11164 15706 11192 17478
rect 11256 16998 11284 17478
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 11716 16946 11744 17682
rect 11888 17604 11940 17610
rect 11888 17546 11940 17552
rect 11716 16918 11836 16946
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 11072 14890 11100 15302
rect 11060 14884 11112 14890
rect 11060 14826 11112 14832
rect 11072 14414 11100 14826
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 11072 14278 11100 14350
rect 11060 14272 11112 14278
rect 11164 14249 11192 14758
rect 11060 14214 11112 14220
rect 11150 14240 11206 14249
rect 11072 13870 11100 14214
rect 11150 14175 11206 14184
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10888 12238 10916 12718
rect 11072 12238 11100 12854
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11164 12306 11192 12582
rect 11152 12300 11204 12306
rect 11152 12242 11204 12248
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11072 12084 11100 12174
rect 11152 12096 11204 12102
rect 11072 12056 11152 12084
rect 11152 12038 11204 12044
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 10796 11614 11008 11642
rect 11072 11626 11100 11766
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10888 11286 10916 11494
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 10704 11104 10916 11132
rect 10782 10976 10838 10985
rect 10782 10911 10838 10920
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10428 9178 10456 9862
rect 10520 9722 10548 9862
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10704 8922 10732 10746
rect 10796 10577 10824 10911
rect 10782 10568 10838 10577
rect 10782 10503 10838 10512
rect 10888 9110 10916 11104
rect 10980 10985 11008 11614
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 11164 11558 11192 12038
rect 11256 11830 11284 16390
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11716 15706 11744 16730
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11716 14618 11744 15302
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11808 13841 11836 16918
rect 11794 13832 11850 13841
rect 11794 13767 11850 13776
rect 11900 13530 11928 17546
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11244 11824 11296 11830
rect 11244 11766 11296 11772
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10966 10976 11022 10985
rect 10966 10911 11022 10920
rect 11072 10690 11100 11154
rect 11164 11150 11192 11494
rect 11256 11150 11284 11766
rect 11336 11688 11388 11694
rect 11716 11642 11744 13466
rect 11992 12968 12020 19858
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 12084 18698 12112 19450
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 12084 16454 12112 16526
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 12084 15162 12112 16390
rect 12176 16017 12204 20198
rect 12544 19802 12572 22200
rect 12624 20460 12676 20466
rect 12624 20402 12676 20408
rect 12452 19774 12572 19802
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12268 18358 12296 19654
rect 12452 19242 12480 19774
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12544 19446 12572 19654
rect 12532 19440 12584 19446
rect 12532 19382 12584 19388
rect 12440 19236 12492 19242
rect 12440 19178 12492 19184
rect 12636 19174 12664 20402
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12728 19961 12756 20198
rect 13096 20058 13124 22200
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 12714 19952 12770 19961
rect 12714 19887 12770 19896
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12728 18630 12756 19887
rect 13648 19786 13676 22200
rect 14200 20482 14228 22200
rect 14200 20454 14320 20482
rect 13728 20324 13780 20330
rect 13728 20266 13780 20272
rect 13636 19780 13688 19786
rect 13636 19722 13688 19728
rect 13740 19446 13768 20266
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13728 19440 13780 19446
rect 13728 19382 13780 19388
rect 13268 18692 13320 18698
rect 13268 18634 13320 18640
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12268 16658 12296 18294
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12360 16998 12388 17206
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 12162 16008 12218 16017
rect 12162 15943 12218 15952
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 11900 12940 12020 12968
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11808 11762 11836 12582
rect 11900 11762 11928 12940
rect 12084 12918 12112 13262
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 11992 11778 12020 12786
rect 12176 11801 12204 15846
rect 12268 14822 12296 16050
rect 12636 15473 12664 18158
rect 12716 17060 12768 17066
rect 12716 17002 12768 17008
rect 12728 16522 12756 17002
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12622 15464 12678 15473
rect 12622 15399 12678 15408
rect 12728 15314 12756 16458
rect 12820 16250 12848 18566
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12912 15337 12940 17138
rect 12992 16788 13044 16794
rect 12992 16730 13044 16736
rect 12636 15286 12756 15314
rect 12898 15328 12954 15337
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12254 13832 12310 13841
rect 12254 13767 12310 13776
rect 12268 13530 12296 13767
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 12162 11792 12218 11801
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11888 11756 11940 11762
rect 11992 11750 12112 11778
rect 11888 11698 11940 11704
rect 11336 11630 11388 11636
rect 11152 11144 11204 11150
rect 11152 11086 11204 11092
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 10980 10662 11100 10690
rect 11256 10674 11284 11086
rect 11348 11082 11376 11630
rect 11440 11614 11744 11642
rect 11440 11218 11468 11614
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11612 10736 11664 10742
rect 11612 10678 11664 10684
rect 11152 10668 11204 10674
rect 10980 10538 11008 10662
rect 11152 10610 11204 10616
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10968 10532 11020 10538
rect 10968 10474 11020 10480
rect 10876 9104 10928 9110
rect 10876 9046 10928 9052
rect 10704 8894 10824 8922
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10600 8424 10652 8430
rect 10704 8401 10732 8774
rect 10600 8366 10652 8372
rect 10690 8392 10746 8401
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10416 8016 10468 8022
rect 10416 7958 10468 7964
rect 10232 6248 10284 6254
rect 10232 6190 10284 6196
rect 10428 5914 10456 7958
rect 10612 7546 10640 8366
rect 10690 8327 10746 8336
rect 10704 7818 10732 8327
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10704 7478 10732 7754
rect 10692 7472 10744 7478
rect 10506 7440 10562 7449
rect 10692 7414 10744 7420
rect 10506 7375 10562 7384
rect 10520 6458 10548 7375
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10612 6662 10640 6734
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 9968 5370 9996 5782
rect 10060 5766 10548 5794
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 10060 4690 10088 5102
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 8864 4282 8892 4558
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 10048 4548 10100 4554
rect 10048 4490 10100 4496
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 9140 3641 9168 4422
rect 9692 4282 9720 4490
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 10060 3942 10088 4490
rect 10048 3936 10100 3942
rect 9770 3904 9826 3913
rect 10048 3878 10100 3884
rect 9770 3839 9826 3848
rect 9220 3664 9272 3670
rect 9126 3632 9182 3641
rect 9220 3606 9272 3612
rect 9126 3567 9182 3576
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 8588 870 8708 898
rect 8588 762 8616 870
rect 8680 800 8708 870
rect 9232 800 9260 3606
rect 9784 3097 9812 3839
rect 10060 3738 10088 3878
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 9862 3224 9918 3233
rect 10152 3194 10180 5238
rect 10414 4720 10470 4729
rect 10324 4684 10376 4690
rect 10414 4655 10470 4664
rect 10324 4626 10376 4632
rect 10336 4282 10364 4626
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 9862 3159 9864 3168
rect 9916 3159 9918 3168
rect 10140 3188 10192 3194
rect 9864 3130 9916 3136
rect 10140 3130 10192 3136
rect 9770 3088 9826 3097
rect 9770 3023 9826 3032
rect 9784 800 9812 3023
rect 10244 2650 10272 3538
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10428 2258 10456 4655
rect 10520 2582 10548 5766
rect 10612 5137 10640 6598
rect 10704 6254 10732 6802
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10796 5370 10824 8894
rect 10888 8430 10916 9046
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10980 8022 11008 8366
rect 10968 8016 11020 8022
rect 10968 7958 11020 7964
rect 11072 7546 11100 10542
rect 11164 10130 11192 10610
rect 11624 10130 11652 10678
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11612 10124 11664 10130
rect 11612 10066 11664 10072
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11256 9722 11284 9862
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11716 9654 11744 11494
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11808 9353 11836 11698
rect 11978 11656 12034 11665
rect 11978 11591 12034 11600
rect 11992 9586 12020 11591
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11888 9376 11940 9382
rect 11794 9344 11850 9353
rect 11940 9336 12020 9364
rect 11888 9318 11940 9324
rect 11794 9279 11850 9288
rect 11992 9178 12020 9336
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11152 8968 11204 8974
rect 12084 8956 12112 11750
rect 12162 11727 12218 11736
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12176 11286 12204 11630
rect 12164 11280 12216 11286
rect 12164 11222 12216 11228
rect 12164 11008 12216 11014
rect 12162 10976 12164 10985
rect 12216 10976 12218 10985
rect 12162 10911 12218 10920
rect 12162 10840 12218 10849
rect 12162 10775 12164 10784
rect 12216 10775 12218 10784
rect 12164 10746 12216 10752
rect 12268 10690 12296 12786
rect 12176 10662 12296 10690
rect 12176 9738 12204 10662
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12268 10062 12296 10542
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12176 9710 12296 9738
rect 12162 9616 12218 9625
rect 12162 9551 12218 9560
rect 12176 9450 12204 9551
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 11152 8910 11204 8916
rect 11992 8928 12112 8956
rect 11164 8838 11192 8910
rect 11992 8888 12020 8928
rect 11992 8860 12112 8888
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11164 7426 11192 8774
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 10980 7398 11192 7426
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 10888 6662 10916 6870
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10980 6474 11008 7398
rect 11150 6896 11206 6905
rect 11150 6831 11152 6840
rect 11204 6831 11206 6840
rect 11152 6802 11204 6808
rect 10888 6446 11008 6474
rect 11164 6458 11192 6802
rect 11256 6798 11284 8230
rect 11900 8129 11928 8298
rect 11886 8120 11942 8129
rect 11886 8055 11942 8064
rect 11992 7750 12020 8434
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 11992 7546 12020 7686
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 12084 7342 12112 8860
rect 12268 8616 12296 9710
rect 12176 8588 12296 8616
rect 12176 7954 12204 8588
rect 12360 8514 12388 15098
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12544 12102 12572 13874
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12636 11626 12664 15286
rect 12898 15263 12954 15272
rect 13004 15144 13032 16730
rect 13280 16590 13308 18634
rect 13832 18358 13860 19654
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13544 18080 13596 18086
rect 13372 18028 13544 18034
rect 13372 18022 13596 18028
rect 13372 18006 13584 18022
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13280 16046 13308 16390
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 13280 15502 13308 15982
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 12820 15116 13032 15144
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12728 12442 12756 12854
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12624 11620 12676 11626
rect 12624 11562 12676 11568
rect 12636 11286 12664 11562
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10810 12480 10950
rect 12544 10849 12572 11154
rect 12624 11144 12676 11150
rect 12622 11112 12624 11121
rect 12676 11112 12678 11121
rect 12622 11047 12678 11056
rect 12530 10840 12586 10849
rect 12440 10804 12492 10810
rect 12530 10775 12586 10784
rect 12440 10746 12492 10752
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12268 8486 12388 8514
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12176 7478 12204 7686
rect 12164 7472 12216 7478
rect 12164 7414 12216 7420
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 11978 7032 12034 7041
rect 11978 6967 12034 6976
rect 11992 6866 12020 6967
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11152 6452 11204 6458
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 10598 5128 10654 5137
rect 10598 5063 10654 5072
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10598 4176 10654 4185
rect 10598 4111 10654 4120
rect 10612 3194 10640 4111
rect 10704 4078 10732 4422
rect 10692 4072 10744 4078
rect 10888 4049 10916 6446
rect 11152 6394 11204 6400
rect 11152 6180 11204 6186
rect 11152 6122 11204 6128
rect 11164 5710 11192 6122
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11900 5914 11928 6054
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 10692 4014 10744 4020
rect 10874 4040 10930 4049
rect 10704 3602 10732 4014
rect 10874 3975 10930 3984
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10704 2854 10732 3538
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 10508 2576 10560 2582
rect 10508 2518 10560 2524
rect 10336 2230 10456 2258
rect 10336 800 10364 2230
rect 10520 1970 10548 2518
rect 10508 1964 10560 1970
rect 10508 1906 10560 1912
rect 10888 800 10916 3538
rect 10980 3534 11008 5510
rect 11164 5370 11192 5510
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 11164 4554 11192 5034
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 11058 4040 11114 4049
rect 11058 3975 11114 3984
rect 11072 3670 11100 3975
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11060 3664 11112 3670
rect 11060 3606 11112 3612
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11072 2961 11100 3402
rect 11164 3058 11192 3402
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11058 2952 11114 2961
rect 11058 2887 11114 2896
rect 11072 2774 11100 2887
rect 11072 2746 11192 2774
rect 11164 2650 11192 2746
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11060 2372 11112 2378
rect 11060 2314 11112 2320
rect 11072 2106 11100 2314
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11060 2100 11112 2106
rect 11060 2042 11112 2048
rect 11440 870 11560 898
rect 11440 800 11468 870
rect 8404 734 8616 762
rect 8666 0 8722 800
rect 9218 0 9274 800
rect 9770 0 9826 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11426 0 11482 800
rect 11532 762 11560 870
rect 11716 762 11744 3878
rect 11900 3058 11928 4422
rect 12084 3534 12112 7142
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12176 6225 12204 6258
rect 12162 6216 12218 6225
rect 12162 6151 12218 6160
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 12176 4282 12204 5102
rect 12268 4690 12296 8486
rect 12452 8378 12480 10406
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12530 9344 12586 9353
rect 12530 9279 12586 9288
rect 12544 9042 12572 9279
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12360 8350 12480 8378
rect 12360 8265 12388 8350
rect 12532 8288 12584 8294
rect 12346 8256 12402 8265
rect 12532 8230 12584 8236
rect 12346 8191 12402 8200
rect 12440 8016 12492 8022
rect 12346 7984 12402 7993
rect 12440 7958 12492 7964
rect 12346 7919 12402 7928
rect 12360 5778 12388 7919
rect 12452 7818 12480 7958
rect 12544 7886 12572 8230
rect 12636 8090 12664 9862
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12728 7954 12756 12038
rect 12820 10470 12848 15116
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12912 11898 12940 14962
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12898 11384 12954 11393
rect 12898 11319 12954 11328
rect 12912 11286 12940 11319
rect 12900 11280 12952 11286
rect 12900 11222 12952 11228
rect 12898 11112 12954 11121
rect 12898 11047 12900 11056
rect 12952 11047 12954 11056
rect 12900 11018 12952 11024
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12898 10432 12954 10441
rect 12898 10367 12954 10376
rect 12806 10296 12862 10305
rect 12806 10231 12808 10240
rect 12860 10231 12862 10240
rect 12808 10202 12860 10208
rect 12806 9616 12862 9625
rect 12806 9551 12862 9560
rect 12820 9518 12848 9551
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12808 8628 12860 8634
rect 12808 8570 12860 8576
rect 12716 7948 12768 7954
rect 12716 7890 12768 7896
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12544 6769 12572 6802
rect 12530 6760 12586 6769
rect 12530 6695 12586 6704
rect 12532 6656 12584 6662
rect 12532 6598 12584 6604
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12346 5672 12402 5681
rect 12346 5607 12402 5616
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12164 4276 12216 4282
rect 12164 4218 12216 4224
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 11888 2916 11940 2922
rect 11888 2858 11940 2864
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11808 2650 11836 2790
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 11808 2378 11836 2586
rect 11796 2372 11848 2378
rect 11796 2314 11848 2320
rect 11900 1442 11928 2858
rect 11992 2446 12020 3402
rect 12072 3120 12124 3126
rect 12070 3088 12072 3097
rect 12124 3088 12126 3097
rect 12070 3023 12126 3032
rect 12164 2984 12216 2990
rect 12164 2926 12216 2932
rect 12176 2446 12204 2926
rect 12360 2774 12388 5607
rect 12452 4146 12480 6394
rect 12544 5710 12572 6598
rect 12636 6458 12664 7754
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12728 6497 12756 6666
rect 12714 6488 12770 6497
rect 12624 6452 12676 6458
rect 12714 6423 12770 6432
rect 12624 6394 12676 6400
rect 12716 6384 12768 6390
rect 12716 6326 12768 6332
rect 12532 5704 12584 5710
rect 12532 5646 12584 5652
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12544 4282 12572 4422
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12728 4146 12756 6326
rect 12820 6225 12848 8570
rect 12912 6390 12940 10367
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 13004 6322 13032 12106
rect 13096 11218 13124 13194
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 13084 11008 13136 11014
rect 13082 10976 13084 10985
rect 13136 10976 13138 10985
rect 13082 10911 13138 10920
rect 13096 7750 13124 10911
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 13096 6934 13124 7346
rect 13188 7018 13216 14010
rect 13280 9738 13308 14554
rect 13372 9926 13400 18006
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13464 16794 13492 16934
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13452 16516 13504 16522
rect 13452 16458 13504 16464
rect 13464 14278 13492 16458
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13648 14074 13676 14962
rect 13740 14822 13768 15302
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13740 14278 13768 14758
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13556 13530 13584 13670
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13280 9710 13400 9738
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13280 9042 13308 9522
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13280 7857 13308 8366
rect 13266 7848 13322 7857
rect 13266 7783 13322 7792
rect 13188 6990 13308 7018
rect 13084 6928 13136 6934
rect 13084 6870 13136 6876
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 12900 6248 12952 6254
rect 12806 6216 12862 6225
rect 12900 6190 12952 6196
rect 12806 6151 12862 6160
rect 12912 5914 12940 6190
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 13004 5250 13032 6258
rect 12820 5222 13032 5250
rect 12820 5166 12848 5222
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 13004 4622 13032 5102
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12452 3534 12480 4082
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12820 3738 12848 3878
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 13096 3398 13124 6870
rect 13174 6760 13230 6769
rect 13174 6695 13230 6704
rect 13188 6458 13216 6695
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 13188 4758 13216 5646
rect 13176 4752 13228 4758
rect 13176 4694 13228 4700
rect 13280 4690 13308 6990
rect 13372 5166 13400 9710
rect 13464 7993 13492 11290
rect 13556 10130 13584 13466
rect 13740 13326 13768 14214
rect 13728 13320 13780 13326
rect 13728 13262 13780 13268
rect 13832 12434 13860 18294
rect 14200 18290 14228 18702
rect 14292 18426 14320 20454
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14660 20262 14688 20402
rect 14648 20256 14700 20262
rect 14646 20224 14648 20233
rect 14700 20224 14702 20233
rect 14646 20159 14702 20168
rect 14648 19780 14700 19786
rect 14648 19722 14700 19728
rect 14660 19514 14688 19722
rect 14648 19508 14700 19514
rect 14648 19450 14700 19456
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 14280 18420 14332 18426
rect 14280 18362 14332 18368
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 14292 15366 14320 16050
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14280 13184 14332 13190
rect 14280 13126 14332 13132
rect 14016 12850 14044 13126
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 14292 12646 14320 13126
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 13832 12406 14320 12434
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13648 11393 13676 11494
rect 13634 11384 13690 11393
rect 13634 11319 13690 11328
rect 13648 10810 13676 11319
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13832 10674 13860 12310
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 14096 11144 14148 11150
rect 14094 11112 14096 11121
rect 14148 11112 14150 11121
rect 14094 11047 14150 11056
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13636 10600 13688 10606
rect 13636 10542 13688 10548
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13542 8664 13598 8673
rect 13542 8599 13544 8608
rect 13596 8599 13598 8608
rect 13544 8570 13596 8576
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13450 7984 13506 7993
rect 13450 7919 13506 7928
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 6769 13492 7686
rect 13556 7426 13584 8230
rect 13648 7546 13676 10542
rect 13740 10130 13768 10610
rect 13924 10470 13952 10746
rect 14200 10470 14228 10950
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13740 9518 13768 9862
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13740 8242 13768 9454
rect 13832 8922 13860 10406
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14188 9172 14240 9178
rect 14188 9114 14240 9120
rect 14016 8974 14044 9114
rect 14200 9081 14228 9114
rect 14186 9072 14242 9081
rect 14186 9007 14242 9016
rect 14004 8968 14056 8974
rect 13832 8894 13952 8922
rect 14004 8910 14056 8916
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13832 8537 13860 8774
rect 13818 8528 13874 8537
rect 13818 8463 13874 8472
rect 13924 8430 13952 8894
rect 14292 8566 14320 12406
rect 14384 11898 14412 15642
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14384 10810 14412 11698
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14476 10146 14504 18566
rect 14660 15910 14688 19450
rect 14752 18970 14780 22200
rect 14740 18964 14792 18970
rect 14740 18906 14792 18912
rect 15304 18873 15332 22200
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15476 19848 15528 19854
rect 15382 19816 15438 19825
rect 15476 19790 15528 19796
rect 15568 19848 15620 19854
rect 15568 19790 15620 19796
rect 15382 19751 15438 19760
rect 15396 19446 15424 19751
rect 15384 19440 15436 19446
rect 15384 19382 15436 19388
rect 15488 19378 15516 19790
rect 15476 19372 15528 19378
rect 15476 19314 15528 19320
rect 15290 18864 15346 18873
rect 15290 18799 15346 18808
rect 15580 17785 15608 19790
rect 15566 17776 15622 17785
rect 15566 17711 15622 17720
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 14740 16448 14792 16454
rect 14844 16436 14872 17138
rect 14792 16408 14872 16436
rect 14740 16390 14792 16396
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14568 12646 14596 14418
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14568 11354 14596 12582
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14660 11150 14688 12786
rect 14752 12730 14780 16390
rect 15120 15450 15148 17478
rect 15476 15972 15528 15978
rect 15476 15914 15528 15920
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 14844 15422 15148 15450
rect 15212 15434 15240 15846
rect 15488 15434 15516 15914
rect 15200 15428 15252 15434
rect 14844 12850 14872 15422
rect 15200 15370 15252 15376
rect 15292 15428 15344 15434
rect 15292 15370 15344 15376
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 14924 14340 14976 14346
rect 14924 14282 14976 14288
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14752 12702 14872 12730
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14568 10266 14596 11086
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14476 10118 14596 10146
rect 14462 9752 14518 9761
rect 14462 9687 14518 9696
rect 14280 8560 14332 8566
rect 14280 8502 14332 8508
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 14292 8378 14320 8502
rect 14292 8350 14412 8378
rect 14280 8288 14332 8294
rect 13740 8214 13860 8242
rect 14280 8230 14332 8236
rect 13726 8120 13782 8129
rect 13726 8055 13728 8064
rect 13780 8055 13782 8064
rect 13728 8026 13780 8032
rect 13740 7818 13768 8026
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13832 7698 13860 8214
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 13740 7670 13860 7698
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13556 7398 13676 7426
rect 13542 7032 13598 7041
rect 13542 6967 13598 6976
rect 13556 6866 13584 6967
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13450 6760 13506 6769
rect 13450 6695 13506 6704
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 13556 6225 13584 6326
rect 13542 6216 13598 6225
rect 13542 6151 13598 6160
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 13464 5370 13492 6054
rect 13556 5778 13584 6151
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 13556 4826 13584 5170
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13280 4146 13308 4626
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13084 3392 13136 3398
rect 13084 3334 13136 3340
rect 13372 3126 13400 3470
rect 13464 3194 13492 4014
rect 13648 3942 13676 7398
rect 13740 6322 13768 7670
rect 14292 7478 14320 8230
rect 14384 7954 14412 8350
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 14476 7342 14504 9687
rect 14568 9518 14596 10118
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14568 8090 14596 9318
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14568 7546 14596 7686
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 13832 7206 13860 7278
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 14280 6724 14332 6730
rect 14280 6666 14332 6672
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13832 5914 13860 6598
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 13818 5808 13874 5817
rect 13740 4282 13768 5782
rect 13818 5743 13874 5752
rect 13832 5710 13860 5743
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13924 5273 13952 5306
rect 13910 5264 13966 5273
rect 13910 5199 13966 5208
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13832 3602 13860 4966
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14200 4282 14228 4422
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14292 4146 14320 6666
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14372 5092 14424 5098
rect 14372 5034 14424 5040
rect 14384 5001 14412 5034
rect 14476 5030 14504 6258
rect 14660 5166 14688 10950
rect 14752 6254 14780 11834
rect 14844 11778 14872 12702
rect 14936 12102 14964 14282
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 15028 13258 15056 13670
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 15120 13138 15148 15302
rect 15212 14822 15240 15370
rect 15304 15162 15332 15370
rect 15488 15314 15516 15370
rect 15672 15337 15700 20402
rect 15856 19174 15884 22200
rect 16304 20324 16356 20330
rect 16304 20266 16356 20272
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 16212 20256 16264 20262
rect 16212 20198 16264 20204
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15948 18970 15976 20198
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 16040 18766 16068 19246
rect 16028 18760 16080 18766
rect 16224 18748 16252 20198
rect 16316 19417 16344 20266
rect 16408 19718 16436 22200
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 16764 20392 16816 20398
rect 16764 20334 16816 20340
rect 16776 20233 16804 20334
rect 16762 20224 16818 20233
rect 16762 20159 16818 20168
rect 16960 19786 16988 22200
rect 17040 19848 17092 19854
rect 17040 19790 17092 19796
rect 17316 19848 17368 19854
rect 17316 19790 17368 19796
rect 16948 19780 17000 19786
rect 16948 19722 17000 19728
rect 16396 19712 16448 19718
rect 16396 19654 16448 19660
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 16302 19408 16358 19417
rect 16302 19343 16358 19352
rect 16304 18760 16356 18766
rect 16224 18720 16304 18748
rect 16028 18702 16080 18708
rect 16304 18702 16356 18708
rect 16486 18728 16542 18737
rect 15844 18624 15896 18630
rect 15844 18566 15896 18572
rect 15856 18290 15884 18566
rect 16040 18426 16068 18702
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15764 16590 15792 17070
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15764 15910 15792 16526
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15396 15286 15516 15314
rect 15658 15328 15714 15337
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15304 13433 15332 13942
rect 15290 13424 15346 13433
rect 15290 13359 15346 13368
rect 15028 13110 15148 13138
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14936 11898 14964 12038
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 14844 11750 14964 11778
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14844 11354 14872 11630
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14844 8480 14872 11086
rect 14936 10849 14964 11750
rect 15028 11014 15056 13110
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15212 11354 15240 11698
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 14922 10840 14978 10849
rect 14922 10775 14978 10784
rect 14936 10606 14964 10775
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 15212 10062 15240 10610
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 15120 9722 15148 9862
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 14922 9616 14978 9625
rect 14922 9551 14924 9560
rect 14976 9551 14978 9560
rect 14924 9522 14976 9528
rect 14936 9178 14964 9522
rect 15120 9518 15148 9549
rect 15108 9512 15160 9518
rect 15106 9480 15108 9489
rect 15160 9480 15162 9489
rect 15106 9415 15162 9424
rect 15120 9178 15148 9415
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 15212 8838 15240 9862
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15198 8664 15254 8673
rect 15198 8599 15200 8608
rect 15252 8599 15254 8608
rect 15200 8570 15252 8576
rect 15212 8514 15240 8570
rect 15120 8486 15240 8514
rect 14844 8452 15056 8480
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14844 7410 14872 8298
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 14936 7546 14964 7822
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14464 5024 14516 5030
rect 14370 4992 14426 5001
rect 14464 4966 14516 4972
rect 14370 4927 14426 4936
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14568 4010 14596 4422
rect 14660 4078 14688 5102
rect 14752 4690 14780 6190
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14556 4004 14608 4010
rect 14556 3946 14608 3952
rect 14844 3890 14872 7346
rect 15028 6866 15056 8452
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 14924 6724 14976 6730
rect 14924 6666 14976 6672
rect 14936 6390 14964 6666
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 14924 6384 14976 6390
rect 14924 6326 14976 6332
rect 14936 5370 14964 6326
rect 15028 6118 15056 6598
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 15028 5234 15056 6054
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 14660 3862 14872 3890
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 13372 2774 13400 3062
rect 13556 3058 13584 3334
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13820 2984 13872 2990
rect 14200 2961 14228 3130
rect 13820 2926 13872 2932
rect 14186 2952 14242 2961
rect 12268 2746 12388 2774
rect 13188 2746 13400 2774
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 12164 2440 12216 2446
rect 12164 2382 12216 2388
rect 12268 2106 12296 2746
rect 13188 2650 13216 2746
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13832 2446 13860 2926
rect 14186 2887 14242 2896
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 12532 2304 12584 2310
rect 12532 2246 12584 2252
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 12256 2100 12308 2106
rect 12256 2042 12308 2048
rect 11900 1414 12020 1442
rect 11992 800 12020 1414
rect 12544 800 12572 2246
rect 13096 800 13124 2246
rect 13556 1170 13584 2246
rect 13556 1142 13676 1170
rect 13648 800 13676 1142
rect 14200 800 14228 2246
rect 14660 2038 14688 3862
rect 14936 3777 14964 4626
rect 14922 3768 14978 3777
rect 14740 3732 14792 3738
rect 14922 3703 14978 3712
rect 14740 3674 14792 3680
rect 14648 2032 14700 2038
rect 14648 1974 14700 1980
rect 14752 800 14780 3674
rect 14832 3392 14884 3398
rect 14832 3334 14884 3340
rect 14844 3194 14872 3334
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 14936 3126 14964 3703
rect 14924 3120 14976 3126
rect 14924 3062 14976 3068
rect 15028 2774 15056 5170
rect 15120 4690 15148 8486
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 15212 6089 15240 8366
rect 15304 6474 15332 13359
rect 15396 9602 15424 15286
rect 15658 15263 15714 15272
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15672 13326 15700 13806
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15660 13320 15712 13326
rect 15856 13274 15884 18226
rect 16040 18222 16068 18362
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 16316 18154 16344 18702
rect 16486 18663 16488 18672
rect 16540 18663 16542 18672
rect 16670 18728 16726 18737
rect 16670 18663 16672 18672
rect 16488 18634 16540 18640
rect 16724 18663 16726 18672
rect 16672 18634 16724 18640
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 16488 18216 16540 18222
rect 16488 18158 16540 18164
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 16028 17876 16080 17882
rect 16028 17818 16080 17824
rect 16040 16998 16068 17818
rect 16500 17678 16528 18158
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 16040 16590 16068 16934
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 15936 16516 15988 16522
rect 15936 16458 15988 16464
rect 15660 13262 15712 13268
rect 15488 12918 15516 13262
rect 15764 13246 15884 13274
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15488 12306 15516 12854
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15488 11898 15516 12242
rect 15568 12164 15620 12170
rect 15568 12106 15620 12112
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15396 9574 15516 9602
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15396 8362 15424 8774
rect 15384 8356 15436 8362
rect 15384 8298 15436 8304
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15396 6730 15424 8026
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 15304 6446 15424 6474
rect 15290 6352 15346 6361
rect 15290 6287 15346 6296
rect 15304 6254 15332 6287
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15198 6080 15254 6089
rect 15198 6015 15254 6024
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 15212 5710 15240 5850
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15212 5370 15240 5510
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 15120 3602 15148 4014
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15212 3126 15240 4966
rect 15304 4826 15332 6190
rect 15396 5846 15424 6446
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15396 4554 15424 5306
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 15488 3670 15516 9574
rect 15580 8922 15608 12106
rect 15764 11830 15792 13246
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15752 11824 15804 11830
rect 15752 11766 15804 11772
rect 15764 11218 15792 11766
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 15672 9586 15700 11018
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15672 9110 15700 9522
rect 15764 9518 15792 10406
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15580 8894 15700 8922
rect 15568 8832 15620 8838
rect 15566 8800 15568 8809
rect 15620 8800 15622 8809
rect 15566 8735 15622 8744
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15580 7002 15608 7346
rect 15672 7206 15700 8894
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15672 4690 15700 5714
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15476 3664 15528 3670
rect 15476 3606 15528 3612
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 15304 3194 15332 3334
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15200 3120 15252 3126
rect 15200 3062 15252 3068
rect 14936 2746 15056 2774
rect 14936 2650 14964 2746
rect 14924 2644 14976 2650
rect 14924 2586 14976 2592
rect 15396 1714 15424 3470
rect 15488 2990 15516 3606
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15580 2514 15608 3470
rect 15672 3058 15700 4626
rect 15764 4486 15792 9114
rect 15856 7342 15884 13126
rect 15948 10130 15976 16458
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16408 15026 16436 15438
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 16408 14414 16436 14962
rect 16396 14408 16448 14414
rect 16396 14350 16448 14356
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 16856 13728 16908 13734
rect 16854 13696 16856 13705
rect 16908 13696 16910 13705
rect 16854 13631 16910 13640
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16028 13252 16080 13258
rect 16028 13194 16080 13200
rect 16040 12714 16068 13194
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 16028 12436 16080 12442
rect 16028 12378 16080 12384
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 15936 9988 15988 9994
rect 15936 9930 15988 9936
rect 15948 8634 15976 9930
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 15948 8344 15976 8570
rect 16040 8566 16068 12378
rect 16132 12374 16160 12786
rect 16120 12368 16172 12374
rect 16120 12310 16172 12316
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16132 11150 16160 11834
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 15948 8316 16068 8344
rect 15934 8256 15990 8265
rect 15934 8191 15990 8200
rect 15948 7750 15976 8191
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 15844 7336 15896 7342
rect 15844 7278 15896 7284
rect 15948 6934 15976 7686
rect 15936 6928 15988 6934
rect 15936 6870 15988 6876
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 15948 5914 15976 6258
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 16040 5778 16068 8316
rect 16132 6866 16160 11086
rect 16224 10606 16252 11086
rect 16316 10742 16344 13262
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16960 12170 16988 19450
rect 17052 19174 17080 19790
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 17040 18080 17092 18086
rect 17040 18022 17092 18028
rect 17052 16182 17080 18022
rect 17144 16561 17172 18566
rect 17328 16574 17356 19790
rect 17512 19417 17540 22200
rect 17592 20528 17644 20534
rect 17592 20470 17644 20476
rect 17604 19990 17632 20470
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17592 19984 17644 19990
rect 17592 19926 17644 19932
rect 17972 19825 18000 20198
rect 18064 20058 18092 22200
rect 18616 20602 18644 22200
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18696 20596 18748 20602
rect 18696 20538 18748 20544
rect 18708 20505 18736 20538
rect 18694 20496 18750 20505
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 18420 20460 18472 20466
rect 18694 20431 18750 20440
rect 18880 20460 18932 20466
rect 18420 20402 18472 20408
rect 18880 20402 18932 20408
rect 18156 20262 18184 20402
rect 18144 20256 18196 20262
rect 18144 20198 18196 20204
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 18234 19952 18290 19961
rect 18432 19922 18460 20402
rect 18786 20360 18842 20369
rect 18786 20295 18842 20304
rect 18696 20052 18748 20058
rect 18696 19994 18748 20000
rect 18602 19952 18658 19961
rect 18234 19887 18290 19896
rect 18420 19916 18472 19922
rect 18248 19854 18276 19887
rect 18602 19887 18658 19896
rect 18420 19858 18472 19864
rect 18236 19848 18288 19854
rect 17958 19816 18014 19825
rect 18236 19790 18288 19796
rect 17958 19751 18014 19760
rect 18420 19780 18472 19786
rect 18420 19722 18472 19728
rect 17498 19408 17554 19417
rect 17498 19343 17554 19352
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 17684 18624 17736 18630
rect 17684 18566 17736 18572
rect 17696 18154 17724 18566
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 17684 18148 17736 18154
rect 17684 18090 17736 18096
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 18064 17610 18092 18022
rect 18156 17882 18184 18158
rect 18144 17876 18196 17882
rect 18144 17818 18196 17824
rect 18052 17604 18104 17610
rect 18052 17546 18104 17552
rect 18064 16574 18092 17546
rect 17130 16552 17186 16561
rect 17328 16546 17448 16574
rect 17130 16487 17186 16496
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 17132 16176 17184 16182
rect 17132 16118 17184 16124
rect 17052 16017 17080 16118
rect 17038 16008 17094 16017
rect 17038 15943 17094 15952
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 17052 13258 17080 13670
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16946 12064 17002 12073
rect 16544 11996 16852 12005
rect 16946 11999 17002 12008
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16960 11898 16988 11999
rect 16948 11892 17000 11898
rect 16948 11834 17000 11840
rect 17052 11830 17080 12174
rect 17040 11824 17092 11830
rect 17040 11766 17092 11772
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 16960 11286 16988 11630
rect 17052 11354 17080 11766
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 16948 11280 17000 11286
rect 16948 11222 17000 11228
rect 17038 11112 17094 11121
rect 17038 11047 17040 11056
rect 17092 11047 17094 11056
rect 17040 11018 17092 11024
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16304 10736 16356 10742
rect 16304 10678 16356 10684
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16224 9178 16252 10542
rect 16592 9994 16620 10542
rect 16684 10198 16712 10610
rect 16672 10192 16724 10198
rect 16672 10134 16724 10140
rect 16946 10160 17002 10169
rect 16946 10095 17002 10104
rect 16960 10062 16988 10095
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16580 9988 16632 9994
rect 16580 9930 16632 9936
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 17052 9722 17080 9862
rect 17040 9716 17092 9722
rect 17040 9658 17092 9664
rect 16946 9616 17002 9625
rect 17144 9586 17172 16118
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17236 11762 17264 12922
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17328 11098 17356 14962
rect 17236 11070 17356 11098
rect 16946 9551 17002 9560
rect 17132 9580 17184 9586
rect 16960 9518 16988 9551
rect 17132 9522 17184 9528
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16580 9512 16632 9518
rect 16580 9454 16632 9460
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16316 9058 16344 9318
rect 16224 9030 16344 9058
rect 16224 8265 16252 9030
rect 16408 8906 16436 9454
rect 16592 9042 16620 9454
rect 16960 9382 16988 9454
rect 17132 9444 17184 9450
rect 17132 9386 17184 9392
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 16304 8832 16356 8838
rect 16948 8832 17000 8838
rect 16356 8780 16436 8786
rect 16304 8774 16436 8780
rect 16948 8774 17000 8780
rect 16316 8758 16436 8774
rect 16210 8256 16266 8265
rect 16210 8191 16266 8200
rect 16224 8022 16252 8053
rect 16212 8016 16264 8022
rect 16408 7970 16436 8758
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 16960 8634 16988 8774
rect 17052 8634 17080 9318
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 16856 8560 16908 8566
rect 16856 8502 16908 8508
rect 16868 8090 16896 8502
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16264 7964 16436 7970
rect 16212 7958 16436 7964
rect 16224 7942 16436 7958
rect 16224 7206 16252 7942
rect 17144 7818 17172 9386
rect 17236 8430 17264 11070
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17328 10810 17356 10950
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17314 10704 17370 10713
rect 17314 10639 17370 10648
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17132 7812 17184 7818
rect 17132 7754 17184 7760
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16316 7546 16344 7686
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16408 7478 16436 7686
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 16396 7472 16448 7478
rect 16396 7414 16448 7420
rect 17328 7410 17356 10639
rect 17420 10266 17448 16546
rect 17972 16546 18092 16574
rect 17682 15056 17738 15065
rect 17682 14991 17738 15000
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17604 14006 17632 14214
rect 17592 14000 17644 14006
rect 17592 13942 17644 13948
rect 17500 13388 17552 13394
rect 17500 13330 17552 13336
rect 17512 10674 17540 13330
rect 17604 12306 17632 13942
rect 17592 12300 17644 12306
rect 17592 12242 17644 12248
rect 17592 12164 17644 12170
rect 17592 12106 17644 12112
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17408 10260 17460 10266
rect 17408 10202 17460 10208
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17420 9081 17448 9930
rect 17406 9072 17462 9081
rect 17406 9007 17462 9016
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16960 7002 16988 7278
rect 16948 6996 17000 7002
rect 16948 6938 17000 6944
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 16118 6760 16174 6769
rect 16118 6695 16174 6704
rect 16304 6724 16356 6730
rect 16132 6322 16160 6695
rect 16304 6666 16356 6672
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 16132 5574 16160 6258
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 15842 5400 15898 5409
rect 15842 5335 15844 5344
rect 15896 5335 15898 5344
rect 15844 5306 15896 5312
rect 15856 4690 15884 5306
rect 16132 5030 16160 5510
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15856 4185 15884 4626
rect 16028 4548 16080 4554
rect 16028 4490 16080 4496
rect 16040 4282 16068 4490
rect 16028 4276 16080 4282
rect 16028 4218 16080 4224
rect 15842 4176 15898 4185
rect 15842 4111 15898 4120
rect 15750 3496 15806 3505
rect 15750 3431 15806 3440
rect 15764 3398 15792 3431
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 15764 2961 15792 3334
rect 15856 3058 15884 4111
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15750 2952 15806 2961
rect 15750 2887 15806 2896
rect 15844 2576 15896 2582
rect 15844 2518 15896 2524
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15752 2372 15804 2378
rect 15752 2314 15804 2320
rect 15476 2304 15528 2310
rect 15568 2304 15620 2310
rect 15528 2252 15568 2258
rect 15476 2246 15620 2252
rect 15488 2230 15608 2246
rect 15488 1970 15516 2230
rect 15764 2038 15792 2314
rect 15752 2032 15804 2038
rect 15752 1974 15804 1980
rect 15476 1964 15528 1970
rect 15476 1906 15528 1912
rect 15304 1686 15424 1714
rect 15304 800 15332 1686
rect 15856 800 15884 2518
rect 16040 2514 16068 4218
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16132 3602 16160 3878
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 16224 2650 16252 5714
rect 16316 4162 16344 6666
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 16960 6338 16988 6598
rect 17038 6488 17094 6497
rect 17038 6423 17094 6432
rect 16868 6310 16988 6338
rect 17052 6322 17080 6423
rect 17040 6316 17092 6322
rect 16764 6180 16816 6186
rect 16764 6122 16816 6128
rect 16408 5642 16528 5658
rect 16408 5636 16540 5642
rect 16408 5630 16488 5636
rect 16408 5370 16436 5630
rect 16488 5578 16540 5584
rect 16776 5574 16804 6122
rect 16868 5794 16896 6310
rect 17040 6258 17092 6264
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 16960 5914 16988 6190
rect 17132 6112 17184 6118
rect 17132 6054 17184 6060
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 17052 5817 17080 5850
rect 17038 5808 17094 5817
rect 16868 5766 16988 5794
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16776 5098 16804 5306
rect 16764 5092 16816 5098
rect 16764 5034 16816 5040
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 16960 4264 16988 5766
rect 17038 5743 17094 5752
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 17052 4622 17080 5510
rect 17144 5302 17172 6054
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 17236 5166 17264 6190
rect 17420 6066 17448 9007
rect 17512 7954 17540 10406
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 17512 6934 17540 7890
rect 17500 6928 17552 6934
rect 17500 6870 17552 6876
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17512 6100 17540 6394
rect 17604 6254 17632 12106
rect 17696 10810 17724 14991
rect 17776 13728 17828 13734
rect 17776 13670 17828 13676
rect 17788 12434 17816 13670
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17880 13433 17908 13466
rect 17866 13424 17922 13433
rect 17866 13359 17922 13368
rect 17788 12406 17908 12434
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 17696 9178 17724 9522
rect 17684 9172 17736 9178
rect 17684 9114 17736 9120
rect 17788 7834 17816 12242
rect 17880 12050 17908 12406
rect 17972 12170 18000 16546
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 18064 14822 18092 15302
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 18156 13138 18184 17818
rect 18340 16590 18368 19314
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 18236 16516 18288 16522
rect 18236 16458 18288 16464
rect 18248 16402 18276 16458
rect 18248 16374 18368 16402
rect 18236 13456 18288 13462
rect 18234 13424 18236 13433
rect 18288 13424 18290 13433
rect 18234 13359 18290 13368
rect 18156 13110 18276 13138
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 18064 12238 18092 12718
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 17960 12164 18012 12170
rect 17960 12106 18012 12112
rect 17880 12022 18000 12050
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 17696 7806 17816 7834
rect 17696 6866 17724 7806
rect 17776 7744 17828 7750
rect 17776 7686 17828 7692
rect 17788 7546 17816 7686
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17776 7404 17828 7410
rect 17776 7346 17828 7352
rect 17684 6860 17736 6866
rect 17684 6802 17736 6808
rect 17788 6338 17816 7346
rect 17696 6310 17816 6338
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17512 6072 17632 6100
rect 17328 6038 17448 6066
rect 17328 5846 17356 6038
rect 17406 5944 17462 5953
rect 17406 5879 17462 5888
rect 17316 5840 17368 5846
rect 17316 5782 17368 5788
rect 17420 5710 17448 5879
rect 17498 5808 17554 5817
rect 17604 5778 17632 6072
rect 17498 5743 17500 5752
rect 17552 5743 17554 5752
rect 17592 5772 17644 5778
rect 17500 5714 17552 5720
rect 17592 5714 17644 5720
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17420 5234 17448 5646
rect 17696 5574 17724 6310
rect 17776 6248 17828 6254
rect 17774 6216 17776 6225
rect 17828 6216 17830 6225
rect 17774 6151 17830 6160
rect 17776 5840 17828 5846
rect 17776 5782 17828 5788
rect 17500 5568 17552 5574
rect 17500 5510 17552 5516
rect 17684 5568 17736 5574
rect 17684 5510 17736 5516
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 16868 4236 16988 4264
rect 16488 4208 16540 4214
rect 16316 4134 16436 4162
rect 16488 4150 16540 4156
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 16316 3466 16344 4014
rect 16304 3460 16356 3466
rect 16304 3402 16356 3408
rect 16408 3398 16436 4134
rect 16500 3534 16528 4150
rect 16868 4049 16896 4236
rect 16948 4072 17000 4078
rect 16854 4040 16910 4049
rect 16948 4014 17000 4020
rect 16854 3975 16910 3984
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 16960 3058 16988 4014
rect 17144 3534 17172 4966
rect 17236 3738 17264 5102
rect 17316 5024 17368 5030
rect 17316 4966 17368 4972
rect 17328 4146 17356 4966
rect 17420 4214 17448 5170
rect 17512 4706 17540 5510
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17696 4826 17724 5170
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 17512 4678 17724 4706
rect 17500 4548 17552 4554
rect 17500 4490 17552 4496
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 17236 2990 17264 3674
rect 17224 2984 17276 2990
rect 17224 2926 17276 2932
rect 16948 2916 17000 2922
rect 16948 2858 17000 2864
rect 16396 2848 16448 2854
rect 16396 2790 16448 2796
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 15948 2106 15976 2382
rect 15936 2100 15988 2106
rect 15936 2042 15988 2048
rect 16408 800 16436 2790
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 16960 800 16988 2858
rect 17236 2774 17264 2926
rect 17052 2746 17264 2774
rect 17052 2310 17080 2746
rect 17420 2582 17448 4150
rect 17512 3058 17540 4490
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17408 2576 17460 2582
rect 17408 2518 17460 2524
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 17512 800 17540 2790
rect 17696 2774 17724 4678
rect 17788 4282 17816 5782
rect 17880 5166 17908 11834
rect 17972 11234 18000 12022
rect 18064 11830 18092 12174
rect 18144 12164 18196 12170
rect 18144 12106 18196 12112
rect 18052 11824 18104 11830
rect 18052 11766 18104 11772
rect 18156 11558 18184 12106
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 17972 11206 18092 11234
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17972 10674 18000 11018
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 18064 10470 18092 11206
rect 18142 10840 18198 10849
rect 18142 10775 18144 10784
rect 18196 10775 18198 10784
rect 18144 10746 18196 10752
rect 18144 10600 18196 10606
rect 18248 10588 18276 13110
rect 18196 10560 18276 10588
rect 18144 10542 18196 10548
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 17958 10160 18014 10169
rect 17958 10095 17960 10104
rect 18012 10095 18014 10104
rect 17960 10066 18012 10072
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 17958 9480 18014 9489
rect 18064 9450 18092 9862
rect 18156 9722 18184 9862
rect 18144 9716 18196 9722
rect 18144 9658 18196 9664
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 17958 9415 18014 9424
rect 18052 9444 18104 9450
rect 17972 9110 18000 9415
rect 18052 9386 18104 9392
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 17972 8634 18000 9046
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 17960 8016 18012 8022
rect 17960 7958 18012 7964
rect 17972 7342 18000 7958
rect 17960 7336 18012 7342
rect 18064 7313 18092 8910
rect 18156 8634 18184 9454
rect 18248 9110 18276 10560
rect 18340 10130 18368 16374
rect 18432 11354 18460 19722
rect 18616 17762 18644 19887
rect 18708 19378 18736 19994
rect 18800 19854 18828 20295
rect 18788 19848 18840 19854
rect 18788 19790 18840 19796
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18694 19272 18750 19281
rect 18694 19207 18750 19216
rect 18708 18970 18736 19207
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 18892 18850 18920 20402
rect 19168 20244 19196 22200
rect 19720 21026 19748 22200
rect 19076 20216 19196 20244
rect 19536 20998 19748 21026
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 18800 18822 18920 18850
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18708 18358 18736 18702
rect 18800 18426 18828 18822
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18788 18420 18840 18426
rect 18788 18362 18840 18368
rect 18696 18352 18748 18358
rect 18696 18294 18748 18300
rect 18616 17734 18736 17762
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18616 17066 18644 17546
rect 18604 17060 18656 17066
rect 18604 17002 18656 17008
rect 18708 16998 18736 17734
rect 18788 17536 18840 17542
rect 18788 17478 18840 17484
rect 18800 17202 18828 17478
rect 18788 17196 18840 17202
rect 18788 17138 18840 17144
rect 18696 16992 18748 16998
rect 18696 16934 18748 16940
rect 18602 16552 18658 16561
rect 18602 16487 18658 16496
rect 18512 16040 18564 16046
rect 18512 15982 18564 15988
rect 18524 15502 18552 15982
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18418 11248 18474 11257
rect 18418 11183 18474 11192
rect 18432 11150 18460 11183
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18420 10804 18472 10810
rect 18420 10746 18472 10752
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18236 9104 18288 9110
rect 18236 9046 18288 9052
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18248 8650 18276 8910
rect 18144 8628 18196 8634
rect 18248 8622 18368 8650
rect 18432 8634 18460 10746
rect 18524 9042 18552 15302
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18144 8570 18196 8576
rect 18236 8560 18288 8566
rect 18236 8502 18288 8508
rect 18144 7336 18196 7342
rect 17960 7278 18012 7284
rect 18050 7304 18106 7313
rect 17972 6866 18000 7278
rect 18144 7278 18196 7284
rect 18050 7239 18106 7248
rect 18156 7177 18184 7278
rect 18142 7168 18198 7177
rect 18142 7103 18198 7112
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 18064 6186 18092 6734
rect 18248 6390 18276 8502
rect 18340 8498 18368 8622
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18328 8492 18380 8498
rect 18328 8434 18380 8440
rect 18524 8362 18552 8978
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 18328 8288 18380 8294
rect 18328 8230 18380 8236
rect 18340 7585 18368 8230
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18326 7576 18382 7585
rect 18432 7546 18460 7686
rect 18326 7511 18382 7520
rect 18420 7540 18472 7546
rect 18340 7410 18368 7511
rect 18420 7482 18472 7488
rect 18328 7404 18380 7410
rect 18328 7346 18380 7352
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 18236 6384 18288 6390
rect 18236 6326 18288 6332
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 18052 6180 18104 6186
rect 18052 6122 18104 6128
rect 17972 5817 18000 6122
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 18156 5914 18184 6054
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 17958 5808 18014 5817
rect 17958 5743 18014 5752
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17958 5128 18014 5137
rect 17958 5063 18014 5072
rect 18052 5092 18104 5098
rect 17972 4758 18000 5063
rect 18052 5034 18104 5040
rect 17960 4752 18012 4758
rect 17960 4694 18012 4700
rect 17960 4616 18012 4622
rect 17958 4584 17960 4593
rect 18012 4584 18014 4593
rect 17958 4519 18014 4528
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 17880 3097 17908 3946
rect 17958 3768 18014 3777
rect 17958 3703 18014 3712
rect 17972 3534 18000 3703
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17866 3088 17922 3097
rect 17866 3023 17868 3032
rect 17920 3023 17922 3032
rect 17868 2994 17920 3000
rect 17696 2746 17816 2774
rect 17788 2514 17816 2746
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 18064 800 18092 5034
rect 18156 5001 18184 5714
rect 18142 4992 18198 5001
rect 18142 4927 18198 4936
rect 18156 4049 18184 4927
rect 18142 4040 18198 4049
rect 18142 3975 18198 3984
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18248 3097 18276 3878
rect 18340 3369 18368 7142
rect 18524 7002 18552 7686
rect 18616 7206 18644 16487
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18708 15366 18736 16390
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18800 14090 18828 17138
rect 18708 14062 18828 14090
rect 18708 12918 18736 14062
rect 18786 13968 18842 13977
rect 18786 13903 18842 13912
rect 18800 13462 18828 13903
rect 18892 13841 18920 18702
rect 18984 17338 19012 19450
rect 19076 19242 19104 20216
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 19064 19236 19116 19242
rect 19064 19178 19116 19184
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 19536 18902 19564 20998
rect 19614 20904 19670 20913
rect 19614 20839 19670 20848
rect 19524 18896 19576 18902
rect 19524 18838 19576 18844
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 19628 17814 19656 20839
rect 20272 20534 20300 22200
rect 20534 21312 20590 21321
rect 20534 21247 20590 21256
rect 20260 20528 20312 20534
rect 20260 20470 20312 20476
rect 20168 20324 20220 20330
rect 20168 20266 20220 20272
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19708 19780 19760 19786
rect 19708 19722 19760 19728
rect 19720 18426 19748 19722
rect 19800 19372 19852 19378
rect 19800 19314 19852 19320
rect 19812 18630 19840 19314
rect 19996 18698 20024 20198
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19800 18624 19852 18630
rect 19800 18566 19852 18572
rect 20076 18624 20128 18630
rect 20076 18566 20128 18572
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 19720 18170 19748 18362
rect 19720 18142 19840 18170
rect 19616 17808 19668 17814
rect 19616 17750 19668 17756
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 18972 16992 19024 16998
rect 18972 16934 19024 16940
rect 18984 16522 19012 16934
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 19536 16794 19564 17614
rect 19708 17264 19760 17270
rect 19708 17206 19760 17212
rect 19614 16824 19670 16833
rect 19524 16788 19576 16794
rect 19614 16759 19670 16768
rect 19524 16730 19576 16736
rect 18972 16516 19024 16522
rect 18972 16458 19024 16464
rect 19156 16448 19208 16454
rect 19156 16390 19208 16396
rect 19168 15994 19196 16390
rect 18984 15966 19196 15994
rect 18878 13832 18934 13841
rect 18878 13767 18934 13776
rect 18788 13456 18840 13462
rect 18788 13398 18840 13404
rect 18696 12912 18748 12918
rect 18696 12854 18748 12860
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18708 11898 18736 12582
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18694 11792 18750 11801
rect 18694 11727 18750 11736
rect 18708 11218 18736 11727
rect 18696 11212 18748 11218
rect 18696 11154 18748 11160
rect 18800 10713 18828 12038
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18786 10704 18842 10713
rect 18696 10668 18748 10674
rect 18786 10639 18842 10648
rect 18696 10610 18748 10616
rect 18708 10130 18736 10610
rect 18786 10568 18842 10577
rect 18786 10503 18842 10512
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18694 9888 18750 9897
rect 18694 9823 18750 9832
rect 18708 8566 18736 9823
rect 18800 9178 18828 10503
rect 18892 9738 18920 10950
rect 18984 10606 19012 15966
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19536 14482 19564 16730
rect 19524 14476 19576 14482
rect 19524 14418 19576 14424
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19352 14074 19380 14214
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 19076 12238 19104 13942
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19444 13818 19472 13874
rect 19444 13790 19564 13818
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 19064 12232 19116 12238
rect 19064 12174 19116 12180
rect 19536 12102 19564 13790
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 18972 10464 19024 10470
rect 18970 10432 18972 10441
rect 19024 10432 19026 10441
rect 18970 10367 19026 10376
rect 18892 9710 19012 9738
rect 18878 9616 18934 9625
rect 18878 9551 18934 9560
rect 18892 9518 18920 9551
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18984 9042 19012 9710
rect 18972 9036 19024 9042
rect 18972 8978 19024 8984
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18696 8560 18748 8566
rect 18696 8502 18748 8508
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18694 8392 18750 8401
rect 18694 8327 18750 8336
rect 18708 7954 18736 8327
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18694 7848 18750 7857
rect 18694 7783 18750 7792
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18708 6914 18736 7783
rect 18616 6886 18736 6914
rect 18616 6662 18644 6886
rect 18604 6656 18656 6662
rect 18604 6598 18656 6604
rect 18418 6080 18474 6089
rect 18418 6015 18474 6024
rect 18432 5778 18460 6015
rect 18420 5772 18472 5778
rect 18420 5714 18472 5720
rect 18432 5137 18460 5714
rect 18512 5704 18564 5710
rect 18512 5646 18564 5652
rect 18418 5128 18474 5137
rect 18418 5063 18474 5072
rect 18326 3360 18382 3369
rect 18326 3295 18382 3304
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 18234 3088 18290 3097
rect 18234 3023 18290 3032
rect 18340 2774 18368 3130
rect 18340 2746 18460 2774
rect 18432 2650 18460 2746
rect 18420 2644 18472 2650
rect 18420 2586 18472 2592
rect 18524 2446 18552 5646
rect 18616 4321 18644 6598
rect 18800 6458 18828 8434
rect 18892 6769 18920 8774
rect 18984 7993 19012 8978
rect 18970 7984 19026 7993
rect 18970 7919 19026 7928
rect 18878 6760 18934 6769
rect 18878 6695 18934 6704
rect 18984 6610 19012 7919
rect 18892 6582 19012 6610
rect 18788 6452 18840 6458
rect 18788 6394 18840 6400
rect 18892 5710 18920 6582
rect 18972 6452 19024 6458
rect 18972 6394 19024 6400
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18880 5568 18932 5574
rect 18880 5510 18932 5516
rect 18892 5370 18920 5510
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 18880 5160 18932 5166
rect 18694 5128 18750 5137
rect 18880 5102 18932 5108
rect 18694 5063 18750 5072
rect 18602 4312 18658 4321
rect 18602 4247 18658 4256
rect 18616 3194 18644 4247
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18604 2916 18656 2922
rect 18604 2858 18656 2864
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18616 800 18644 2858
rect 18708 2310 18736 5063
rect 18892 4690 18920 5102
rect 18880 4684 18932 4690
rect 18880 4626 18932 4632
rect 18984 4162 19012 6394
rect 19076 5846 19104 12038
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 19352 10810 19380 10950
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19524 10532 19576 10538
rect 19524 10474 19576 10480
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19536 10062 19564 10474
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 19340 9512 19392 9518
rect 19340 9454 19392 9460
rect 19352 9382 19380 9454
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19444 8344 19472 9114
rect 19524 8900 19576 8906
rect 19524 8842 19576 8848
rect 19536 8498 19564 8842
rect 19628 8634 19656 16759
rect 19720 16522 19748 17206
rect 19708 16516 19760 16522
rect 19708 16458 19760 16464
rect 19720 15366 19748 16458
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19720 14958 19748 15302
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 19720 14414 19748 14894
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19708 12844 19760 12850
rect 19708 12786 19760 12792
rect 19720 11558 19748 12786
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19812 11218 19840 18142
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 19996 16522 20024 17138
rect 19984 16516 20036 16522
rect 19984 16458 20036 16464
rect 20088 16454 20116 18566
rect 20180 17202 20208 20266
rect 20548 19514 20576 21247
rect 20824 20466 20852 22200
rect 21376 20602 21404 22200
rect 21364 20596 21416 20602
rect 21364 20538 21416 20544
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 21100 20058 21128 20402
rect 21364 20392 21416 20398
rect 21364 20334 21416 20340
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 21376 19922 21404 20334
rect 21364 19916 21416 19922
rect 21364 19858 21416 19864
rect 20536 19508 20588 19514
rect 20536 19450 20588 19456
rect 20548 19378 20576 19450
rect 21376 19446 21404 19858
rect 20628 19440 20680 19446
rect 20628 19382 20680 19388
rect 21364 19440 21416 19446
rect 21364 19382 21416 19388
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20260 19304 20312 19310
rect 20260 19246 20312 19252
rect 20168 17196 20220 17202
rect 20168 17138 20220 17144
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 20168 16448 20220 16454
rect 20168 16390 20220 16396
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 19982 15600 20038 15609
rect 19982 15535 20038 15544
rect 19892 15360 19944 15366
rect 19890 15328 19892 15337
rect 19944 15328 19946 15337
rect 19890 15263 19946 15272
rect 19892 14272 19944 14278
rect 19892 14214 19944 14220
rect 19904 13297 19932 14214
rect 19890 13288 19946 13297
rect 19890 13223 19946 13232
rect 19892 12640 19944 12646
rect 19892 12582 19944 12588
rect 19904 11694 19932 12582
rect 19892 11688 19944 11694
rect 19892 11630 19944 11636
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 19708 11076 19760 11082
rect 19708 11018 19760 11024
rect 19720 9178 19748 11018
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 19812 10742 19840 10950
rect 19800 10736 19852 10742
rect 19800 10678 19852 10684
rect 19904 10146 19932 11630
rect 19812 10118 19932 10146
rect 19708 9172 19760 9178
rect 19708 9114 19760 9120
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19444 8316 19564 8344
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19536 7936 19564 8316
rect 19444 7908 19564 7936
rect 19444 7256 19472 7908
rect 19524 7812 19576 7818
rect 19524 7754 19576 7760
rect 19536 7410 19564 7754
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19616 7336 19668 7342
rect 19614 7304 19616 7313
rect 19668 7304 19670 7313
rect 19444 7228 19564 7256
rect 19614 7239 19670 7248
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19246 6896 19302 6905
rect 19536 6866 19564 7228
rect 19246 6831 19302 6840
rect 19340 6860 19392 6866
rect 19260 6458 19288 6831
rect 19340 6802 19392 6808
rect 19524 6860 19576 6866
rect 19524 6802 19576 6808
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19352 6118 19380 6802
rect 19524 6384 19576 6390
rect 19524 6326 19576 6332
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 19064 5840 19116 5846
rect 19064 5782 19116 5788
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 18892 4134 19196 4162
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18800 3505 18828 3878
rect 18786 3496 18842 3505
rect 18786 3431 18842 3440
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18800 2496 18828 3334
rect 18892 2650 18920 4134
rect 19168 4078 19196 4134
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 19156 4072 19208 4078
rect 19156 4014 19208 4020
rect 18970 3632 19026 3641
rect 18970 3567 19026 3576
rect 18880 2644 18932 2650
rect 18880 2586 18932 2592
rect 18800 2468 18920 2496
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 18892 2009 18920 2468
rect 18878 2000 18934 2009
rect 18878 1935 18934 1944
rect 18984 1850 19012 3567
rect 19076 3058 19104 4014
rect 19536 3942 19564 6326
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19616 6248 19668 6254
rect 19616 6190 19668 6196
rect 19628 4826 19656 6190
rect 19720 5273 19748 6258
rect 19812 5778 19840 10118
rect 19892 9988 19944 9994
rect 19892 9930 19944 9936
rect 19904 9586 19932 9930
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19996 9382 20024 15535
rect 20088 15094 20116 15846
rect 20180 15178 20208 16390
rect 20272 15366 20300 19246
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 20364 18766 20392 19110
rect 20640 18834 20668 19382
rect 21086 18864 21142 18873
rect 20628 18828 20680 18834
rect 21086 18799 21142 18808
rect 20628 18770 20680 18776
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20180 15150 20300 15178
rect 20076 15088 20128 15094
rect 20076 15030 20128 15036
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 20088 10674 20116 14418
rect 20168 14340 20220 14346
rect 20168 14282 20220 14288
rect 20180 13938 20208 14282
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20168 12912 20220 12918
rect 20168 12854 20220 12860
rect 20180 11082 20208 12854
rect 20168 11076 20220 11082
rect 20168 11018 20220 11024
rect 20076 10668 20128 10674
rect 20076 10610 20128 10616
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19890 8528 19946 8537
rect 19890 8463 19946 8472
rect 19984 8492 20036 8498
rect 19904 6254 19932 8463
rect 19984 8434 20036 8440
rect 19996 6390 20024 8434
rect 20180 7886 20208 10406
rect 20272 10146 20300 15150
rect 20364 11218 20392 18702
rect 20640 18358 20668 18770
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20628 18352 20680 18358
rect 20442 18320 20498 18329
rect 20628 18294 20680 18300
rect 20442 18255 20498 18264
rect 20456 16250 20484 18255
rect 20640 17678 20668 18294
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 20640 17218 20668 17614
rect 20548 17202 20668 17218
rect 20536 17196 20668 17202
rect 20588 17190 20668 17196
rect 20536 17138 20588 17144
rect 20534 17096 20590 17105
rect 20534 17031 20590 17040
rect 20444 16244 20496 16250
rect 20444 16186 20496 16192
rect 20548 12458 20576 17031
rect 20732 16289 20760 18702
rect 20902 17640 20958 17649
rect 20902 17575 20958 17584
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20718 16280 20774 16289
rect 20718 16215 20774 16224
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20626 14784 20682 14793
rect 20626 14719 20682 14728
rect 20640 13530 20668 14719
rect 20628 13524 20680 13530
rect 20628 13466 20680 13472
rect 20456 12442 20576 12458
rect 20444 12436 20576 12442
rect 20496 12430 20576 12436
rect 20444 12378 20496 12384
rect 20456 12347 20484 12378
rect 20352 11212 20404 11218
rect 20352 11154 20404 11160
rect 20364 10538 20392 11154
rect 20626 11112 20682 11121
rect 20536 11076 20588 11082
rect 20626 11047 20682 11056
rect 20536 11018 20588 11024
rect 20444 10600 20496 10606
rect 20444 10542 20496 10548
rect 20352 10532 20404 10538
rect 20352 10474 20404 10480
rect 20272 10118 20392 10146
rect 20260 10056 20312 10062
rect 20258 10024 20260 10033
rect 20312 10024 20314 10033
rect 20258 9959 20314 9968
rect 20260 9648 20312 9654
rect 20260 9590 20312 9596
rect 20272 9330 20300 9590
rect 20364 9450 20392 10118
rect 20352 9444 20404 9450
rect 20352 9386 20404 9392
rect 20272 9302 20392 9330
rect 20258 8664 20314 8673
rect 20258 8599 20260 8608
rect 20312 8599 20314 8608
rect 20260 8570 20312 8576
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 19984 6384 20036 6390
rect 19984 6326 20036 6332
rect 19892 6248 19944 6254
rect 19892 6190 19944 6196
rect 19892 6112 19944 6118
rect 19892 6054 19944 6060
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 19904 5710 19932 6054
rect 19984 5840 20036 5846
rect 19984 5782 20036 5788
rect 19892 5704 19944 5710
rect 19892 5646 19944 5652
rect 19706 5264 19762 5273
rect 19706 5199 19762 5208
rect 19996 5166 20024 5782
rect 19800 5160 19852 5166
rect 19800 5102 19852 5108
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 19616 4208 19668 4214
rect 19616 4150 19668 4156
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19352 3058 19380 3334
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19352 2961 19380 2994
rect 19536 2990 19564 3878
rect 19628 3738 19656 4150
rect 19812 4010 19840 5102
rect 19890 4176 19946 4185
rect 19890 4111 19946 4120
rect 19800 4004 19852 4010
rect 19800 3946 19852 3952
rect 19616 3732 19668 3738
rect 19616 3674 19668 3680
rect 19524 2984 19576 2990
rect 19338 2952 19394 2961
rect 19524 2926 19576 2932
rect 19338 2887 19394 2896
rect 19904 2774 19932 4111
rect 19984 4072 20036 4078
rect 19982 4040 19984 4049
rect 20036 4040 20038 4049
rect 19982 3975 20038 3984
rect 20088 3466 20116 6734
rect 20364 6662 20392 9302
rect 20456 6866 20484 10542
rect 20548 9722 20576 11018
rect 20640 10810 20668 11047
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20444 6860 20496 6866
rect 20444 6802 20496 6808
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 20260 5568 20312 5574
rect 20166 5536 20222 5545
rect 20260 5510 20312 5516
rect 20166 5471 20222 5480
rect 20180 4826 20208 5471
rect 20272 5302 20300 5510
rect 20260 5296 20312 5302
rect 20260 5238 20312 5244
rect 20364 5148 20392 6598
rect 20456 5166 20484 6802
rect 20536 5568 20588 5574
rect 20536 5510 20588 5516
rect 20548 5370 20576 5510
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20272 5120 20392 5148
rect 20444 5160 20496 5166
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20272 4729 20300 5120
rect 20444 5102 20496 5108
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20258 4720 20314 4729
rect 20258 4655 20260 4664
rect 20312 4655 20314 4664
rect 20260 4626 20312 4632
rect 20364 4146 20392 4966
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20352 4004 20404 4010
rect 20352 3946 20404 3952
rect 20260 3664 20312 3670
rect 20260 3606 20312 3612
rect 20076 3460 20128 3466
rect 20076 3402 20128 3408
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19904 2746 20024 2774
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 19996 2650 20024 2746
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 19708 2576 19760 2582
rect 19154 2544 19210 2553
rect 19708 2518 19760 2524
rect 19154 2479 19210 2488
rect 19168 2378 19196 2479
rect 19156 2372 19208 2378
rect 19156 2314 19208 2320
rect 18984 1822 19196 1850
rect 19168 800 19196 1822
rect 19720 800 19748 2518
rect 20272 800 20300 3606
rect 20364 1737 20392 3946
rect 20456 3058 20484 5102
rect 20640 4593 20668 10610
rect 20732 7954 20760 16050
rect 20824 9926 20852 16526
rect 20916 16250 20944 17575
rect 21100 16454 21128 18799
rect 21180 18692 21232 18698
rect 21180 18634 21232 18640
rect 21192 16998 21220 18634
rect 21456 18080 21508 18086
rect 21456 18022 21508 18028
rect 21468 17610 21496 18022
rect 21456 17604 21508 17610
rect 21456 17546 21508 17552
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 20996 16040 21048 16046
rect 20996 15982 21048 15988
rect 21362 16008 21418 16017
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 20916 11898 20944 13262
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 20812 9920 20864 9926
rect 20812 9862 20864 9868
rect 20812 8968 20864 8974
rect 20812 8910 20864 8916
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20824 7886 20852 8910
rect 20904 8832 20956 8838
rect 20904 8774 20956 8780
rect 21008 8786 21036 15982
rect 21362 15943 21418 15952
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21284 15502 21312 15846
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 21088 15428 21140 15434
rect 21088 15370 21140 15376
rect 21100 14822 21128 15370
rect 21088 14816 21140 14822
rect 21088 14758 21140 14764
rect 21284 14414 21312 15438
rect 21272 14408 21324 14414
rect 21178 14376 21234 14385
rect 21088 14340 21140 14346
rect 21272 14350 21324 14356
rect 21178 14311 21234 14320
rect 21088 14282 21140 14288
rect 21100 11558 21128 14282
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 21100 10146 21128 11494
rect 21192 10266 21220 14311
rect 21284 13938 21312 14350
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21284 13394 21312 13874
rect 21272 13388 21324 13394
rect 21272 13330 21324 13336
rect 21284 12850 21312 13330
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 21284 12238 21312 12786
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21284 11830 21312 12174
rect 21272 11824 21324 11830
rect 21272 11766 21324 11772
rect 21284 11082 21312 11766
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 21180 10260 21232 10266
rect 21180 10202 21232 10208
rect 21100 10118 21220 10146
rect 20916 8634 20944 8774
rect 21008 8758 21128 8786
rect 20904 8628 20956 8634
rect 20904 8570 20956 8576
rect 20996 8628 21048 8634
rect 20996 8570 21048 8576
rect 20904 8492 20956 8498
rect 20904 8434 20956 8440
rect 20812 7880 20864 7886
rect 20916 7857 20944 8434
rect 20812 7822 20864 7828
rect 20902 7848 20958 7857
rect 20902 7783 20958 7792
rect 20718 7440 20774 7449
rect 20718 7375 20720 7384
rect 20772 7375 20774 7384
rect 20720 7346 20772 7352
rect 20812 7336 20864 7342
rect 20812 7278 20864 7284
rect 20824 6798 20852 7278
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20916 6390 20944 7783
rect 20904 6384 20956 6390
rect 20718 6352 20774 6361
rect 20718 6287 20774 6296
rect 20902 6352 20904 6361
rect 20956 6352 20958 6361
rect 20902 6287 20958 6296
rect 20626 4584 20682 4593
rect 20626 4519 20682 4528
rect 20536 4480 20588 4486
rect 20536 4422 20588 4428
rect 20548 4146 20576 4422
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20732 3210 20760 6287
rect 20904 5704 20956 5710
rect 20902 5672 20904 5681
rect 20956 5672 20958 5681
rect 20824 5630 20902 5658
rect 20824 3738 20852 5630
rect 20902 5607 20958 5616
rect 20904 5568 20956 5574
rect 20904 5510 20956 5516
rect 20916 4690 20944 5510
rect 21008 5166 21036 8570
rect 21100 7478 21128 8758
rect 21192 8634 21220 10118
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 21088 7472 21140 7478
rect 21088 7414 21140 7420
rect 21192 7324 21220 8366
rect 21100 7296 21220 7324
rect 21100 6254 21128 7296
rect 21088 6248 21140 6254
rect 21088 6190 21140 6196
rect 21180 6248 21232 6254
rect 21180 6190 21232 6196
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 21100 5001 21128 6190
rect 21192 5234 21220 6190
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 21086 4992 21142 5001
rect 21086 4927 21142 4936
rect 21100 4758 21128 4927
rect 21284 4826 21312 11018
rect 21376 8090 21404 15943
rect 21468 8430 21496 17546
rect 21560 17542 21588 22222
rect 21836 22114 21864 22222
rect 21914 22200 21970 23000
rect 22466 22200 22522 23000
rect 21928 22114 21956 22200
rect 21836 22086 21956 22114
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 22480 18970 22508 22200
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 21548 17536 21600 17542
rect 21548 17478 21600 17484
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21548 14884 21600 14890
rect 21548 14826 21600 14832
rect 21560 12170 21588 14826
rect 22192 14816 22244 14822
rect 22192 14758 22244 14764
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21640 14068 21692 14074
rect 21640 14010 21692 14016
rect 21652 12918 21680 14010
rect 22006 13288 22062 13297
rect 22006 13223 22062 13232
rect 22020 13190 22048 13223
rect 22008 13184 22060 13190
rect 22008 13126 22060 13132
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21640 12912 21692 12918
rect 21640 12854 21692 12860
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21548 11620 21600 11626
rect 21548 11562 21600 11568
rect 21456 8424 21508 8430
rect 21456 8366 21508 8372
rect 21364 8084 21416 8090
rect 21364 8026 21416 8032
rect 21560 6254 21588 11562
rect 21548 6248 21600 6254
rect 21548 6190 21600 6196
rect 21652 5098 21680 12854
rect 22100 12164 22152 12170
rect 22100 12106 22152 12112
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 22006 11520 22062 11529
rect 22006 11455 22062 11464
rect 22020 11082 22048 11455
rect 22008 11076 22060 11082
rect 22008 11018 22060 11024
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 22006 10704 22062 10713
rect 22006 10639 22008 10648
rect 22060 10639 22062 10648
rect 22008 10610 22060 10616
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 21640 5092 21692 5098
rect 21640 5034 21692 5040
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 21088 4752 21140 4758
rect 21088 4694 21140 4700
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 21178 4584 21234 4593
rect 21178 4519 21234 4528
rect 21192 4146 21220 4519
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 21180 4140 21232 4146
rect 21180 4082 21232 4088
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 22112 3670 22140 12106
rect 22204 8022 22232 14758
rect 22560 13184 22612 13190
rect 22560 13126 22612 13132
rect 22376 11076 22428 11082
rect 22376 11018 22428 11024
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22296 8906 22324 10610
rect 22284 8900 22336 8906
rect 22284 8842 22336 8848
rect 22192 8016 22244 8022
rect 22192 7958 22244 7964
rect 22296 5710 22324 8842
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22100 3664 22152 3670
rect 22100 3606 22152 3612
rect 22388 3602 22416 11018
rect 22572 6662 22600 13126
rect 22560 6656 22612 6662
rect 22560 6598 22612 6604
rect 22376 3596 22428 3602
rect 22376 3538 22428 3544
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 20640 3182 20760 3210
rect 20902 3224 20958 3233
rect 21742 3227 22050 3236
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20640 2802 20668 3182
rect 20902 3159 20958 3168
rect 22468 3188 22520 3194
rect 20720 3120 20772 3126
rect 20720 3062 20772 3068
rect 20732 2938 20760 3062
rect 20916 2961 20944 3159
rect 22468 3130 22520 3136
rect 20902 2952 20958 2961
rect 20732 2910 20852 2938
rect 20640 2774 20760 2802
rect 20732 2650 20760 2774
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20350 1728 20406 1737
rect 20350 1663 20406 1672
rect 20824 800 20852 2910
rect 20902 2887 20958 2896
rect 21364 2916 21416 2922
rect 21364 2858 21416 2864
rect 21376 800 21404 2858
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 11532 734 11744 762
rect 11978 0 12034 800
rect 12530 0 12586 800
rect 13082 0 13138 800
rect 13634 0 13690 800
rect 14186 0 14242 800
rect 14738 0 14794 800
rect 15290 0 15346 800
rect 15842 0 15898 800
rect 16394 0 16450 800
rect 16946 0 17002 800
rect 17498 0 17554 800
rect 18050 0 18106 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19706 0 19762 800
rect 20258 0 20314 800
rect 20810 0 20866 800
rect 21362 0 21418 800
rect 21560 762 21588 2790
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 21836 870 21956 898
rect 21836 762 21864 870
rect 21928 800 21956 870
rect 22480 800 22508 3130
rect 21560 734 21864 762
rect 21914 0 21970 800
rect 22466 0 22522 800
<< via2 >>
rect 386 18672 442 18728
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 5630 20204 5632 20224
rect 5632 20204 5684 20224
rect 5684 20204 5686 20224
rect 5630 20168 5686 20204
rect 4618 18808 4674 18864
rect 4066 17176 4122 17232
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 1490 3032 1546 3088
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3514 5752 3570 5808
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 4618 9016 4674 9072
rect 4526 6840 4582 6896
rect 5446 13368 5502 13424
rect 5078 11192 5134 11248
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 5998 17312 6054 17368
rect 5722 13232 5778 13288
rect 5630 12280 5686 12336
rect 5354 6840 5410 6896
rect 4802 3984 4858 4040
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6090 15428 6146 15464
rect 6090 15408 6092 15428
rect 6092 15408 6144 15428
rect 6144 15408 6146 15428
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 6550 12688 6606 12744
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6182 11736 6238 11792
rect 6090 11056 6146 11112
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 5998 9968 6054 10024
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 7562 15952 7618 16008
rect 7286 14864 7342 14920
rect 6826 9968 6882 10024
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 5906 7248 5962 7304
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 7562 15428 7618 15464
rect 7562 15408 7564 15428
rect 7564 15408 7616 15428
rect 7616 15408 7618 15428
rect 7654 11872 7710 11928
rect 8206 17584 8262 17640
rect 7838 12824 7894 12880
rect 7838 11872 7894 11928
rect 8482 12416 8538 12472
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6550 3848 6606 3904
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 8206 11736 8262 11792
rect 8114 10104 8170 10160
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 9034 18672 9090 18728
rect 9310 19760 9366 19816
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8758 17040 8814 17096
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 8390 10784 8446 10840
rect 8390 6996 8446 7032
rect 8390 6976 8392 6996
rect 8392 6976 8444 6996
rect 8444 6976 8446 6996
rect 8574 10648 8630 10704
rect 8574 9968 8630 10024
rect 9218 12688 9274 12744
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 9034 10920 9090 10976
rect 8850 10512 8906 10568
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 9310 9580 9366 9616
rect 9310 9560 9312 9580
rect 9312 9560 9364 9580
rect 9364 9560 9366 9580
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 9218 6296 9274 6352
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 10506 19896 10562 19952
rect 9770 17992 9826 18048
rect 9678 10376 9734 10432
rect 9862 9424 9918 9480
rect 9678 8372 9680 8392
rect 9680 8372 9732 8392
rect 9732 8372 9734 8392
rect 9678 8336 9734 8372
rect 10138 14184 10194 14240
rect 10322 14048 10378 14104
rect 10138 10804 10194 10840
rect 10138 10784 10140 10804
rect 10140 10784 10192 10804
rect 10192 10784 10194 10804
rect 10138 8200 10194 8256
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 12162 20304 12218 20360
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11334 18128 11390 18184
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11150 14184 11206 14240
rect 10782 10920 10838 10976
rect 10782 10512 10838 10568
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11794 13776 11850 13832
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 10966 10920 11022 10976
rect 12714 19896 12770 19952
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 12162 15952 12218 16008
rect 12622 15408 12678 15464
rect 12254 13776 12310 13832
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 10690 8336 10746 8392
rect 10506 7384 10562 7440
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 9770 3848 9826 3904
rect 9126 3576 9182 3632
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 9862 3188 9918 3224
rect 10414 4664 10470 4720
rect 9862 3168 9864 3188
rect 9864 3168 9916 3188
rect 9916 3168 9918 3188
rect 9770 3032 9826 3088
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11978 11600 12034 11656
rect 11794 9288 11850 9344
rect 12162 11736 12218 11792
rect 12162 10956 12164 10976
rect 12164 10956 12216 10976
rect 12216 10956 12218 10976
rect 12162 10920 12218 10956
rect 12162 10804 12218 10840
rect 12162 10784 12164 10804
rect 12164 10784 12216 10804
rect 12216 10784 12218 10804
rect 12162 9560 12218 9616
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11150 6860 11206 6896
rect 11150 6840 11152 6860
rect 11152 6840 11204 6860
rect 11204 6840 11206 6860
rect 11886 8064 11942 8120
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 12898 15272 12954 15328
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 12622 11092 12624 11112
rect 12624 11092 12676 11112
rect 12676 11092 12678 11112
rect 12622 11056 12678 11092
rect 12530 10784 12586 10840
rect 11978 6976 12034 7032
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 10598 5072 10654 5128
rect 10598 4120 10654 4176
rect 10874 3984 10930 4040
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11058 3984 11114 4040
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11058 2896 11114 2952
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12162 6160 12218 6216
rect 12530 9288 12586 9344
rect 12346 8200 12402 8256
rect 12346 7928 12402 7984
rect 12898 11328 12954 11384
rect 12898 11076 12954 11112
rect 12898 11056 12900 11076
rect 12900 11056 12952 11076
rect 12952 11056 12954 11076
rect 12898 10376 12954 10432
rect 12806 10260 12862 10296
rect 12806 10240 12808 10260
rect 12808 10240 12860 10260
rect 12860 10240 12862 10260
rect 12806 9560 12862 9616
rect 12530 6704 12586 6760
rect 12346 5616 12402 5672
rect 12070 3068 12072 3088
rect 12072 3068 12124 3088
rect 12124 3068 12126 3088
rect 12070 3032 12126 3068
rect 12714 6432 12770 6488
rect 13082 10956 13084 10976
rect 13084 10956 13136 10976
rect 13136 10956 13138 10976
rect 13082 10920 13138 10956
rect 13266 7792 13322 7848
rect 12806 6160 12862 6216
rect 13174 6704 13230 6760
rect 14646 20204 14648 20224
rect 14648 20204 14700 20224
rect 14700 20204 14702 20224
rect 14646 20168 14702 20204
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13634 11328 13690 11384
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 14094 11092 14096 11112
rect 14096 11092 14148 11112
rect 14148 11092 14150 11112
rect 14094 11056 14150 11092
rect 13542 8628 13598 8664
rect 13542 8608 13544 8628
rect 13544 8608 13596 8628
rect 13596 8608 13598 8628
rect 13450 7928 13506 7984
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 14186 9016 14242 9072
rect 13818 8472 13874 8528
rect 15382 19760 15438 19816
rect 15290 18808 15346 18864
rect 15566 17720 15622 17776
rect 14462 9696 14518 9752
rect 13726 8084 13782 8120
rect 13726 8064 13728 8084
rect 13728 8064 13780 8084
rect 13780 8064 13782 8084
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13542 6976 13598 7032
rect 13450 6704 13506 6760
rect 13542 6160 13598 6216
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 13818 5752 13874 5808
rect 13910 5208 13966 5264
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 16762 20168 16818 20224
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 16302 19352 16358 19408
rect 15290 13368 15346 13424
rect 14922 10784 14978 10840
rect 14922 9580 14978 9616
rect 14922 9560 14924 9580
rect 14924 9560 14976 9580
rect 14976 9560 14978 9580
rect 15106 9460 15108 9480
rect 15108 9460 15160 9480
rect 15160 9460 15162 9480
rect 15106 9424 15162 9460
rect 15198 8628 15254 8664
rect 15198 8608 15200 8628
rect 15200 8608 15252 8628
rect 15252 8608 15254 8628
rect 14370 4936 14426 4992
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 14186 2896 14242 2952
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 14922 3712 14978 3768
rect 15658 15272 15714 15328
rect 16486 18692 16542 18728
rect 16486 18672 16488 18692
rect 16488 18672 16540 18692
rect 16540 18672 16542 18692
rect 16670 18692 16726 18728
rect 16670 18672 16672 18692
rect 16672 18672 16724 18692
rect 16724 18672 16726 18692
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 15290 6296 15346 6352
rect 15198 6024 15254 6080
rect 15566 8780 15568 8800
rect 15568 8780 15620 8800
rect 15620 8780 15622 8800
rect 15566 8744 15622 8780
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16854 13676 16856 13696
rect 16856 13676 16908 13696
rect 16908 13676 16910 13696
rect 16854 13640 16910 13676
rect 15934 8200 15990 8256
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 18694 20440 18750 20496
rect 18234 19896 18290 19952
rect 18786 20304 18842 20360
rect 18602 19896 18658 19952
rect 17958 19760 18014 19816
rect 17498 19352 17554 19408
rect 17130 16496 17186 16552
rect 17038 15952 17094 16008
rect 16946 12008 17002 12064
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 17038 11076 17094 11112
rect 17038 11056 17040 11076
rect 17040 11056 17092 11076
rect 17092 11056 17094 11076
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16946 10104 17002 10160
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16946 9560 17002 9616
rect 16210 8200 16266 8256
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 17314 10648 17370 10704
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 17682 15000 17738 15056
rect 17406 9016 17462 9072
rect 16118 6704 16174 6760
rect 15842 5364 15898 5400
rect 15842 5344 15844 5364
rect 15844 5344 15896 5364
rect 15896 5344 15898 5364
rect 15842 4120 15898 4176
rect 15750 3440 15806 3496
rect 15750 2896 15806 2952
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 17038 6432 17094 6488
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 17038 5752 17094 5808
rect 17866 13368 17922 13424
rect 18234 13404 18236 13424
rect 18236 13404 18288 13424
rect 18288 13404 18290 13424
rect 18234 13368 18290 13404
rect 17406 5888 17462 5944
rect 17498 5772 17554 5808
rect 17498 5752 17500 5772
rect 17500 5752 17552 5772
rect 17552 5752 17554 5772
rect 17774 6196 17776 6216
rect 17776 6196 17828 6216
rect 17828 6196 17830 6216
rect 17774 6160 17830 6196
rect 16854 3984 16910 4040
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 18142 10804 18198 10840
rect 18142 10784 18144 10804
rect 18144 10784 18196 10804
rect 18196 10784 18198 10804
rect 17958 10124 18014 10160
rect 17958 10104 17960 10124
rect 17960 10104 18012 10124
rect 18012 10104 18014 10124
rect 17958 9424 18014 9480
rect 18694 19216 18750 19272
rect 18602 16496 18658 16552
rect 18418 11192 18474 11248
rect 18050 7248 18106 7304
rect 18142 7112 18198 7168
rect 18326 7520 18382 7576
rect 17958 5752 18014 5808
rect 17958 5072 18014 5128
rect 17958 4564 17960 4584
rect 17960 4564 18012 4584
rect 18012 4564 18014 4584
rect 17958 4528 18014 4564
rect 17958 3712 18014 3768
rect 17866 3052 17922 3088
rect 17866 3032 17868 3052
rect 17868 3032 17920 3052
rect 17920 3032 17922 3052
rect 18142 4936 18198 4992
rect 18142 3984 18198 4040
rect 18786 13912 18842 13968
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19614 20848 19670 20904
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 20534 21256 20590 21312
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19614 16768 19670 16824
rect 18878 13776 18934 13832
rect 18694 11736 18750 11792
rect 18786 10648 18842 10704
rect 18786 10512 18842 10568
rect 18694 9832 18750 9888
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 18970 10412 18972 10432
rect 18972 10412 19024 10432
rect 19024 10412 19026 10432
rect 18970 10376 19026 10412
rect 18878 9560 18934 9616
rect 18694 8336 18750 8392
rect 18694 7792 18750 7848
rect 18418 6024 18474 6080
rect 18418 5072 18474 5128
rect 18326 3304 18382 3360
rect 18234 3032 18290 3088
rect 18970 7928 19026 7984
rect 18878 6704 18934 6760
rect 18694 5072 18750 5128
rect 18602 4256 18658 4312
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19982 15544 20038 15600
rect 19890 15308 19892 15328
rect 19892 15308 19944 15328
rect 19944 15308 19946 15328
rect 19890 15272 19946 15308
rect 19890 13232 19946 13288
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19614 7284 19616 7304
rect 19616 7284 19668 7304
rect 19668 7284 19670 7304
rect 19614 7248 19670 7284
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19246 6840 19302 6896
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 18786 3440 18842 3496
rect 18970 3576 19026 3632
rect 18878 1944 18934 2000
rect 21086 18808 21142 18864
rect 19890 8472 19946 8528
rect 20442 18264 20498 18320
rect 20534 17040 20590 17096
rect 20902 17584 20958 17640
rect 20718 16224 20774 16280
rect 20626 14728 20682 14784
rect 20626 11056 20682 11112
rect 20258 10004 20260 10024
rect 20260 10004 20312 10024
rect 20312 10004 20314 10024
rect 20258 9968 20314 10004
rect 20258 8628 20314 8664
rect 20258 8608 20260 8628
rect 20260 8608 20312 8628
rect 20312 8608 20314 8628
rect 19706 5208 19762 5264
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 19890 4120 19946 4176
rect 19338 2896 19394 2952
rect 19982 4020 19984 4040
rect 19984 4020 20036 4040
rect 20036 4020 20038 4040
rect 19982 3984 20038 4020
rect 20166 5480 20222 5536
rect 20258 4684 20314 4720
rect 20258 4664 20260 4684
rect 20260 4664 20312 4684
rect 20312 4664 20314 4684
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 19154 2488 19210 2544
rect 21362 15952 21418 16008
rect 21178 14320 21234 14376
rect 20902 7792 20958 7848
rect 20718 7404 20774 7440
rect 20718 7384 20720 7404
rect 20720 7384 20772 7404
rect 20772 7384 20774 7404
rect 20718 6296 20774 6352
rect 20902 6332 20904 6352
rect 20904 6332 20956 6352
rect 20956 6332 20958 6352
rect 20902 6296 20958 6332
rect 20626 4528 20682 4584
rect 20902 5652 20904 5672
rect 20904 5652 20956 5672
rect 20956 5652 20958 5672
rect 20902 5616 20958 5652
rect 21086 4936 21142 4992
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 22006 13232 22062 13288
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 22006 11464 22062 11520
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 22006 10668 22062 10704
rect 22006 10648 22008 10668
rect 22008 10648 22060 10668
rect 22060 10648 22062 10668
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 21178 4528 21234 4584
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 20902 3168 20958 3224
rect 20350 1672 20406 1728
rect 20902 2896 20958 2952
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
<< metal3 >>
rect 20529 21314 20595 21317
rect 22200 21314 23000 21344
rect 20529 21312 23000 21314
rect 20529 21256 20534 21312
rect 20590 21256 23000 21312
rect 20529 21254 23000 21256
rect 20529 21251 20595 21254
rect 22200 21224 23000 21254
rect 19609 20906 19675 20909
rect 22200 20906 23000 20936
rect 19609 20904 23000 20906
rect 19609 20848 19614 20904
rect 19670 20848 23000 20904
rect 19609 20846 23000 20848
rect 19609 20843 19675 20846
rect 22200 20816 23000 20846
rect 6144 20704 6460 20705
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 18689 20498 18755 20501
rect 22200 20498 23000 20528
rect 18689 20496 23000 20498
rect 18689 20440 18694 20496
rect 18750 20440 23000 20496
rect 18689 20438 23000 20440
rect 18689 20435 18755 20438
rect 22200 20408 23000 20438
rect 12157 20362 12223 20365
rect 18781 20362 18847 20365
rect 12157 20360 18847 20362
rect 12157 20304 12162 20360
rect 12218 20304 18786 20360
rect 18842 20304 18847 20360
rect 12157 20302 18847 20304
rect 12157 20299 12223 20302
rect 18781 20299 18847 20302
rect 5625 20226 5691 20229
rect 5942 20226 5948 20228
rect 5625 20224 5948 20226
rect 5625 20168 5630 20224
rect 5686 20168 5948 20224
rect 5625 20166 5948 20168
rect 5625 20163 5691 20166
rect 5942 20164 5948 20166
rect 6012 20164 6018 20228
rect 14406 20164 14412 20228
rect 14476 20226 14482 20228
rect 14641 20226 14707 20229
rect 14476 20224 14707 20226
rect 14476 20168 14646 20224
rect 14702 20168 14707 20224
rect 14476 20166 14707 20168
rect 14476 20164 14482 20166
rect 14641 20163 14707 20166
rect 16757 20226 16823 20229
rect 17350 20226 17356 20228
rect 16757 20224 17356 20226
rect 16757 20168 16762 20224
rect 16818 20168 17356 20224
rect 16757 20166 17356 20168
rect 16757 20163 16823 20166
rect 17350 20164 17356 20166
rect 17420 20164 17426 20228
rect 3545 20160 3861 20161
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 19139 20095 19455 20096
rect 22200 20090 23000 20120
rect 19566 20030 23000 20090
rect 10501 19954 10567 19957
rect 12198 19954 12204 19956
rect 10501 19952 12204 19954
rect 10501 19896 10506 19952
rect 10562 19896 12204 19952
rect 10501 19894 12204 19896
rect 10501 19891 10567 19894
rect 12198 19892 12204 19894
rect 12268 19892 12274 19956
rect 12709 19954 12775 19957
rect 18229 19954 18295 19957
rect 12709 19952 18295 19954
rect 12709 19896 12714 19952
rect 12770 19896 18234 19952
rect 18290 19896 18295 19952
rect 12709 19894 18295 19896
rect 12709 19891 12775 19894
rect 18229 19891 18295 19894
rect 18597 19954 18663 19957
rect 19566 19954 19626 20030
rect 22200 20000 23000 20030
rect 18597 19952 19626 19954
rect 18597 19896 18602 19952
rect 18658 19896 19626 19952
rect 18597 19894 19626 19896
rect 18597 19891 18663 19894
rect 9305 19818 9371 19821
rect 15377 19818 15443 19821
rect 9305 19816 15443 19818
rect 9305 19760 9310 19816
rect 9366 19760 15382 19816
rect 15438 19760 15443 19816
rect 9305 19758 15443 19760
rect 9305 19755 9371 19758
rect 15377 19755 15443 19758
rect 17953 19818 18019 19821
rect 17953 19816 22202 19818
rect 17953 19760 17958 19816
rect 18014 19760 22202 19816
rect 17953 19758 22202 19760
rect 17953 19755 18019 19758
rect 22142 19712 22202 19758
rect 22142 19622 23000 19712
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 22200 19592 23000 19622
rect 21738 19551 22054 19552
rect 16297 19410 16363 19413
rect 17493 19410 17559 19413
rect 16297 19408 17559 19410
rect 16297 19352 16302 19408
rect 16358 19352 17498 19408
rect 17554 19352 17559 19408
rect 16297 19350 17559 19352
rect 16297 19347 16363 19350
rect 17493 19347 17559 19350
rect 18689 19274 18755 19277
rect 22200 19274 23000 19304
rect 18689 19272 23000 19274
rect 18689 19216 18694 19272
rect 18750 19216 23000 19272
rect 18689 19214 23000 19216
rect 18689 19211 18755 19214
rect 22200 19184 23000 19214
rect 3545 19072 3861 19073
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 4613 18866 4679 18869
rect 15285 18866 15351 18869
rect 4613 18864 15351 18866
rect 4613 18808 4618 18864
rect 4674 18808 15290 18864
rect 15346 18808 15351 18864
rect 4613 18806 15351 18808
rect 4613 18803 4679 18806
rect 15285 18803 15351 18806
rect 21081 18866 21147 18869
rect 22200 18866 23000 18896
rect 21081 18864 23000 18866
rect 21081 18808 21086 18864
rect 21142 18808 23000 18864
rect 21081 18806 23000 18808
rect 21081 18803 21147 18806
rect 22200 18776 23000 18806
rect 381 18730 447 18733
rect 9029 18730 9095 18733
rect 381 18728 9095 18730
rect 381 18672 386 18728
rect 442 18672 9034 18728
rect 9090 18672 9095 18728
rect 381 18670 9095 18672
rect 381 18667 447 18670
rect 9029 18667 9095 18670
rect 16481 18730 16547 18733
rect 16665 18730 16731 18733
rect 16481 18728 16731 18730
rect 16481 18672 16486 18728
rect 16542 18672 16670 18728
rect 16726 18672 16731 18728
rect 16481 18670 16731 18672
rect 16481 18667 16547 18670
rect 16665 18667 16731 18670
rect 6144 18528 6460 18529
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 21738 18463 22054 18464
rect 22200 18458 23000 18488
rect 22142 18368 23000 18458
rect 20437 18322 20503 18325
rect 22142 18322 22202 18368
rect 20437 18320 22202 18322
rect 20437 18264 20442 18320
rect 20498 18264 22202 18320
rect 20437 18262 22202 18264
rect 20437 18259 20503 18262
rect 9438 18124 9444 18188
rect 9508 18186 9514 18188
rect 11329 18186 11395 18189
rect 9508 18184 11395 18186
rect 9508 18128 11334 18184
rect 11390 18128 11395 18184
rect 9508 18126 11395 18128
rect 9508 18124 9514 18126
rect 11329 18123 11395 18126
rect 9765 18052 9831 18053
rect 9765 18048 9812 18052
rect 9876 18050 9882 18052
rect 9765 17992 9770 18048
rect 9765 17988 9812 17992
rect 9876 17990 9922 18050
rect 9876 17988 9882 17990
rect 20294 17988 20300 18052
rect 20364 18050 20370 18052
rect 22200 18050 23000 18080
rect 20364 17990 23000 18050
rect 20364 17988 20370 17990
rect 9765 17987 9831 17988
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 22200 17960 23000 17990
rect 19139 17919 19455 17920
rect 10358 17716 10364 17780
rect 10428 17778 10434 17780
rect 15561 17778 15627 17781
rect 10428 17776 15627 17778
rect 10428 17720 15566 17776
rect 15622 17720 15627 17776
rect 10428 17718 15627 17720
rect 10428 17716 10434 17718
rect 15561 17715 15627 17718
rect 8201 17642 8267 17645
rect 13670 17642 13676 17644
rect 8201 17640 13676 17642
rect 8201 17584 8206 17640
rect 8262 17584 13676 17640
rect 8201 17582 13676 17584
rect 8201 17579 8267 17582
rect 13670 17580 13676 17582
rect 13740 17580 13746 17644
rect 20897 17642 20963 17645
rect 22200 17642 23000 17672
rect 20897 17640 23000 17642
rect 20897 17584 20902 17640
rect 20958 17584 23000 17640
rect 20897 17582 23000 17584
rect 20897 17579 20963 17582
rect 22200 17552 23000 17582
rect 6144 17440 6460 17441
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 5993 17370 6059 17373
rect 5950 17368 6059 17370
rect 5950 17312 5998 17368
rect 6054 17312 6059 17368
rect 5950 17307 6059 17312
rect 0 17234 800 17264
rect 4061 17234 4127 17237
rect 0 17232 4127 17234
rect 0 17176 4066 17232
rect 4122 17176 4127 17232
rect 0 17174 4127 17176
rect 5950 17234 6010 17307
rect 15878 17234 15884 17236
rect 5950 17174 15884 17234
rect 0 17144 800 17174
rect 4061 17171 4127 17174
rect 15878 17172 15884 17174
rect 15948 17172 15954 17236
rect 22200 17234 23000 17264
rect 20670 17174 23000 17234
rect 8753 17098 8819 17101
rect 15510 17098 15516 17100
rect 8753 17096 15516 17098
rect 8753 17040 8758 17096
rect 8814 17040 15516 17096
rect 8753 17038 15516 17040
rect 8753 17035 8819 17038
rect 15510 17036 15516 17038
rect 15580 17036 15586 17100
rect 20529 17098 20595 17101
rect 20670 17098 20730 17174
rect 22200 17144 23000 17174
rect 20529 17096 20730 17098
rect 20529 17040 20534 17096
rect 20590 17040 20730 17096
rect 20529 17038 20730 17040
rect 20529 17035 20595 17038
rect 3545 16896 3861 16897
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 19139 16831 19455 16832
rect 19609 16826 19675 16829
rect 22200 16826 23000 16856
rect 19609 16824 23000 16826
rect 19609 16768 19614 16824
rect 19670 16768 23000 16824
rect 19609 16766 23000 16768
rect 19609 16763 19675 16766
rect 22200 16736 23000 16766
rect 12934 16492 12940 16556
rect 13004 16554 13010 16556
rect 17125 16554 17191 16557
rect 13004 16552 17191 16554
rect 13004 16496 17130 16552
rect 17186 16496 17191 16552
rect 13004 16494 17191 16496
rect 13004 16492 13010 16494
rect 17125 16491 17191 16494
rect 18597 16554 18663 16557
rect 18597 16552 22202 16554
rect 18597 16496 18602 16552
rect 18658 16496 22202 16552
rect 18597 16494 22202 16496
rect 18597 16491 18663 16494
rect 22142 16448 22202 16494
rect 22142 16358 23000 16448
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 22200 16328 23000 16358
rect 21738 16287 22054 16288
rect 20713 16282 20779 16285
rect 18600 16280 20779 16282
rect 18600 16224 20718 16280
rect 20774 16224 20779 16280
rect 18600 16222 20779 16224
rect 13118 16084 13124 16148
rect 13188 16146 13194 16148
rect 18600 16146 18660 16222
rect 20713 16219 20779 16222
rect 13188 16086 18660 16146
rect 13188 16084 13194 16086
rect 7557 16010 7623 16013
rect 12157 16010 12223 16013
rect 7557 16008 12223 16010
rect 7557 15952 7562 16008
rect 7618 15952 12162 16008
rect 12218 15952 12223 16008
rect 7557 15950 12223 15952
rect 7557 15947 7623 15950
rect 12157 15947 12223 15950
rect 14774 15948 14780 16012
rect 14844 16010 14850 16012
rect 17033 16010 17099 16013
rect 14844 16008 17099 16010
rect 14844 15952 17038 16008
rect 17094 15952 17099 16008
rect 14844 15950 17099 15952
rect 14844 15948 14850 15950
rect 17033 15947 17099 15950
rect 21357 16010 21423 16013
rect 22200 16010 23000 16040
rect 21357 16008 23000 16010
rect 21357 15952 21362 16008
rect 21418 15952 23000 16008
rect 21357 15950 23000 15952
rect 21357 15947 21423 15950
rect 22200 15920 23000 15950
rect 3545 15808 3861 15809
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 19977 15602 20043 15605
rect 22200 15602 23000 15632
rect 19977 15600 23000 15602
rect 19977 15544 19982 15600
rect 20038 15544 23000 15600
rect 19977 15542 23000 15544
rect 19977 15539 20043 15542
rect 22200 15512 23000 15542
rect 6085 15466 6151 15469
rect 6678 15466 6684 15468
rect 6085 15464 6684 15466
rect 6085 15408 6090 15464
rect 6146 15408 6684 15464
rect 6085 15406 6684 15408
rect 6085 15403 6151 15406
rect 6678 15404 6684 15406
rect 6748 15466 6754 15468
rect 7557 15466 7623 15469
rect 6748 15464 7623 15466
rect 6748 15408 7562 15464
rect 7618 15408 7623 15464
rect 6748 15406 7623 15408
rect 6748 15404 6754 15406
rect 7557 15403 7623 15406
rect 12617 15466 12683 15469
rect 17166 15466 17172 15468
rect 12617 15464 17172 15466
rect 12617 15408 12622 15464
rect 12678 15408 17172 15464
rect 12617 15406 17172 15408
rect 12617 15403 12683 15406
rect 17166 15404 17172 15406
rect 17236 15404 17242 15468
rect 11830 15268 11836 15332
rect 11900 15330 11906 15332
rect 12893 15330 12959 15333
rect 11900 15328 12959 15330
rect 11900 15272 12898 15328
rect 12954 15272 12959 15328
rect 11900 15270 12959 15272
rect 11900 15268 11906 15270
rect 12893 15267 12959 15270
rect 15142 15268 15148 15332
rect 15212 15330 15218 15332
rect 15653 15330 15719 15333
rect 15212 15328 15719 15330
rect 15212 15272 15658 15328
rect 15714 15272 15719 15328
rect 15212 15270 15719 15272
rect 15212 15268 15218 15270
rect 15653 15267 15719 15270
rect 19742 15268 19748 15332
rect 19812 15330 19818 15332
rect 19885 15330 19951 15333
rect 19812 15328 19951 15330
rect 19812 15272 19890 15328
rect 19946 15272 19951 15328
rect 19812 15270 19951 15272
rect 19812 15268 19818 15270
rect 19885 15267 19951 15270
rect 6144 15264 6460 15265
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 21738 15199 22054 15200
rect 22200 15194 23000 15224
rect 22142 15104 23000 15194
rect 17677 15058 17743 15061
rect 22142 15058 22202 15104
rect 17677 15056 22202 15058
rect 17677 15000 17682 15056
rect 17738 15000 22202 15056
rect 17677 14998 22202 15000
rect 17677 14995 17743 14998
rect 7281 14922 7347 14925
rect 19006 14922 19012 14924
rect 7281 14920 19012 14922
rect 7281 14864 7286 14920
rect 7342 14864 19012 14920
rect 7281 14862 19012 14864
rect 7281 14859 7347 14862
rect 19006 14860 19012 14862
rect 19076 14860 19082 14924
rect 20621 14786 20687 14789
rect 22200 14786 23000 14816
rect 20621 14784 23000 14786
rect 20621 14728 20626 14784
rect 20682 14728 23000 14784
rect 20621 14726 23000 14728
rect 20621 14723 20687 14726
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 22200 14696 23000 14726
rect 19139 14655 19455 14656
rect 21173 14378 21239 14381
rect 22200 14378 23000 14408
rect 21173 14376 23000 14378
rect 21173 14320 21178 14376
rect 21234 14320 23000 14376
rect 21173 14318 23000 14320
rect 21173 14315 21239 14318
rect 22200 14288 23000 14318
rect 10133 14242 10199 14245
rect 11145 14242 11211 14245
rect 10133 14240 11211 14242
rect 10133 14184 10138 14240
rect 10194 14184 11150 14240
rect 11206 14184 11211 14240
rect 10133 14182 11211 14184
rect 10133 14179 10199 14182
rect 11145 14179 11211 14182
rect 6144 14176 6460 14177
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 8150 14044 8156 14108
rect 8220 14106 8226 14108
rect 10317 14106 10383 14109
rect 8220 14104 10383 14106
rect 8220 14048 10322 14104
rect 10378 14048 10383 14104
rect 8220 14046 10383 14048
rect 8220 14044 8226 14046
rect 10317 14043 10383 14046
rect 18781 13970 18847 13973
rect 22200 13970 23000 14000
rect 18781 13968 23000 13970
rect 18781 13912 18786 13968
rect 18842 13912 23000 13968
rect 18781 13910 23000 13912
rect 18781 13907 18847 13910
rect 22200 13880 23000 13910
rect 11789 13834 11855 13837
rect 12249 13834 12315 13837
rect 18873 13836 18939 13837
rect 15326 13834 15332 13836
rect 11789 13832 15332 13834
rect 11789 13776 11794 13832
rect 11850 13776 12254 13832
rect 12310 13776 15332 13832
rect 11789 13774 15332 13776
rect 11789 13771 11855 13774
rect 12249 13771 12315 13774
rect 15326 13772 15332 13774
rect 15396 13772 15402 13836
rect 18822 13772 18828 13836
rect 18892 13834 18939 13836
rect 18892 13832 18984 13834
rect 18934 13776 18984 13832
rect 18892 13774 18984 13776
rect 18892 13772 18939 13774
rect 18873 13771 18939 13772
rect 16849 13698 16915 13701
rect 17534 13698 17540 13700
rect 16849 13696 17540 13698
rect 16849 13640 16854 13696
rect 16910 13640 17540 13696
rect 16849 13638 17540 13640
rect 16849 13635 16915 13638
rect 17534 13636 17540 13638
rect 17604 13636 17610 13700
rect 3545 13632 3861 13633
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 19139 13567 19455 13568
rect 22200 13562 23000 13592
rect 20302 13502 23000 13562
rect 5441 13426 5507 13429
rect 11094 13426 11100 13428
rect 5441 13424 11100 13426
rect 5441 13368 5446 13424
rect 5502 13368 11100 13424
rect 5441 13366 11100 13368
rect 5441 13363 5507 13366
rect 11094 13364 11100 13366
rect 11164 13364 11170 13428
rect 15285 13426 15351 13429
rect 17861 13426 17927 13429
rect 15285 13424 17927 13426
rect 15285 13368 15290 13424
rect 15346 13368 17866 13424
rect 17922 13368 17927 13424
rect 15285 13366 17927 13368
rect 15285 13363 15351 13366
rect 17861 13363 17927 13366
rect 18229 13426 18295 13429
rect 20302 13426 20362 13502
rect 22200 13472 23000 13502
rect 18229 13424 20362 13426
rect 18229 13368 18234 13424
rect 18290 13368 20362 13424
rect 18229 13366 20362 13368
rect 18229 13363 18295 13366
rect 5717 13290 5783 13293
rect 5717 13288 6010 13290
rect 5717 13232 5722 13288
rect 5778 13232 6010 13288
rect 5717 13230 6010 13232
rect 5717 13227 5783 13230
rect 5950 12746 6010 13230
rect 17534 13228 17540 13292
rect 17604 13290 17610 13292
rect 19885 13290 19951 13293
rect 17604 13288 19951 13290
rect 17604 13232 19890 13288
rect 19946 13232 19951 13288
rect 17604 13230 19951 13232
rect 17604 13228 17610 13230
rect 19885 13227 19951 13230
rect 22001 13290 22067 13293
rect 22001 13288 22202 13290
rect 22001 13232 22006 13288
rect 22062 13232 22202 13288
rect 22001 13230 22202 13232
rect 22001 13227 22067 13230
rect 22142 13184 22202 13230
rect 22142 13094 23000 13184
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 22200 13064 23000 13094
rect 21738 13023 22054 13024
rect 7833 12882 7899 12885
rect 7966 12882 7972 12884
rect 7833 12880 7972 12882
rect 7833 12824 7838 12880
rect 7894 12824 7972 12880
rect 7833 12822 7972 12824
rect 7833 12819 7899 12822
rect 7966 12820 7972 12822
rect 8036 12820 8042 12884
rect 6545 12746 6611 12749
rect 9213 12746 9279 12749
rect 5950 12744 6611 12746
rect 5950 12688 6550 12744
rect 6606 12688 6611 12744
rect 5950 12686 6611 12688
rect 6545 12683 6611 12686
rect 8526 12744 9279 12746
rect 8526 12688 9218 12744
rect 9274 12688 9279 12744
rect 8526 12686 9279 12688
rect 3545 12544 3861 12545
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8526 12477 8586 12686
rect 9213 12683 9279 12686
rect 19926 12684 19932 12748
rect 19996 12746 20002 12748
rect 22200 12746 23000 12776
rect 19996 12686 23000 12746
rect 19996 12684 20002 12686
rect 22200 12656 23000 12686
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 8477 12472 8586 12477
rect 8477 12416 8482 12472
rect 8538 12416 8586 12472
rect 8477 12414 8586 12416
rect 8477 12411 8543 12414
rect 5625 12338 5691 12341
rect 22200 12338 23000 12368
rect 5625 12336 5826 12338
rect 5625 12280 5630 12336
rect 5686 12280 5826 12336
rect 5625 12278 5826 12280
rect 5625 12275 5691 12278
rect 5766 11794 5826 12278
rect 18094 12278 23000 12338
rect 16941 12066 17007 12069
rect 18094 12066 18154 12278
rect 22200 12248 23000 12278
rect 16941 12064 18154 12066
rect 16941 12008 16946 12064
rect 17002 12008 18154 12064
rect 16941 12006 18154 12008
rect 16941 12003 17007 12006
rect 6144 12000 6460 12001
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 21738 11935 22054 11936
rect 7649 11930 7715 11933
rect 7833 11930 7899 11933
rect 22200 11930 23000 11960
rect 7649 11928 7899 11930
rect 7649 11872 7654 11928
rect 7710 11872 7838 11928
rect 7894 11872 7899 11928
rect 7649 11870 7899 11872
rect 7649 11867 7715 11870
rect 7833 11867 7899 11870
rect 22142 11840 23000 11930
rect 6177 11794 6243 11797
rect 8201 11796 8267 11797
rect 8150 11794 8156 11796
rect 5766 11792 6243 11794
rect 5766 11736 6182 11792
rect 6238 11736 6243 11792
rect 5766 11734 6243 11736
rect 8110 11734 8156 11794
rect 8220 11792 8267 11796
rect 12157 11794 12223 11797
rect 8262 11736 8267 11792
rect 6177 11731 6243 11734
rect 8150 11732 8156 11734
rect 8220 11732 8267 11736
rect 8201 11731 8267 11732
rect 12022 11792 12223 11794
rect 12022 11736 12162 11792
rect 12218 11736 12223 11792
rect 12022 11734 12223 11736
rect 12022 11661 12082 11734
rect 12157 11731 12223 11734
rect 18689 11794 18755 11797
rect 22142 11794 22202 11840
rect 18689 11792 22202 11794
rect 18689 11736 18694 11792
rect 18750 11736 22202 11792
rect 18689 11734 22202 11736
rect 18689 11731 18755 11734
rect 11973 11656 12082 11661
rect 11973 11600 11978 11656
rect 12034 11600 12082 11656
rect 11973 11598 12082 11600
rect 11973 11595 12039 11598
rect 22001 11522 22067 11525
rect 22200 11522 23000 11552
rect 22001 11520 23000 11522
rect 22001 11464 22006 11520
rect 22062 11464 23000 11520
rect 22001 11462 23000 11464
rect 22001 11459 22067 11462
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 22200 11432 23000 11462
rect 19139 11391 19455 11392
rect 12893 11386 12959 11389
rect 13629 11386 13695 11389
rect 12893 11384 13695 11386
rect 12893 11328 12898 11384
rect 12954 11328 13634 11384
rect 13690 11328 13695 11384
rect 12893 11326 13695 11328
rect 12893 11323 12959 11326
rect 13629 11323 13695 11326
rect 5073 11250 5139 11253
rect 18413 11250 18479 11253
rect 5073 11248 18479 11250
rect 5073 11192 5078 11248
rect 5134 11192 18418 11248
rect 18474 11192 18479 11248
rect 5073 11190 18479 11192
rect 5073 11187 5139 11190
rect 18413 11187 18479 11190
rect 6085 11114 6151 11117
rect 8150 11114 8156 11116
rect 6085 11112 8156 11114
rect 6085 11056 6090 11112
rect 6146 11056 8156 11112
rect 6085 11054 8156 11056
rect 6085 11051 6151 11054
rect 8150 11052 8156 11054
rect 8220 11052 8226 11116
rect 12617 11114 12683 11117
rect 12893 11114 12959 11117
rect 14089 11114 14155 11117
rect 12617 11112 14155 11114
rect 12617 11056 12622 11112
rect 12678 11056 12898 11112
rect 12954 11056 14094 11112
rect 14150 11056 14155 11112
rect 12617 11054 14155 11056
rect 12617 11051 12683 11054
rect 12893 11051 12959 11054
rect 14089 11051 14155 11054
rect 17033 11114 17099 11117
rect 19558 11114 19564 11116
rect 17033 11112 19564 11114
rect 17033 11056 17038 11112
rect 17094 11056 19564 11112
rect 17033 11054 19564 11056
rect 17033 11051 17099 11054
rect 19558 11052 19564 11054
rect 19628 11114 19634 11116
rect 20621 11114 20687 11117
rect 22200 11114 23000 11144
rect 19628 11112 23000 11114
rect 19628 11056 20626 11112
rect 20682 11056 23000 11112
rect 19628 11054 23000 11056
rect 19628 11052 19634 11054
rect 20621 11051 20687 11054
rect 22200 11024 23000 11054
rect 9029 10978 9095 10981
rect 10777 10978 10843 10981
rect 10961 10978 11027 10981
rect 9029 10976 11027 10978
rect 9029 10920 9034 10976
rect 9090 10920 10782 10976
rect 10838 10920 10966 10976
rect 11022 10920 11027 10976
rect 9029 10918 11027 10920
rect 9029 10915 9095 10918
rect 10777 10915 10843 10918
rect 10961 10915 11027 10918
rect 12157 10978 12223 10981
rect 13077 10978 13143 10981
rect 12157 10976 13143 10978
rect 12157 10920 12162 10976
rect 12218 10920 13082 10976
rect 13138 10920 13143 10976
rect 12157 10918 13143 10920
rect 12157 10915 12223 10918
rect 13077 10915 13143 10918
rect 6144 10912 6460 10913
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 8385 10842 8451 10845
rect 10133 10842 10199 10845
rect 10358 10842 10364 10844
rect 8385 10840 8586 10842
rect 8385 10784 8390 10840
rect 8446 10784 8586 10840
rect 8385 10782 8586 10784
rect 8385 10779 8451 10782
rect 8526 10709 8586 10782
rect 10133 10840 10364 10842
rect 10133 10784 10138 10840
rect 10194 10784 10364 10840
rect 10133 10782 10364 10784
rect 10133 10779 10199 10782
rect 10358 10780 10364 10782
rect 10428 10780 10434 10844
rect 11830 10780 11836 10844
rect 11900 10842 11906 10844
rect 12157 10842 12223 10845
rect 11900 10840 12223 10842
rect 11900 10784 12162 10840
rect 12218 10784 12223 10840
rect 11900 10782 12223 10784
rect 11900 10780 11906 10782
rect 12157 10779 12223 10782
rect 12525 10842 12591 10845
rect 14917 10842 14983 10845
rect 18137 10842 18203 10845
rect 12525 10840 14983 10842
rect 12525 10784 12530 10840
rect 12586 10784 14922 10840
rect 14978 10784 14983 10840
rect 12525 10782 14983 10784
rect 12525 10779 12591 10782
rect 14917 10779 14983 10782
rect 17174 10840 18203 10842
rect 17174 10784 18142 10840
rect 18198 10784 18203 10840
rect 17174 10782 18203 10784
rect 8526 10704 8635 10709
rect 17174 10706 17234 10782
rect 18137 10779 18203 10782
rect 8526 10648 8574 10704
rect 8630 10648 8635 10704
rect 8526 10646 8635 10648
rect 8569 10643 8635 10646
rect 8710 10646 17234 10706
rect 17309 10706 17375 10709
rect 18781 10706 18847 10709
rect 17309 10704 18847 10706
rect 17309 10648 17314 10704
rect 17370 10648 18786 10704
rect 18842 10648 18847 10704
rect 17309 10646 18847 10648
rect 6678 10508 6684 10572
rect 6748 10570 6754 10572
rect 8710 10570 8770 10646
rect 17309 10643 17375 10646
rect 18781 10643 18847 10646
rect 22001 10706 22067 10709
rect 22200 10706 23000 10736
rect 22001 10704 23000 10706
rect 22001 10648 22006 10704
rect 22062 10648 23000 10704
rect 22001 10646 23000 10648
rect 22001 10643 22067 10646
rect 22200 10616 23000 10646
rect 6748 10510 8770 10570
rect 8845 10570 8911 10573
rect 9438 10570 9444 10572
rect 8845 10568 9444 10570
rect 8845 10512 8850 10568
rect 8906 10512 9444 10568
rect 8845 10510 9444 10512
rect 6748 10508 6754 10510
rect 8845 10507 8911 10510
rect 9438 10508 9444 10510
rect 9508 10508 9514 10572
rect 10777 10570 10843 10573
rect 18781 10570 18847 10573
rect 19926 10570 19932 10572
rect 10777 10568 18706 10570
rect 10777 10512 10782 10568
rect 10838 10512 18706 10568
rect 10777 10510 18706 10512
rect 10777 10507 10843 10510
rect 9673 10434 9739 10437
rect 12893 10434 12959 10437
rect 9673 10432 12959 10434
rect 9673 10376 9678 10432
rect 9734 10376 12898 10432
rect 12954 10376 12959 10432
rect 9673 10374 12959 10376
rect 18646 10434 18706 10510
rect 18781 10568 19932 10570
rect 18781 10512 18786 10568
rect 18842 10512 19932 10568
rect 18781 10510 19932 10512
rect 18781 10507 18847 10510
rect 19926 10508 19932 10510
rect 19996 10508 20002 10572
rect 18965 10434 19031 10437
rect 18646 10432 19031 10434
rect 18646 10376 18970 10432
rect 19026 10376 19031 10432
rect 18646 10374 19031 10376
rect 9673 10371 9739 10374
rect 12893 10371 12959 10374
rect 18965 10371 19031 10374
rect 3545 10368 3861 10369
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 19139 10303 19455 10304
rect 12801 10298 12867 10301
rect 13118 10298 13124 10300
rect 12801 10296 13124 10298
rect 12801 10240 12806 10296
rect 12862 10240 13124 10296
rect 12801 10238 13124 10240
rect 12801 10235 12867 10238
rect 13118 10236 13124 10238
rect 13188 10236 13194 10300
rect 22200 10298 23000 10328
rect 19566 10238 23000 10298
rect 8109 10162 8175 10165
rect 16941 10162 17007 10165
rect 8109 10160 17007 10162
rect 8109 10104 8114 10160
rect 8170 10104 16946 10160
rect 17002 10104 17007 10160
rect 8109 10102 17007 10104
rect 8109 10099 8175 10102
rect 16941 10099 17007 10102
rect 17953 10162 18019 10165
rect 19566 10162 19626 10238
rect 22200 10208 23000 10238
rect 17953 10160 19626 10162
rect 17953 10104 17958 10160
rect 18014 10104 19626 10160
rect 17953 10102 19626 10104
rect 17953 10099 18019 10102
rect 5993 10026 6059 10029
rect 6821 10026 6887 10029
rect 5993 10024 6887 10026
rect 5993 9968 5998 10024
rect 6054 9968 6826 10024
rect 6882 9968 6887 10024
rect 5993 9966 6887 9968
rect 5993 9963 6059 9966
rect 6821 9963 6887 9966
rect 8569 10026 8635 10029
rect 13670 10026 13676 10028
rect 8569 10024 13676 10026
rect 8569 9968 8574 10024
rect 8630 9968 13676 10024
rect 8569 9966 13676 9968
rect 8569 9963 8635 9966
rect 13670 9964 13676 9966
rect 13740 10026 13746 10028
rect 14406 10026 14412 10028
rect 13740 9966 14412 10026
rect 13740 9964 13746 9966
rect 14406 9964 14412 9966
rect 14476 9964 14482 10028
rect 19006 9964 19012 10028
rect 19076 10026 19082 10028
rect 20110 10026 20116 10028
rect 19076 9966 20116 10026
rect 19076 9964 19082 9966
rect 20110 9964 20116 9966
rect 20180 10026 20186 10028
rect 20253 10026 20319 10029
rect 20180 10024 20319 10026
rect 20180 9968 20258 10024
rect 20314 9968 20319 10024
rect 20180 9966 20319 9968
rect 20180 9964 20186 9966
rect 20253 9963 20319 9966
rect 20486 9966 22202 10026
rect 18689 9890 18755 9893
rect 20486 9890 20546 9966
rect 18689 9888 20546 9890
rect 18689 9832 18694 9888
rect 18750 9832 20546 9888
rect 18689 9830 20546 9832
rect 22142 9920 22202 9966
rect 22142 9830 23000 9920
rect 18689 9827 18755 9830
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 22200 9800 23000 9830
rect 21738 9759 22054 9760
rect 14457 9754 14523 9757
rect 14774 9754 14780 9756
rect 14457 9752 14780 9754
rect 14457 9696 14462 9752
rect 14518 9696 14780 9752
rect 14457 9694 14780 9696
rect 14457 9691 14523 9694
rect 14774 9692 14780 9694
rect 14844 9692 14850 9756
rect 9305 9618 9371 9621
rect 12157 9620 12223 9621
rect 9438 9618 9444 9620
rect 9305 9616 9444 9618
rect 9305 9560 9310 9616
rect 9366 9560 9444 9616
rect 9305 9558 9444 9560
rect 9305 9555 9371 9558
rect 9438 9556 9444 9558
rect 9508 9556 9514 9620
rect 12157 9618 12204 9620
rect 12112 9616 12204 9618
rect 12112 9560 12162 9616
rect 12112 9558 12204 9560
rect 12157 9556 12204 9558
rect 12268 9556 12274 9620
rect 12801 9618 12867 9621
rect 12934 9618 12940 9620
rect 12801 9616 12940 9618
rect 12801 9560 12806 9616
rect 12862 9560 12940 9616
rect 12801 9558 12940 9560
rect 12157 9555 12223 9556
rect 12801 9555 12867 9558
rect 12934 9556 12940 9558
rect 13004 9556 13010 9620
rect 14917 9618 14983 9621
rect 15142 9618 15148 9620
rect 14917 9616 15148 9618
rect 14917 9560 14922 9616
rect 14978 9560 15148 9616
rect 14917 9558 15148 9560
rect 14917 9555 14983 9558
rect 15142 9556 15148 9558
rect 15212 9556 15218 9620
rect 16941 9618 17007 9621
rect 18873 9620 18939 9621
rect 17350 9618 17356 9620
rect 16941 9616 17356 9618
rect 16941 9560 16946 9616
rect 17002 9560 17356 9616
rect 16941 9558 17356 9560
rect 16941 9555 17007 9558
rect 17350 9556 17356 9558
rect 17420 9556 17426 9620
rect 18822 9618 18828 9620
rect 18782 9558 18828 9618
rect 18892 9616 18939 9620
rect 18934 9560 18939 9616
rect 18822 9556 18828 9558
rect 18892 9556 18939 9560
rect 18873 9555 18939 9556
rect 7966 9420 7972 9484
rect 8036 9482 8042 9484
rect 9857 9482 9923 9485
rect 15101 9482 15167 9485
rect 8036 9480 15167 9482
rect 8036 9424 9862 9480
rect 9918 9424 15106 9480
rect 15162 9424 15167 9480
rect 8036 9422 15167 9424
rect 8036 9420 8042 9422
rect 9857 9419 9923 9422
rect 15101 9419 15167 9422
rect 17953 9482 18019 9485
rect 22200 9482 23000 9512
rect 17953 9480 23000 9482
rect 17953 9424 17958 9480
rect 18014 9424 23000 9480
rect 17953 9422 23000 9424
rect 17953 9419 18019 9422
rect 22200 9392 23000 9422
rect 11789 9346 11855 9349
rect 12525 9346 12591 9349
rect 11789 9344 12591 9346
rect 11789 9288 11794 9344
rect 11850 9288 12530 9344
rect 12586 9288 12591 9344
rect 11789 9286 12591 9288
rect 11789 9283 11855 9286
rect 12525 9283 12591 9286
rect 3545 9280 3861 9281
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 4613 9074 4679 9077
rect 14181 9074 14247 9077
rect 4613 9072 14247 9074
rect 4613 9016 4618 9072
rect 4674 9016 14186 9072
rect 14242 9016 14247 9072
rect 4613 9014 14247 9016
rect 4613 9011 4679 9014
rect 14181 9011 14247 9014
rect 17401 9074 17467 9077
rect 22200 9074 23000 9104
rect 17401 9072 23000 9074
rect 17401 9016 17406 9072
rect 17462 9016 23000 9072
rect 17401 9014 23000 9016
rect 17401 9011 17467 9014
rect 22200 8984 23000 9014
rect 15561 8804 15627 8805
rect 15510 8740 15516 8804
rect 15580 8802 15627 8804
rect 15580 8800 15672 8802
rect 15622 8744 15672 8800
rect 15580 8742 15672 8744
rect 15580 8740 15627 8742
rect 15518 8739 15627 8740
rect 6144 8736 6460 8737
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 13537 8668 13603 8669
rect 13486 8604 13492 8668
rect 13556 8666 13603 8668
rect 15193 8666 15259 8669
rect 15518 8666 15578 8739
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 21738 8671 22054 8672
rect 20253 8668 20319 8669
rect 20253 8666 20300 8668
rect 13556 8664 13648 8666
rect 13598 8608 13648 8664
rect 13556 8606 13648 8608
rect 15193 8664 15578 8666
rect 15193 8608 15198 8664
rect 15254 8608 15578 8664
rect 15193 8606 15578 8608
rect 20208 8664 20300 8666
rect 20208 8608 20258 8664
rect 20208 8606 20300 8608
rect 13556 8604 13603 8606
rect 13537 8603 13603 8604
rect 15193 8603 15259 8606
rect 20253 8604 20300 8606
rect 20364 8604 20370 8668
rect 22200 8666 23000 8696
rect 20253 8603 20319 8604
rect 22142 8576 23000 8666
rect 13813 8530 13879 8533
rect 16982 8530 16988 8532
rect 13813 8528 16988 8530
rect 13813 8472 13818 8528
rect 13874 8472 16988 8528
rect 13813 8470 16988 8472
rect 13813 8467 13879 8470
rect 16982 8468 16988 8470
rect 17052 8468 17058 8532
rect 19885 8530 19951 8533
rect 22142 8530 22202 8576
rect 19885 8528 22202 8530
rect 19885 8472 19890 8528
rect 19946 8472 22202 8528
rect 19885 8470 22202 8472
rect 19885 8467 19951 8470
rect 9673 8394 9739 8397
rect 10685 8394 10751 8397
rect 9673 8392 10751 8394
rect 9673 8336 9678 8392
rect 9734 8336 10690 8392
rect 10746 8336 10751 8392
rect 9673 8334 10751 8336
rect 9673 8331 9739 8334
rect 10685 8331 10751 8334
rect 18689 8394 18755 8397
rect 19742 8394 19748 8396
rect 18689 8392 19748 8394
rect 18689 8336 18694 8392
rect 18750 8336 19748 8392
rect 18689 8334 19748 8336
rect 18689 8331 18755 8334
rect 19742 8332 19748 8334
rect 19812 8332 19818 8396
rect 10133 8258 10199 8261
rect 12341 8258 12407 8261
rect 10133 8256 12407 8258
rect 10133 8200 10138 8256
rect 10194 8200 12346 8256
rect 12402 8200 12407 8256
rect 10133 8198 12407 8200
rect 10133 8195 10199 8198
rect 12341 8195 12407 8198
rect 15929 8258 15995 8261
rect 16205 8258 16271 8261
rect 22200 8258 23000 8288
rect 15929 8256 16271 8258
rect 15929 8200 15934 8256
rect 15990 8200 16210 8256
rect 16266 8200 16271 8256
rect 15929 8198 16271 8200
rect 15929 8195 15995 8198
rect 16205 8195 16271 8198
rect 19566 8198 23000 8258
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 9622 8060 9628 8124
rect 9692 8122 9698 8124
rect 11881 8122 11947 8125
rect 13721 8124 13787 8125
rect 9692 8120 11947 8122
rect 9692 8064 11886 8120
rect 11942 8064 11947 8120
rect 9692 8062 11947 8064
rect 9692 8060 9698 8062
rect 11881 8059 11947 8062
rect 13670 8060 13676 8124
rect 13740 8122 13787 8124
rect 13740 8120 13832 8122
rect 13782 8064 13832 8120
rect 13740 8062 13832 8064
rect 13740 8060 13787 8062
rect 13721 8059 13787 8060
rect 12341 7986 12407 7989
rect 13445 7986 13511 7989
rect 12341 7984 13511 7986
rect 12341 7928 12346 7984
rect 12402 7928 13450 7984
rect 13506 7928 13511 7984
rect 12341 7926 13511 7928
rect 12341 7923 12407 7926
rect 13445 7923 13511 7926
rect 18965 7986 19031 7989
rect 19566 7986 19626 8198
rect 22200 8168 23000 8198
rect 18965 7984 19626 7986
rect 18965 7928 18970 7984
rect 19026 7928 19626 7984
rect 18965 7926 19626 7928
rect 18965 7923 19031 7926
rect 13261 7850 13327 7853
rect 18689 7850 18755 7853
rect 13261 7848 18755 7850
rect 13261 7792 13266 7848
rect 13322 7792 18694 7848
rect 18750 7792 18755 7848
rect 13261 7790 18755 7792
rect 13261 7787 13327 7790
rect 18689 7787 18755 7790
rect 20897 7850 20963 7853
rect 22200 7850 23000 7880
rect 20897 7848 23000 7850
rect 20897 7792 20902 7848
rect 20958 7792 23000 7848
rect 20897 7790 23000 7792
rect 20897 7787 20963 7790
rect 22200 7760 23000 7790
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 18321 7578 18387 7581
rect 18321 7576 20914 7578
rect 18321 7520 18326 7576
rect 18382 7520 20914 7576
rect 18321 7518 20914 7520
rect 18321 7515 18387 7518
rect 10501 7442 10567 7445
rect 20713 7442 20779 7445
rect 10501 7440 20779 7442
rect 10501 7384 10506 7440
rect 10562 7384 20718 7440
rect 20774 7384 20779 7440
rect 10501 7382 20779 7384
rect 20854 7442 20914 7518
rect 22200 7442 23000 7472
rect 20854 7382 23000 7442
rect 10501 7379 10567 7382
rect 20713 7379 20779 7382
rect 22200 7352 23000 7382
rect 5901 7308 5967 7309
rect 5901 7304 5948 7308
rect 6012 7306 6018 7308
rect 18045 7306 18111 7309
rect 19609 7306 19675 7309
rect 5901 7248 5906 7304
rect 5901 7244 5948 7248
rect 6012 7246 6058 7306
rect 15150 7304 19675 7306
rect 15150 7248 18050 7304
rect 18106 7248 19614 7304
rect 19670 7248 19675 7304
rect 15150 7246 19675 7248
rect 6012 7244 6018 7246
rect 5901 7243 5967 7244
rect 3545 7104 3861 7105
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 8150 6972 8156 7036
rect 8220 7034 8226 7036
rect 8385 7034 8451 7037
rect 8220 7032 8451 7034
rect 8220 6976 8390 7032
rect 8446 6976 8451 7032
rect 8220 6974 8451 6976
rect 8220 6972 8226 6974
rect 8385 6971 8451 6974
rect 11973 7034 12039 7037
rect 13537 7034 13603 7037
rect 11973 7032 13603 7034
rect 11973 6976 11978 7032
rect 12034 6976 13542 7032
rect 13598 6976 13603 7032
rect 11973 6974 13603 6976
rect 11973 6971 12039 6974
rect 13537 6971 13603 6974
rect 4521 6898 4587 6901
rect 5349 6898 5415 6901
rect 11145 6900 11211 6901
rect 4521 6896 10978 6898
rect 4521 6840 4526 6896
rect 4582 6840 5354 6896
rect 5410 6840 10978 6896
rect 4521 6838 10978 6840
rect 4521 6835 4587 6838
rect 5349 6835 5415 6838
rect 10918 6762 10978 6838
rect 11094 6836 11100 6900
rect 11164 6898 11211 6900
rect 15150 6898 15210 7246
rect 18045 7243 18111 7246
rect 19609 7243 19675 7246
rect 18137 7172 18203 7173
rect 18086 7108 18092 7172
rect 18156 7170 18203 7172
rect 18156 7168 18248 7170
rect 18198 7112 18248 7168
rect 18156 7110 18248 7112
rect 18156 7108 18203 7110
rect 18137 7107 18203 7108
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 19139 7039 19455 7040
rect 22200 7034 23000 7064
rect 19566 6974 23000 7034
rect 11164 6896 11256 6898
rect 11206 6840 11256 6896
rect 11164 6838 11256 6840
rect 12390 6838 15210 6898
rect 19241 6898 19307 6901
rect 19566 6898 19626 6974
rect 22200 6944 23000 6974
rect 19241 6896 19626 6898
rect 19241 6840 19246 6896
rect 19302 6840 19626 6896
rect 19241 6838 19626 6840
rect 11164 6836 11211 6838
rect 11145 6835 11211 6836
rect 12390 6762 12450 6838
rect 19241 6835 19307 6838
rect 10918 6702 12450 6762
rect 12525 6762 12591 6765
rect 13169 6762 13235 6765
rect 12525 6760 13235 6762
rect 12525 6704 12530 6760
rect 12586 6704 13174 6760
rect 13230 6704 13235 6760
rect 12525 6702 13235 6704
rect 12525 6699 12591 6702
rect 13169 6699 13235 6702
rect 13445 6762 13511 6765
rect 16113 6762 16179 6765
rect 13445 6760 16179 6762
rect 13445 6704 13450 6760
rect 13506 6704 16118 6760
rect 16174 6704 16179 6760
rect 13445 6702 16179 6704
rect 13445 6699 13511 6702
rect 16113 6699 16179 6702
rect 18873 6762 18939 6765
rect 18873 6760 22202 6762
rect 18873 6704 18878 6760
rect 18934 6704 22202 6760
rect 18873 6702 22202 6704
rect 18873 6699 18939 6702
rect 22142 6656 22202 6702
rect 22142 6566 23000 6656
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 22200 6536 23000 6566
rect 21738 6495 22054 6496
rect 12709 6490 12775 6493
rect 17033 6490 17099 6493
rect 12709 6488 15578 6490
rect 12709 6432 12714 6488
rect 12770 6432 15578 6488
rect 12709 6430 15578 6432
rect 12709 6427 12775 6430
rect 9213 6354 9279 6357
rect 15285 6356 15351 6357
rect 15285 6354 15332 6356
rect 9213 6352 13370 6354
rect 9213 6296 9218 6352
rect 9274 6296 13370 6352
rect 9213 6294 13370 6296
rect 15240 6352 15332 6354
rect 15240 6296 15290 6352
rect 15240 6294 15332 6296
rect 9213 6291 9279 6294
rect 12157 6218 12223 6221
rect 12801 6218 12867 6221
rect 12157 6216 12867 6218
rect 12157 6160 12162 6216
rect 12218 6160 12806 6216
rect 12862 6160 12867 6216
rect 12157 6158 12867 6160
rect 12157 6155 12223 6158
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 0 5810 800 5840
rect 3509 5810 3575 5813
rect 0 5808 3575 5810
rect 0 5752 3514 5808
rect 3570 5752 3575 5808
rect 0 5750 3575 5752
rect 0 5720 800 5750
rect 3509 5747 3575 5750
rect 12390 5677 12450 6158
rect 12801 6155 12867 6158
rect 12341 5672 12450 5677
rect 12341 5616 12346 5672
rect 12402 5616 12450 5672
rect 12341 5614 12450 5616
rect 13310 5674 13370 6294
rect 15285 6292 15332 6294
rect 15396 6292 15402 6356
rect 15518 6354 15578 6430
rect 17033 6488 21098 6490
rect 17033 6432 17038 6488
rect 17094 6432 21098 6488
rect 17033 6430 21098 6432
rect 17033 6427 17099 6430
rect 20713 6354 20779 6357
rect 20897 6354 20963 6357
rect 15518 6352 20963 6354
rect 15518 6296 20718 6352
rect 20774 6296 20902 6352
rect 20958 6296 20963 6352
rect 15518 6294 20963 6296
rect 15285 6291 15351 6292
rect 20713 6291 20779 6294
rect 20897 6291 20963 6294
rect 13537 6218 13603 6221
rect 17769 6218 17835 6221
rect 13537 6216 17835 6218
rect 13537 6160 13542 6216
rect 13598 6160 17774 6216
rect 17830 6160 17835 6216
rect 13537 6158 17835 6160
rect 21038 6218 21098 6430
rect 22200 6218 23000 6248
rect 21038 6158 23000 6218
rect 13537 6155 13603 6158
rect 17769 6155 17835 6158
rect 22200 6128 23000 6158
rect 15193 6082 15259 6085
rect 18413 6082 18479 6085
rect 15193 6080 18479 6082
rect 15193 6024 15198 6080
rect 15254 6024 18418 6080
rect 18474 6024 18479 6080
rect 15193 6022 18479 6024
rect 15193 6019 15259 6022
rect 18413 6019 18479 6022
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 17166 5884 17172 5948
rect 17236 5946 17242 5948
rect 17401 5946 17467 5949
rect 17236 5944 17467 5946
rect 17236 5888 17406 5944
rect 17462 5888 17467 5944
rect 17236 5886 17467 5888
rect 17236 5884 17242 5886
rect 17401 5883 17467 5886
rect 13813 5810 13879 5813
rect 17033 5810 17099 5813
rect 17493 5812 17559 5813
rect 17493 5810 17540 5812
rect 13813 5808 17099 5810
rect 13813 5752 13818 5808
rect 13874 5752 17038 5808
rect 17094 5752 17099 5808
rect 13813 5750 17099 5752
rect 17448 5808 17540 5810
rect 17448 5752 17498 5808
rect 17448 5750 17540 5752
rect 13813 5747 13879 5750
rect 17033 5747 17099 5750
rect 17493 5748 17540 5750
rect 17604 5748 17610 5812
rect 17953 5810 18019 5813
rect 22200 5810 23000 5840
rect 17953 5808 23000 5810
rect 17953 5752 17958 5808
rect 18014 5752 23000 5808
rect 17953 5750 23000 5752
rect 17493 5747 17559 5748
rect 17953 5747 18019 5750
rect 22200 5720 23000 5750
rect 20897 5674 20963 5677
rect 13310 5672 20963 5674
rect 13310 5616 20902 5672
rect 20958 5616 20963 5672
rect 13310 5614 20963 5616
rect 12341 5611 12407 5614
rect 20897 5611 20963 5614
rect 20161 5540 20227 5541
rect 20110 5538 20116 5540
rect 20070 5478 20116 5538
rect 20180 5536 20227 5540
rect 20222 5480 20227 5536
rect 20110 5476 20116 5478
rect 20180 5476 20227 5480
rect 20161 5475 20227 5476
rect 6144 5472 6460 5473
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 21738 5407 22054 5408
rect 15837 5404 15903 5405
rect 15837 5402 15884 5404
rect 15792 5400 15884 5402
rect 15792 5344 15842 5400
rect 15792 5342 15884 5344
rect 15837 5340 15884 5342
rect 15948 5340 15954 5404
rect 22200 5402 23000 5432
rect 15837 5339 15903 5340
rect 22142 5312 23000 5402
rect 13905 5266 13971 5269
rect 19701 5266 19767 5269
rect 22142 5266 22202 5312
rect 13905 5264 19767 5266
rect 13905 5208 13910 5264
rect 13966 5208 19706 5264
rect 19762 5208 19767 5264
rect 13905 5206 19767 5208
rect 13905 5203 13971 5206
rect 19701 5203 19767 5206
rect 21958 5206 22202 5266
rect 10593 5130 10659 5133
rect 17953 5130 18019 5133
rect 10593 5128 18019 5130
rect 10593 5072 10598 5128
rect 10654 5072 17958 5128
rect 18014 5072 18019 5128
rect 10593 5070 18019 5072
rect 10593 5067 10659 5070
rect 17953 5067 18019 5070
rect 18413 5130 18479 5133
rect 18689 5130 18755 5133
rect 21958 5130 22018 5206
rect 18413 5128 22018 5130
rect 18413 5072 18418 5128
rect 18474 5072 18694 5128
rect 18750 5072 22018 5128
rect 18413 5070 22018 5072
rect 18413 5067 18479 5070
rect 18689 5067 18755 5070
rect 14365 4994 14431 4997
rect 18137 4994 18203 4997
rect 14365 4992 18203 4994
rect 14365 4936 14370 4992
rect 14426 4936 18142 4992
rect 18198 4936 18203 4992
rect 14365 4934 18203 4936
rect 14365 4931 14431 4934
rect 18137 4931 18203 4934
rect 21081 4994 21147 4997
rect 22200 4994 23000 5024
rect 21081 4992 23000 4994
rect 21081 4936 21086 4992
rect 21142 4936 23000 4992
rect 21081 4934 23000 4936
rect 21081 4931 21147 4934
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 22200 4904 23000 4934
rect 19139 4863 19455 4864
rect 10409 4722 10475 4725
rect 20253 4722 20319 4725
rect 10409 4720 20319 4722
rect 10409 4664 10414 4720
rect 10470 4664 20258 4720
rect 20314 4664 20319 4720
rect 10409 4662 20319 4664
rect 10409 4659 10475 4662
rect 20253 4659 20319 4662
rect 17953 4586 18019 4589
rect 19558 4586 19564 4588
rect 16254 4584 19564 4586
rect 16254 4528 17958 4584
rect 18014 4528 19564 4584
rect 16254 4526 19564 4528
rect 16254 4450 16314 4526
rect 17953 4523 18019 4526
rect 19558 4524 19564 4526
rect 19628 4524 19634 4588
rect 20621 4586 20687 4589
rect 21173 4586 21239 4589
rect 22200 4586 23000 4616
rect 20621 4584 23000 4586
rect 20621 4528 20626 4584
rect 20682 4528 21178 4584
rect 21234 4528 23000 4584
rect 20621 4526 23000 4528
rect 20621 4523 20687 4526
rect 21173 4523 21239 4526
rect 22200 4496 23000 4526
rect 12390 4390 16314 4450
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 10593 4178 10659 4181
rect 12390 4178 12450 4390
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 18597 4314 18663 4317
rect 18597 4312 20178 4314
rect 18597 4256 18602 4312
rect 18658 4256 20178 4312
rect 18597 4254 20178 4256
rect 18597 4251 18663 4254
rect 10593 4176 12450 4178
rect 10593 4120 10598 4176
rect 10654 4120 12450 4176
rect 10593 4118 12450 4120
rect 15837 4178 15903 4181
rect 19885 4178 19951 4181
rect 15837 4176 19951 4178
rect 15837 4120 15842 4176
rect 15898 4120 19890 4176
rect 19946 4120 19951 4176
rect 15837 4118 19951 4120
rect 20118 4178 20178 4254
rect 22200 4178 23000 4208
rect 20118 4118 23000 4178
rect 10593 4115 10659 4118
rect 15837 4115 15903 4118
rect 19885 4115 19951 4118
rect 22200 4088 23000 4118
rect 4797 4042 4863 4045
rect 10869 4042 10935 4045
rect 4797 4040 10935 4042
rect 4797 3984 4802 4040
rect 4858 3984 10874 4040
rect 10930 3984 10935 4040
rect 4797 3982 10935 3984
rect 4797 3979 4863 3982
rect 10869 3979 10935 3982
rect 11053 4042 11119 4045
rect 16849 4042 16915 4045
rect 11053 4040 16915 4042
rect 11053 3984 11058 4040
rect 11114 3984 16854 4040
rect 16910 3984 16915 4040
rect 11053 3982 16915 3984
rect 11053 3979 11119 3982
rect 16849 3979 16915 3982
rect 18137 4042 18203 4045
rect 19977 4042 20043 4045
rect 18137 4040 20043 4042
rect 18137 3984 18142 4040
rect 18198 3984 19982 4040
rect 20038 3984 20043 4040
rect 18137 3982 20043 3984
rect 18137 3979 18203 3982
rect 19977 3979 20043 3982
rect 6545 3906 6611 3909
rect 6678 3906 6684 3908
rect 6545 3904 6684 3906
rect 6545 3848 6550 3904
rect 6606 3848 6684 3904
rect 6545 3846 6684 3848
rect 6545 3843 6611 3846
rect 6678 3844 6684 3846
rect 6748 3844 6754 3908
rect 9438 3844 9444 3908
rect 9508 3906 9514 3908
rect 9765 3906 9831 3909
rect 9508 3904 9831 3906
rect 9508 3848 9770 3904
rect 9826 3848 9831 3904
rect 9508 3846 9831 3848
rect 9508 3844 9514 3846
rect 9765 3843 9831 3846
rect 3545 3840 3861 3841
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 19139 3775 19455 3776
rect 14917 3770 14983 3773
rect 17953 3770 18019 3773
rect 22200 3770 23000 3800
rect 14917 3768 18019 3770
rect 14917 3712 14922 3768
rect 14978 3712 17958 3768
rect 18014 3712 18019 3768
rect 14917 3710 18019 3712
rect 14917 3707 14983 3710
rect 17953 3707 18019 3710
rect 19566 3710 23000 3770
rect 9121 3634 9187 3637
rect 18965 3634 19031 3637
rect 9121 3632 19031 3634
rect 9121 3576 9126 3632
rect 9182 3576 18970 3632
rect 19026 3576 19031 3632
rect 9121 3574 19031 3576
rect 9121 3571 9187 3574
rect 18965 3571 19031 3574
rect 9806 3436 9812 3500
rect 9876 3498 9882 3500
rect 15745 3498 15811 3501
rect 18086 3498 18092 3500
rect 9876 3496 15811 3498
rect 9876 3440 15750 3496
rect 15806 3440 15811 3496
rect 9876 3438 15811 3440
rect 9876 3436 9882 3438
rect 15745 3435 15811 3438
rect 16254 3438 18092 3498
rect 16254 3362 16314 3438
rect 18086 3436 18092 3438
rect 18156 3498 18162 3500
rect 18781 3498 18847 3501
rect 18156 3496 18847 3498
rect 18156 3440 18786 3496
rect 18842 3440 18847 3496
rect 18156 3438 18847 3440
rect 18156 3436 18162 3438
rect 18781 3435 18847 3438
rect 12390 3302 16314 3362
rect 18321 3362 18387 3365
rect 19566 3362 19626 3710
rect 22200 3680 23000 3710
rect 18321 3360 19626 3362
rect 18321 3304 18326 3360
rect 18382 3304 19626 3360
rect 18321 3302 19626 3304
rect 21038 3438 22202 3498
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 9857 3228 9923 3229
rect 9806 3164 9812 3228
rect 9876 3226 9923 3228
rect 12390 3226 12450 3302
rect 18321 3299 18387 3302
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 9876 3224 9968 3226
rect 9918 3168 9968 3224
rect 9876 3166 9968 3168
rect 11838 3166 12450 3226
rect 9876 3164 9923 3166
rect 9857 3163 9923 3164
rect 1485 3090 1551 3093
rect 9622 3090 9628 3092
rect 1485 3088 9628 3090
rect 1485 3032 1490 3088
rect 1546 3032 9628 3088
rect 1485 3030 9628 3032
rect 1485 3027 1551 3030
rect 9622 3028 9628 3030
rect 9692 3028 9698 3092
rect 9765 3090 9831 3093
rect 11838 3090 11898 3166
rect 16982 3164 16988 3228
rect 17052 3226 17058 3228
rect 20897 3226 20963 3229
rect 17052 3224 20963 3226
rect 17052 3168 20902 3224
rect 20958 3168 20963 3224
rect 17052 3166 20963 3168
rect 17052 3164 17058 3166
rect 20897 3163 20963 3166
rect 9765 3088 11898 3090
rect 9765 3032 9770 3088
rect 9826 3032 11898 3088
rect 9765 3030 11898 3032
rect 12065 3090 12131 3093
rect 17861 3090 17927 3093
rect 12065 3088 17927 3090
rect 12065 3032 12070 3088
rect 12126 3032 17866 3088
rect 17922 3032 17927 3088
rect 12065 3030 17927 3032
rect 9765 3027 9831 3030
rect 12065 3027 12131 3030
rect 17861 3027 17927 3030
rect 18229 3090 18295 3093
rect 21038 3090 21098 3438
rect 22142 3392 22202 3438
rect 22142 3302 23000 3392
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 22200 3272 23000 3302
rect 21738 3231 22054 3232
rect 18229 3088 21098 3090
rect 18229 3032 18234 3088
rect 18290 3032 21098 3088
rect 18229 3030 21098 3032
rect 18229 3027 18295 3030
rect 11053 2954 11119 2957
rect 14181 2954 14247 2957
rect 11053 2952 14247 2954
rect 11053 2896 11058 2952
rect 11114 2896 14186 2952
rect 14242 2896 14247 2952
rect 11053 2894 14247 2896
rect 11053 2891 11119 2894
rect 14181 2891 14247 2894
rect 15745 2954 15811 2957
rect 19333 2954 19399 2957
rect 15745 2952 19399 2954
rect 15745 2896 15750 2952
rect 15806 2896 19338 2952
rect 19394 2896 19399 2952
rect 15745 2894 19399 2896
rect 15745 2891 15811 2894
rect 19333 2891 19399 2894
rect 20897 2954 20963 2957
rect 22200 2954 23000 2984
rect 20897 2952 23000 2954
rect 20897 2896 20902 2952
rect 20958 2896 23000 2952
rect 20897 2894 23000 2896
rect 20897 2891 20963 2894
rect 22200 2864 23000 2894
rect 3545 2752 3861 2753
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 19149 2546 19215 2549
rect 22200 2546 23000 2576
rect 19149 2544 23000 2546
rect 19149 2488 19154 2544
rect 19210 2488 23000 2544
rect 19149 2486 23000 2488
rect 19149 2483 19215 2486
rect 22200 2456 23000 2486
rect 6144 2208 6460 2209
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 21738 2143 22054 2144
rect 22200 2138 23000 2168
rect 22142 2048 23000 2138
rect 18873 2002 18939 2005
rect 22142 2002 22202 2048
rect 18873 2000 22202 2002
rect 18873 1944 18878 2000
rect 18934 1944 22202 2000
rect 18873 1942 22202 1944
rect 18873 1939 18939 1942
rect 20345 1730 20411 1733
rect 22200 1730 23000 1760
rect 20345 1728 23000 1730
rect 20345 1672 20350 1728
rect 20406 1672 23000 1728
rect 20345 1670 23000 1672
rect 20345 1667 20411 1670
rect 22200 1640 23000 1670
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 5948 20164 6012 20228
rect 14412 20164 14476 20228
rect 17356 20164 17420 20228
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 12204 19892 12268 19956
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 9444 18124 9508 18188
rect 9812 18048 9876 18052
rect 9812 17992 9826 18048
rect 9826 17992 9876 18048
rect 9812 17988 9876 17992
rect 20300 17988 20364 18052
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 10364 17716 10428 17780
rect 13676 17580 13740 17644
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 15884 17172 15948 17236
rect 15516 17036 15580 17100
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 12940 16492 13004 16556
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 13124 16084 13188 16148
rect 14780 15948 14844 16012
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 6684 15404 6748 15468
rect 17172 15404 17236 15468
rect 11836 15268 11900 15332
rect 15148 15268 15212 15332
rect 19748 15268 19812 15332
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 19012 14860 19076 14924
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 8156 14044 8220 14108
rect 15332 13772 15396 13836
rect 18828 13832 18892 13836
rect 18828 13776 18878 13832
rect 18878 13776 18892 13832
rect 18828 13772 18892 13776
rect 17540 13636 17604 13700
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 11100 13364 11164 13428
rect 17540 13228 17604 13292
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 7972 12820 8036 12884
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 19932 12684 19996 12748
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 8156 11792 8220 11796
rect 8156 11736 8206 11792
rect 8206 11736 8220 11792
rect 8156 11732 8220 11736
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 8156 11052 8220 11116
rect 19564 11052 19628 11116
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 10364 10780 10428 10844
rect 11836 10780 11900 10844
rect 6684 10508 6748 10572
rect 9444 10508 9508 10572
rect 19932 10508 19996 10572
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 13124 10236 13188 10300
rect 13676 9964 13740 10028
rect 14412 9964 14476 10028
rect 19012 9964 19076 10028
rect 20116 9964 20180 10028
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 14780 9692 14844 9756
rect 9444 9556 9508 9620
rect 12204 9616 12268 9620
rect 12204 9560 12218 9616
rect 12218 9560 12268 9616
rect 12204 9556 12268 9560
rect 12940 9556 13004 9620
rect 15148 9556 15212 9620
rect 17356 9556 17420 9620
rect 18828 9616 18892 9620
rect 18828 9560 18878 9616
rect 18878 9560 18892 9616
rect 18828 9556 18892 9560
rect 7972 9420 8036 9484
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 15516 8800 15580 8804
rect 15516 8744 15566 8800
rect 15566 8744 15580 8800
rect 15516 8740 15580 8744
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 13492 8664 13556 8668
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 13492 8608 13542 8664
rect 13542 8608 13556 8664
rect 13492 8604 13556 8608
rect 20300 8664 20364 8668
rect 20300 8608 20314 8664
rect 20314 8608 20364 8664
rect 20300 8604 20364 8608
rect 16988 8468 17052 8532
rect 19748 8332 19812 8396
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 9628 8060 9692 8124
rect 13676 8120 13740 8124
rect 13676 8064 13726 8120
rect 13726 8064 13740 8120
rect 13676 8060 13740 8064
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 5948 7304 6012 7308
rect 5948 7248 5962 7304
rect 5962 7248 6012 7304
rect 5948 7244 6012 7248
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 8156 6972 8220 7036
rect 11100 6896 11164 6900
rect 18092 7168 18156 7172
rect 18092 7112 18142 7168
rect 18142 7112 18156 7168
rect 18092 7108 18156 7112
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 11100 6840 11150 6896
rect 11150 6840 11164 6896
rect 11100 6836 11164 6840
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 15332 6352 15396 6356
rect 15332 6296 15346 6352
rect 15346 6296 15396 6352
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 15332 6292 15396 6296
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 17172 5884 17236 5948
rect 17540 5808 17604 5812
rect 17540 5752 17554 5808
rect 17554 5752 17604 5808
rect 17540 5748 17604 5752
rect 20116 5536 20180 5540
rect 20116 5480 20166 5536
rect 20166 5480 20180 5536
rect 20116 5476 20180 5480
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 15884 5400 15948 5404
rect 15884 5344 15898 5400
rect 15898 5344 15948 5400
rect 15884 5340 15948 5344
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 19564 4524 19628 4588
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 6684 3844 6748 3908
rect 9444 3844 9508 3908
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 9812 3436 9876 3500
rect 18092 3436 18156 3500
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 9812 3224 9876 3228
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 9812 3168 9862 3224
rect 9862 3168 9876 3224
rect 9812 3164 9876 3168
rect 9628 3028 9692 3092
rect 16988 3164 17052 3228
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 5947 20228 6013 20229
rect 5947 20164 5948 20228
rect 6012 20164 6013 20228
rect 5947 20163 6013 20164
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 5950 7309 6010 20163
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 13939 20160 14259 20720
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 14411 20228 14477 20229
rect 14411 20164 14412 20228
rect 14476 20164 14477 20228
rect 14411 20163 14477 20164
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 12203 19956 12269 19957
rect 12203 19892 12204 19956
rect 12268 19892 12269 19956
rect 12203 19891 12269 19892
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 9443 18188 9509 18189
rect 9443 18124 9444 18188
rect 9508 18124 9509 18188
rect 9443 18123 9509 18124
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 6683 15468 6749 15469
rect 6683 15404 6684 15468
rect 6748 15404 6749 15468
rect 6683 15403 6749 15404
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6686 10573 6746 15403
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8155 14108 8221 14109
rect 8155 14044 8156 14108
rect 8220 14044 8221 14108
rect 8155 14043 8221 14044
rect 7971 12884 8037 12885
rect 7971 12820 7972 12884
rect 8036 12820 8037 12884
rect 7971 12819 8037 12820
rect 6683 10572 6749 10573
rect 6683 10508 6684 10572
rect 6748 10508 6749 10572
rect 6683 10507 6749 10508
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 5947 7308 6013 7309
rect 5947 7244 5948 7308
rect 6012 7244 6013 7308
rect 5947 7243 6013 7244
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6686 3909 6746 10507
rect 7974 9485 8034 12819
rect 8158 11797 8218 14043
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8155 11796 8221 11797
rect 8155 11732 8156 11796
rect 8220 11732 8221 11796
rect 8155 11731 8221 11732
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8155 11116 8221 11117
rect 8155 11052 8156 11116
rect 8220 11052 8221 11116
rect 8155 11051 8221 11052
rect 7971 9484 8037 9485
rect 7971 9420 7972 9484
rect 8036 9420 8037 9484
rect 7971 9419 8037 9420
rect 8158 7037 8218 11051
rect 8741 10368 9061 11392
rect 9446 10573 9506 18123
rect 9811 18052 9877 18053
rect 9811 17988 9812 18052
rect 9876 17988 9877 18052
rect 9811 17987 9877 17988
rect 9443 10572 9509 10573
rect 9443 10508 9444 10572
rect 9508 10508 9509 10572
rect 9443 10507 9509 10508
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 9446 9621 9506 10507
rect 9443 9620 9509 9621
rect 9443 9556 9444 9620
rect 9508 9556 9509 9620
rect 9443 9555 9509 9556
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8155 7036 8221 7037
rect 8155 6972 8156 7036
rect 8220 6972 8221 7036
rect 8155 6971 8221 6972
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 6683 3908 6749 3909
rect 6683 3844 6684 3908
rect 6748 3844 6749 3908
rect 6683 3843 6749 3844
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 3840 9061 4864
rect 9446 3909 9506 9555
rect 9627 8124 9693 8125
rect 9627 8060 9628 8124
rect 9692 8060 9693 8124
rect 9627 8059 9693 8060
rect 9443 3908 9509 3909
rect 9443 3844 9444 3908
rect 9508 3844 9509 3908
rect 9443 3843 9509 3844
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 2752 9061 3776
rect 9630 3093 9690 8059
rect 9814 3501 9874 17987
rect 10363 17780 10429 17781
rect 10363 17716 10364 17780
rect 10428 17716 10429 17780
rect 10363 17715 10429 17716
rect 10366 10845 10426 17715
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11835 15332 11901 15333
rect 11835 15268 11836 15332
rect 11900 15268 11901 15332
rect 11835 15267 11901 15268
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11099 13428 11165 13429
rect 11099 13364 11100 13428
rect 11164 13364 11165 13428
rect 11099 13363 11165 13364
rect 10363 10844 10429 10845
rect 10363 10780 10364 10844
rect 10428 10780 10429 10844
rect 10363 10779 10429 10780
rect 11102 6901 11162 13363
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11838 10845 11898 15267
rect 11835 10844 11901 10845
rect 11835 10780 11836 10844
rect 11900 10780 11901 10844
rect 11835 10779 11901 10780
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 12206 9621 12266 19891
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13675 17644 13741 17645
rect 13675 17580 13676 17644
rect 13740 17580 13741 17644
rect 13675 17579 13741 17580
rect 12939 16556 13005 16557
rect 12939 16492 12940 16556
rect 13004 16492 13005 16556
rect 12939 16491 13005 16492
rect 12942 9621 13002 16491
rect 13123 16148 13189 16149
rect 13123 16084 13124 16148
rect 13188 16084 13189 16148
rect 13123 16083 13189 16084
rect 13126 10301 13186 16083
rect 13678 12450 13738 17579
rect 13494 12390 13738 12450
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13123 10300 13189 10301
rect 13123 10236 13124 10300
rect 13188 10236 13189 10300
rect 13123 10235 13189 10236
rect 12203 9620 12269 9621
rect 12203 9556 12204 9620
rect 12268 9556 12269 9620
rect 12203 9555 12269 9556
rect 12939 9620 13005 9621
rect 12939 9556 12940 9620
rect 13004 9556 13005 9620
rect 12939 9555 13005 9556
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 13494 8669 13554 12390
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13675 10028 13741 10029
rect 13675 9964 13676 10028
rect 13740 9964 13741 10028
rect 13675 9963 13741 9964
rect 13491 8668 13557 8669
rect 13491 8604 13492 8668
rect 13556 8604 13557 8668
rect 13491 8603 13557 8604
rect 13678 8125 13738 9963
rect 13939 9280 14259 10304
rect 14414 10029 14474 20163
rect 16538 19616 16858 20640
rect 17355 20228 17421 20229
rect 17355 20164 17356 20228
rect 17420 20164 17421 20228
rect 17355 20163 17421 20164
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 15883 17236 15949 17237
rect 15883 17172 15884 17236
rect 15948 17172 15949 17236
rect 15883 17171 15949 17172
rect 15515 17100 15581 17101
rect 15515 17036 15516 17100
rect 15580 17036 15581 17100
rect 15515 17035 15581 17036
rect 14779 16012 14845 16013
rect 14779 15948 14780 16012
rect 14844 15948 14845 16012
rect 14779 15947 14845 15948
rect 14411 10028 14477 10029
rect 14411 9964 14412 10028
rect 14476 9964 14477 10028
rect 14411 9963 14477 9964
rect 14782 9757 14842 15947
rect 15147 15332 15213 15333
rect 15147 15268 15148 15332
rect 15212 15268 15213 15332
rect 15147 15267 15213 15268
rect 14779 9756 14845 9757
rect 14779 9692 14780 9756
rect 14844 9692 14845 9756
rect 14779 9691 14845 9692
rect 15150 9621 15210 15267
rect 15331 13836 15397 13837
rect 15331 13772 15332 13836
rect 15396 13772 15397 13836
rect 15331 13771 15397 13772
rect 15147 9620 15213 9621
rect 15147 9556 15148 9620
rect 15212 9556 15213 9620
rect 15147 9555 15213 9556
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13675 8124 13741 8125
rect 13675 8060 13676 8124
rect 13740 8060 13741 8124
rect 13675 8059 13741 8060
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11099 6900 11165 6901
rect 11099 6836 11100 6900
rect 11164 6836 11165 6900
rect 11099 6835 11165 6836
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 9811 3500 9877 3501
rect 9811 3436 9812 3500
rect 9876 3436 9877 3500
rect 9811 3435 9877 3436
rect 9814 3229 9874 3435
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 9811 3228 9877 3229
rect 9811 3164 9812 3228
rect 9876 3164 9877 3228
rect 9811 3163 9877 3164
rect 9627 3092 9693 3093
rect 9627 3028 9628 3092
rect 9692 3028 9693 3092
rect 9627 3027 9693 3028
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 15334 6357 15394 13771
rect 15518 8805 15578 17035
rect 15515 8804 15581 8805
rect 15515 8740 15516 8804
rect 15580 8740 15581 8804
rect 15515 8739 15581 8740
rect 15331 6356 15397 6357
rect 15331 6292 15332 6356
rect 15396 6292 15397 6356
rect 15331 6291 15397 6292
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 15886 5405 15946 17171
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 17171 15468 17237 15469
rect 17171 15404 17172 15468
rect 17236 15404 17237 15468
rect 17171 15403 17237 15404
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16987 8532 17053 8533
rect 16987 8468 16988 8532
rect 17052 8468 17053 8532
rect 16987 8467 17053 8468
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 15883 5404 15949 5405
rect 15883 5340 15884 5404
rect 15948 5340 15949 5404
rect 15883 5339 15949 5340
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16990 3229 17050 8467
rect 17174 5949 17234 15403
rect 17358 9621 17418 20163
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 20299 18052 20365 18053
rect 20299 17988 20300 18052
rect 20364 17988 20365 18052
rect 20299 17987 20365 17988
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19011 14924 19077 14925
rect 19011 14860 19012 14924
rect 19076 14860 19077 14924
rect 19011 14859 19077 14860
rect 18827 13836 18893 13837
rect 18827 13772 18828 13836
rect 18892 13772 18893 13836
rect 18827 13771 18893 13772
rect 17539 13700 17605 13701
rect 17539 13636 17540 13700
rect 17604 13636 17605 13700
rect 17539 13635 17605 13636
rect 17542 13293 17602 13635
rect 17539 13292 17605 13293
rect 17539 13228 17540 13292
rect 17604 13228 17605 13292
rect 17539 13227 17605 13228
rect 17355 9620 17421 9621
rect 17355 9556 17356 9620
rect 17420 9556 17421 9620
rect 17355 9555 17421 9556
rect 17171 5948 17237 5949
rect 17171 5884 17172 5948
rect 17236 5884 17237 5948
rect 17171 5883 17237 5884
rect 17542 5813 17602 13227
rect 18830 9621 18890 13771
rect 19014 10029 19074 14859
rect 19137 14720 19457 15744
rect 19747 15332 19813 15333
rect 19747 15268 19748 15332
rect 19812 15268 19813 15332
rect 19747 15267 19813 15268
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19563 11116 19629 11117
rect 19563 11052 19564 11116
rect 19628 11052 19629 11116
rect 19563 11051 19629 11052
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19011 10028 19077 10029
rect 19011 9964 19012 10028
rect 19076 9964 19077 10028
rect 19011 9963 19077 9964
rect 18827 9620 18893 9621
rect 18827 9556 18828 9620
rect 18892 9556 18893 9620
rect 18827 9555 18893 9556
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 18091 7172 18157 7173
rect 18091 7108 18092 7172
rect 18156 7108 18157 7172
rect 18091 7107 18157 7108
rect 17539 5812 17605 5813
rect 17539 5748 17540 5812
rect 17604 5748 17605 5812
rect 17539 5747 17605 5748
rect 18094 3501 18154 7107
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19566 4589 19626 11051
rect 19750 8397 19810 15267
rect 19931 12748 19997 12749
rect 19931 12684 19932 12748
rect 19996 12684 19997 12748
rect 19931 12683 19997 12684
rect 19934 10573 19994 12683
rect 19931 10572 19997 10573
rect 19931 10508 19932 10572
rect 19996 10508 19997 10572
rect 19931 10507 19997 10508
rect 20115 10028 20181 10029
rect 20115 9964 20116 10028
rect 20180 9964 20181 10028
rect 20115 9963 20181 9964
rect 19747 8396 19813 8397
rect 19747 8332 19748 8396
rect 19812 8332 19813 8396
rect 19747 8331 19813 8332
rect 20118 5541 20178 9963
rect 20302 8669 20362 17987
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 20299 8668 20365 8669
rect 20299 8604 20300 8668
rect 20364 8604 20365 8668
rect 20299 8603 20365 8604
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 20115 5540 20181 5541
rect 20115 5476 20116 5540
rect 20180 5476 20181 5540
rect 20115 5475 20181 5476
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 19563 4588 19629 4589
rect 19563 4524 19564 4588
rect 19628 4524 19629 4588
rect 19563 4523 19629 4524
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 18091 3500 18157 3501
rect 18091 3436 18092 3500
rect 18156 3436 18157 3500
rect 18091 3435 18157 3436
rect 16987 3228 17053 3229
rect 16987 3164 16988 3228
rect 17052 3164 17053 3228
rect 16987 3163 17053 3164
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13340 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1649977179
transform 1 0 11592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1649977179
transform 1 0 12512 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1649977179
transform -1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1649977179
transform 1 0 10672 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1649977179
transform -1 0 10304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1649977179
transform -1 0 20148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1649977179
transform -1 0 19780 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1649977179
transform -1 0 8924 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1649977179
transform 1 0 9936 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1649977179
transform 1 0 9844 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1649977179
transform -1 0 9936 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1649977179
transform -1 0 9568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1649977179
transform -1 0 10488 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1649977179
transform -1 0 5796 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1649977179
transform 1 0 5520 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1649977179
transform -1 0 5152 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1649977179
transform 1 0 5888 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1649977179
transform -1 0 12696 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1649977179
transform 1 0 13248 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1649977179
transform -1 0 12328 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1649977179
transform -1 0 13064 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1649977179
transform 1 0 14628 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1649977179
transform 1 0 12880 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1649977179
transform 1 0 11868 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1649977179
transform -1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1649977179
transform -1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7912 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7728 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19596 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 19412 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 17020 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15640 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15180 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 17480 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 18952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19596 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13248 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18584 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19320 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 21252 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 11868 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 8096 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 9016 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8648 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10672 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10672 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12512 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10948 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13064 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10580 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13616 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18124 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17572 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14536 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11776 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16928 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17940 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18124 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19596 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12880 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10764 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 8648 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12144 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13432 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16744 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10856 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15548 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12328 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13616 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14720 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17204 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12972 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12972 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14168 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12144 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10580 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 20424 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 19780 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 14260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11040 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 10672 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 17848 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 18676 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 15088 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 19228 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 16836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 17388 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 20608 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 20148 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10212 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 19872 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 16008 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 17664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 20884 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1649977179
transform -1 0 20516 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 8556 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8740 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 20884 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 20516 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 10672 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 15640 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16468 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 9384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 10488 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 9108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 19412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 16928 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 17296 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 16284 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9568 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 9936 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 10488 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 9108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 10304 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 10488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5152 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 4968 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 5060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 4692 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 10028 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 10396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 3772 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7360 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 7820 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 7912 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8280 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 4508 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4508 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 5060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6164 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 10120 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 10856 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 4692 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5704 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 5060 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 6164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 6072 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 6900 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6072 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 4600 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 8648 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7084 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 7544 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 7912 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1649977179
transform -1 0 20240 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 11684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 7544 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 8464 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 8096 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14352 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12972 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15088 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 15732 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 18860 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 18952 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 21252 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 20424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 20056 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 20056 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17572 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 14168 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 14628 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 19780 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 18676 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13248 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14720 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 11684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13524 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12512 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 12144 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13156 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12328 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 14076 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 21252 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 19964 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 5520 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 4968 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 18676 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16100 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 11408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 13616 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 16192 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16100 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 5612 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 4876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 14720 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7728 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 19320 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 19688 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 19780 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 20424 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15456 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 14904 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 19320 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 12052 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_93
timestamp 1649977179
transform 1 0 9660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_98 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_102
timestamp 1649977179
transform 1 0 10488 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_106
timestamp 1649977179
transform 1 0 10856 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1649977179
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1649977179
transform 1 0 11776 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1649977179
transform 1 0 12328 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_128
timestamp 1649977179
transform 1 0 12880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1649977179
transform 1 0 13432 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1649977179
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_145 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149
timestamp 1649977179
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_154
timestamp 1649977179
transform 1 0 15272 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_158
timestamp 1649977179
transform 1 0 15640 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_162
timestamp 1649977179
transform 1 0 16008 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1649977179
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_172
timestamp 1649977179
transform 1 0 16928 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_176
timestamp 1649977179
transform 1 0 17296 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_180
timestamp 1649977179
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_184
timestamp 1649977179
transform 1 0 18032 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_189
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_199
timestamp 1649977179
transform 1 0 19412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_203
timestamp 1649977179
transform 1 0 19780 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_207
timestamp 1649977179
transform 1 0 20148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_211
timestamp 1649977179
transform 1 0 20516 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_215
timestamp 1649977179
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_89
timestamp 1649977179
transform 1 0 9292 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_92
timestamp 1649977179
transform 1 0 9568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_96
timestamp 1649977179
transform 1 0 9936 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_100
timestamp 1649977179
transform 1 0 10304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_104
timestamp 1649977179
transform 1 0 10672 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1649977179
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_115
timestamp 1649977179
transform 1 0 11684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_123
timestamp 1649977179
transform 1 0 12420 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_133
timestamp 1649977179
transform 1 0 13340 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_147
timestamp 1649977179
transform 1 0 14628 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_158
timestamp 1649977179
transform 1 0 15640 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1649977179
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_173
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_177
timestamp 1649977179
transform 1 0 17388 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_182
timestamp 1649977179
transform 1 0 17848 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1649977179
transform 1 0 18400 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_194
timestamp 1649977179
transform 1 0 18952 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_200
timestamp 1649977179
transform 1 0 19504 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_206
timestamp 1649977179
transform 1 0 20056 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_210
timestamp 1649977179
transform 1 0 20424 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_218
timestamp 1649977179
transform 1 0 21160 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_222
timestamp 1649977179
transform 1 0 21528 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1649977179
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1649977179
transform 1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_105
timestamp 1649977179
transform 1 0 10764 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_113
timestamp 1649977179
transform 1 0 11500 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_125
timestamp 1649977179
transform 1 0 12604 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_130
timestamp 1649977179
transform 1 0 13064 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1649977179
transform 1 0 14996 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_162
timestamp 1649977179
transform 1 0 16008 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_173
timestamp 1649977179
transform 1 0 17020 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_181
timestamp 1649977179
transform 1 0 17756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_193
timestamp 1649977179
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_199
timestamp 1649977179
transform 1 0 19412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_203
timestamp 1649977179
transform 1 0 19780 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_207
timestamp 1649977179
transform 1 0 20148 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_211
timestamp 1649977179
transform 1 0 20516 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1649977179
transform 1 0 20884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_85
timestamp 1649977179
transform 1 0 8924 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_91
timestamp 1649977179
transform 1 0 9476 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_94
timestamp 1649977179
transform 1 0 9752 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_98
timestamp 1649977179
transform 1 0 10120 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_102
timestamp 1649977179
transform 1 0 10488 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1649977179
transform 1 0 10856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1649977179
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_122
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_126
timestamp 1649977179
transform 1 0 12696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_138
timestamp 1649977179
transform 1 0 13800 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_143
timestamp 1649977179
transform 1 0 14260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_147
timestamp 1649977179
transform 1 0 14628 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_153
timestamp 1649977179
transform 1 0 15180 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1649977179
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_171
timestamp 1649977179
transform 1 0 16836 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_175
timestamp 1649977179
transform 1 0 17204 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_182
timestamp 1649977179
transform 1 0 17848 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_192
timestamp 1649977179
transform 1 0 18768 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_196
timestamp 1649977179
transform 1 0 19136 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1649977179
transform 1 0 19504 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_204
timestamp 1649977179
transform 1 0 19872 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_208
timestamp 1649977179
transform 1 0 20240 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_212
timestamp 1649977179
transform 1 0 20608 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_216
timestamp 1649977179
transform 1 0 20976 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1649977179
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1649977179
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_89
timestamp 1649977179
transform 1 0 9292 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_100
timestamp 1649977179
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_112
timestamp 1649977179
transform 1 0 11408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_123
timestamp 1649977179
transform 1 0 12420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_134
timestamp 1649977179
transform 1 0 13432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1649977179
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_150
timestamp 1649977179
transform 1 0 14904 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_161
timestamp 1649977179
transform 1 0 15916 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_169
timestamp 1649977179
transform 1 0 16652 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_173
timestamp 1649977179
transform 1 0 17020 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_180
timestamp 1649977179
transform 1 0 17664 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_191
timestamp 1649977179
transform 1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_200
timestamp 1649977179
transform 1 0 19504 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_204
timestamp 1649977179
transform 1 0 19872 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_208
timestamp 1649977179
transform 1 0 20240 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1649977179
transform 1 0 20608 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_217
timestamp 1649977179
transform 1 0 21068 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_77
timestamp 1649977179
transform 1 0 8188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_85
timestamp 1649977179
transform 1 0 8924 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_89
timestamp 1649977179
transform 1 0 9292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_100
timestamp 1649977179
transform 1 0 10304 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_104
timestamp 1649977179
transform 1 0 10672 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_124
timestamp 1649977179
transform 1 0 12512 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_129
timestamp 1649977179
transform 1 0 12972 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_140
timestamp 1649977179
transform 1 0 13984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_144
timestamp 1649977179
transform 1 0 14352 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_155
timestamp 1649977179
transform 1 0 15364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1649977179
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_173
timestamp 1649977179
transform 1 0 17020 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_185
timestamp 1649977179
transform 1 0 18124 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_196
timestamp 1649977179
transform 1 0 19136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_207
timestamp 1649977179
transform 1 0 20148 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_218
timestamp 1649977179
transform 1 0 21160 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1649977179
transform 1 0 21528 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_87
timestamp 1649977179
transform 1 0 9108 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_98
timestamp 1649977179
transform 1 0 10120 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_102
timestamp 1649977179
transform 1 0 10488 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_113
timestamp 1649977179
transform 1 0 11500 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_126
timestamp 1649977179
transform 1 0 12696 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_137
timestamp 1649977179
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_143
timestamp 1649977179
transform 1 0 14260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_148
timestamp 1649977179
transform 1 0 14720 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_159
timestamp 1649977179
transform 1 0 15732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_170
timestamp 1649977179
transform 1 0 16744 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_181
timestamp 1649977179
transform 1 0 17756 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_220
timestamp 1649977179
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_92
timestamp 1649977179
transform 1 0 9568 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_103
timestamp 1649977179
transform 1 0 10580 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_107
timestamp 1649977179
transform 1 0 10948 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1649977179
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_136
timestamp 1649977179
transform 1 0 13616 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_140
timestamp 1649977179
transform 1 0 13984 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_150
timestamp 1649977179
transform 1 0 14904 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_165
timestamp 1649977179
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_178
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_189
timestamp 1649977179
transform 1 0 18492 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_197
timestamp 1649977179
transform 1 0 19228 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_201
timestamp 1649977179
transform 1 0 19596 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_208
timestamp 1649977179
transform 1 0 20240 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1649977179
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_56
timestamp 1649977179
transform 1 0 6256 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_68
timestamp 1649977179
transform 1 0 7360 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1649977179
transform 1 0 9384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_95
timestamp 1649977179
transform 1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_99
timestamp 1649977179
transform 1 0 10212 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1649977179
transform 1 0 10488 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_106
timestamp 1649977179
transform 1 0 10856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_110
timestamp 1649977179
transform 1 0 11224 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_114
timestamp 1649977179
transform 1 0 11592 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_125
timestamp 1649977179
transform 1 0 12604 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_130
timestamp 1649977179
transform 1 0 13064 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_134
timestamp 1649977179
transform 1 0 13432 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1649977179
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_150
timestamp 1649977179
transform 1 0 14904 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_155
timestamp 1649977179
transform 1 0 15364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_166
timestamp 1649977179
transform 1 0 16376 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_181
timestamp 1649977179
transform 1 0 17756 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_191
timestamp 1649977179
transform 1 0 18676 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_199
timestamp 1649977179
transform 1 0 19412 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_203
timestamp 1649977179
transform 1 0 19780 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_208
timestamp 1649977179
transform 1 0 20240 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1649977179
transform 1 0 20608 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_218
timestamp 1649977179
transform 1 0 21160 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_222
timestamp 1649977179
transform 1 0 21528 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_35
timestamp 1649977179
transform 1 0 4324 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_50
timestamp 1649977179
transform 1 0 5704 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1649977179
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_66
timestamp 1649977179
transform 1 0 7176 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_78
timestamp 1649977179
transform 1 0 8280 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_95
timestamp 1649977179
transform 1 0 9844 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_99
timestamp 1649977179
transform 1 0 10212 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_103
timestamp 1649977179
transform 1 0 10580 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_107
timestamp 1649977179
transform 1 0 10948 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1649977179
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_122
timestamp 1649977179
transform 1 0 12328 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_126
timestamp 1649977179
transform 1 0 12696 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_130
timestamp 1649977179
transform 1 0 13064 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_140
timestamp 1649977179
transform 1 0 13984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_151
timestamp 1649977179
transform 1 0 14996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_162
timestamp 1649977179
transform 1 0 16008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1649977179
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_178
timestamp 1649977179
transform 1 0 17480 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_191
timestamp 1649977179
transform 1 0 18676 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_199
timestamp 1649977179
transform 1 0 19412 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_203
timestamp 1649977179
transform 1 0 19780 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_211
timestamp 1649977179
transform 1 0 20516 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_219
timestamp 1649977179
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_37
timestamp 1649977179
transform 1 0 4508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_52
timestamp 1649977179
transform 1 0 5888 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_63
timestamp 1649977179
transform 1 0 6900 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_75
timestamp 1649977179
transform 1 0 8004 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_94
timestamp 1649977179
transform 1 0 9752 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_100
timestamp 1649977179
transform 1 0 10304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_104
timestamp 1649977179
transform 1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_115
timestamp 1649977179
transform 1 0 11684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_119
timestamp 1649977179
transform 1 0 12052 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_129
timestamp 1649977179
transform 1 0 12972 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_150
timestamp 1649977179
transform 1 0 14904 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_155
timestamp 1649977179
transform 1 0 15364 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_161
timestamp 1649977179
transform 1 0 15916 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_166
timestamp 1649977179
transform 1 0 16376 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_182
timestamp 1649977179
transform 1 0 17848 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1649977179
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_203
timestamp 1649977179
transform 1 0 19780 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_213
timestamp 1649977179
transform 1 0 20700 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_219
timestamp 1649977179
transform 1 0 21252 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_45
timestamp 1649977179
transform 1 0 5244 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_49
timestamp 1649977179
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_60
timestamp 1649977179
transform 1 0 6624 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_72
timestamp 1649977179
transform 1 0 7728 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_76
timestamp 1649977179
transform 1 0 8096 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_80
timestamp 1649977179
transform 1 0 8464 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_86
timestamp 1649977179
transform 1 0 9016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_96
timestamp 1649977179
transform 1 0 9936 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1649977179
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_116
timestamp 1649977179
transform 1 0 11776 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1649977179
transform 1 0 12144 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_124
timestamp 1649977179
transform 1 0 12512 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_128
timestamp 1649977179
transform 1 0 12880 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_131
timestamp 1649977179
transform 1 0 13156 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_142
timestamp 1649977179
transform 1 0 14168 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_146
timestamp 1649977179
transform 1 0 14536 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_150
timestamp 1649977179
transform 1 0 14904 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_154
timestamp 1649977179
transform 1 0 15272 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_158
timestamp 1649977179
transform 1 0 15640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1649977179
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_178
timestamp 1649977179
transform 1 0 17480 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_182
timestamp 1649977179
transform 1 0 17848 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_194
timestamp 1649977179
transform 1 0 18952 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_198
timestamp 1649977179
transform 1 0 19320 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_204
timestamp 1649977179
transform 1 0 19872 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_210
timestamp 1649977179
transform 1 0 20424 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1649977179
transform 1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_57
timestamp 1649977179
transform 1 0 6348 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_61
timestamp 1649977179
transform 1 0 6716 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_71
timestamp 1649977179
transform 1 0 7636 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_75
timestamp 1649977179
transform 1 0 8004 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_79
timestamp 1649977179
transform 1 0 8372 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_102
timestamp 1649977179
transform 1 0 10488 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_106
timestamp 1649977179
transform 1 0 10856 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_112
timestamp 1649977179
transform 1 0 11408 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_115
timestamp 1649977179
transform 1 0 11684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_126
timestamp 1649977179
transform 1 0 12696 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1649977179
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_143
timestamp 1649977179
transform 1 0 14260 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_147
timestamp 1649977179
transform 1 0 14628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_150
timestamp 1649977179
transform 1 0 14904 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_154
timestamp 1649977179
transform 1 0 15272 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_158
timestamp 1649977179
transform 1 0 15640 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_168
timestamp 1649977179
transform 1 0 16560 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp 1649977179
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_203
timestamp 1649977179
transform 1 0 19780 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_207
timestamp 1649977179
transform 1 0 20148 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1649977179
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_35
timestamp 1649977179
transform 1 0 4324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_43
timestamp 1649977179
transform 1 0 5060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1649977179
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_66
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_77
timestamp 1649977179
transform 1 0 8188 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_88
timestamp 1649977179
transform 1 0 9200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_92
timestamp 1649977179
transform 1 0 9568 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_104
timestamp 1649977179
transform 1 0 10672 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1649977179
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115
timestamp 1649977179
transform 1 0 11684 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1649977179
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_129
timestamp 1649977179
transform 1 0 12972 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_140
timestamp 1649977179
transform 1 0 13984 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_152
timestamp 1649977179
transform 1 0 15088 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_163
timestamp 1649977179
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_178
timestamp 1649977179
transform 1 0 17480 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_189
timestamp 1649977179
transform 1 0 18492 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_197
timestamp 1649977179
transform 1 0 19228 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_216
timestamp 1649977179
transform 1 0 20976 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_45
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_55
timestamp 1649977179
transform 1 0 6164 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_66
timestamp 1649977179
transform 1 0 7176 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_70
timestamp 1649977179
transform 1 0 7544 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_74
timestamp 1649977179
transform 1 0 7912 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_78
timestamp 1649977179
transform 1 0 8280 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_96
timestamp 1649977179
transform 1 0 9936 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_107
timestamp 1649977179
transform 1 0 10948 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_112
timestamp 1649977179
transform 1 0 11408 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_117
timestamp 1649977179
transform 1 0 11868 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_131
timestamp 1649977179
transform 1 0 13156 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp 1649977179
transform 1 0 13524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_144
timestamp 1649977179
transform 1 0 14352 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_148
timestamp 1649977179
transform 1 0 14720 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_161
timestamp 1649977179
transform 1 0 15916 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1649977179
transform 1 0 16744 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_178
timestamp 1649977179
transform 1 0 17480 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1649977179
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_206
timestamp 1649977179
transform 1 0 20056 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_214
timestamp 1649977179
transform 1 0 20792 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_220
timestamp 1649977179
transform 1 0 21344 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1649977179
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_66
timestamp 1649977179
transform 1 0 7176 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_71
timestamp 1649977179
transform 1 0 7636 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_76
timestamp 1649977179
transform 1 0 8096 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_87
timestamp 1649977179
transform 1 0 9108 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_99
timestamp 1649977179
transform 1 0 10212 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1649977179
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_115
timestamp 1649977179
transform 1 0 11684 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1649977179
transform 1 0 12144 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_131
timestamp 1649977179
transform 1 0 13156 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_142
timestamp 1649977179
transform 1 0 14168 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_153
timestamp 1649977179
transform 1 0 15180 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_157
timestamp 1649977179
transform 1 0 15548 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1649977179
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_175
timestamp 1649977179
transform 1 0 17204 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_192
timestamp 1649977179
transform 1 0 18768 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_196
timestamp 1649977179
transform 1 0 19136 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_206
timestamp 1649977179
transform 1 0 20056 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1649977179
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_49
timestamp 1649977179
transform 1 0 5612 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_60
timestamp 1649977179
transform 1 0 6624 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_71
timestamp 1649977179
transform 1 0 7636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_88
timestamp 1649977179
transform 1 0 9200 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_107
timestamp 1649977179
transform 1 0 10948 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_111
timestamp 1649977179
transform 1 0 11316 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_132
timestamp 1649977179
transform 1 0 13248 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1649977179
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1649977179
transform 1 0 14996 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_162
timestamp 1649977179
transform 1 0 16008 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_166
timestamp 1649977179
transform 1 0 16376 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1649977179
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1649977179
transform 1 0 17112 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_185
timestamp 1649977179
transform 1 0 18124 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1649977179
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_206
timestamp 1649977179
transform 1 0 20056 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_217
timestamp 1649977179
transform 1 0 21068 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_43
timestamp 1649977179
transform 1 0 5060 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1649977179
transform 1 0 6808 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_73
timestamp 1649977179
transform 1 0 7820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_85
timestamp 1649977179
transform 1 0 8924 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_104
timestamp 1649977179
transform 1 0 10672 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1649977179
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_115
timestamp 1649977179
transform 1 0 11684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_119
timestamp 1649977179
transform 1 0 12052 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_123
timestamp 1649977179
transform 1 0 12420 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_127
timestamp 1649977179
transform 1 0 12788 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_141
timestamp 1649977179
transform 1 0 14076 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1649977179
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_159
timestamp 1649977179
transform 1 0 15732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_163
timestamp 1649977179
transform 1 0 16100 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_173
timestamp 1649977179
transform 1 0 17020 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_199
timestamp 1649977179
transform 1 0 19412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_203
timestamp 1649977179
transform 1 0 19780 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1649977179
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_44
timestamp 1649977179
transform 1 0 5152 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_48
timestamp 1649977179
transform 1 0 5520 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_64
timestamp 1649977179
transform 1 0 6992 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_103
timestamp 1649977179
transform 1 0 10580 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_107
timestamp 1649977179
transform 1 0 10948 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_126
timestamp 1649977179
transform 1 0 12696 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_130
timestamp 1649977179
transform 1 0 13064 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_134
timestamp 1649977179
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_157
timestamp 1649977179
transform 1 0 15548 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_175
timestamp 1649977179
transform 1 0 17204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1649977179
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_203
timestamp 1649977179
transform 1 0 19780 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_74
timestamp 1649977179
transform 1 0 7912 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_92
timestamp 1649977179
transform 1 0 9568 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1649977179
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_115
timestamp 1649977179
transform 1 0 11684 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1649977179
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_122
timestamp 1649977179
transform 1 0 12328 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_126
timestamp 1649977179
transform 1 0 12696 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_144
timestamp 1649977179
transform 1 0 14352 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_162
timestamp 1649977179
transform 1 0 16008 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1649977179
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_185
timestamp 1649977179
transform 1 0 18124 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_203
timestamp 1649977179
transform 1 0 19780 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1649977179
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_51
timestamp 1649977179
transform 1 0 5796 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_55
timestamp 1649977179
transform 1 0 6164 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_63
timestamp 1649977179
transform 1 0 6900 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1649977179
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1649977179
transform 1 0 10488 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_120
timestamp 1649977179
transform 1 0 12144 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1649977179
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_157
timestamp 1649977179
transform 1 0 15548 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_161
timestamp 1649977179
transform 1 0 15916 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_180
timestamp 1649977179
transform 1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_188
timestamp 1649977179
transform 1 0 18400 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1649977179
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_213
timestamp 1649977179
transform 1 0 20700 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_219
timestamp 1649977179
transform 1 0 21252 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_29
timestamp 1649977179
transform 1 0 3772 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_37
timestamp 1649977179
transform 1 0 4508 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_42
timestamp 1649977179
transform 1 0 4968 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_46
timestamp 1649977179
transform 1 0 5336 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_74
timestamp 1649977179
transform 1 0 7912 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_78
timestamp 1649977179
transform 1 0 8280 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_82
timestamp 1649977179
transform 1 0 8648 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_86
timestamp 1649977179
transform 1 0 9016 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_104
timestamp 1649977179
transform 1 0 10672 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1649977179
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_141
timestamp 1649977179
transform 1 0 14076 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_159
timestamp 1649977179
transform 1 0 15732 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_163
timestamp 1649977179
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_185
timestamp 1649977179
transform 1 0 18124 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_203
timestamp 1649977179
transform 1 0 19780 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1649977179
transform 1 0 21436 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_23
timestamp 1649977179
transform 1 0 3220 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1649977179
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_40
timestamp 1649977179
transform 1 0 4784 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_51
timestamp 1649977179
transform 1 0 5796 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_62
timestamp 1649977179
transform 1 0 6808 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_72
timestamp 1649977179
transform 1 0 7728 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_104
timestamp 1649977179
transform 1 0 10672 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_108
timestamp 1649977179
transform 1 0 11040 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_120
timestamp 1649977179
transform 1 0 12144 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_132
timestamp 1649977179
transform 1 0 13248 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1649977179
transform 1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_147
timestamp 1649977179
transform 1 0 14628 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_183
timestamp 1649977179
transform 1 0 17940 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_187
timestamp 1649977179
transform 1 0 18308 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_191
timestamp 1649977179
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_199
timestamp 1649977179
transform 1 0 19412 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_203
timestamp 1649977179
transform 1 0 19780 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_33
timestamp 1649977179
transform 1 0 4140 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_43
timestamp 1649977179
transform 1 0 5060 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_60
timestamp 1649977179
transform 1 0 6624 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_71
timestamp 1649977179
transform 1 0 7636 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_83
timestamp 1649977179
transform 1 0 8740 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_91
timestamp 1649977179
transform 1 0 9476 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1649977179
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_115
timestamp 1649977179
transform 1 0 11684 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_127
timestamp 1649977179
transform 1 0 12788 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_139
timestamp 1649977179
transform 1 0 13892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_144
timestamp 1649977179
transform 1 0 14352 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_148
timestamp 1649977179
transform 1 0 14720 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1649977179
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_171
timestamp 1649977179
transform 1 0 16836 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_175
timestamp 1649977179
transform 1 0 17204 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_185
timestamp 1649977179
transform 1 0 18124 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_189
timestamp 1649977179
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_192
timestamp 1649977179
transform 1 0 18768 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_196
timestamp 1649977179
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_200
timestamp 1649977179
transform 1 0 19504 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_218
timestamp 1649977179
transform 1 0 21160 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_222
timestamp 1649977179
transform 1 0 21528 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_37
timestamp 1649977179
transform 1 0 4508 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_40
timestamp 1649977179
transform 1 0 4784 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_57
timestamp 1649977179
transform 1 0 6348 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_68
timestamp 1649977179
transform 1 0 7360 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_72
timestamp 1649977179
transform 1 0 7728 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_76
timestamp 1649977179
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_88
timestamp 1649977179
transform 1 0 9200 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_110
timestamp 1649977179
transform 1 0 11224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_114
timestamp 1649977179
transform 1 0 11592 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_134
timestamp 1649977179
transform 1 0 13432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1649977179
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_158
timestamp 1649977179
transform 1 0 15640 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_176
timestamp 1649977179
transform 1 0 17296 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_180
timestamp 1649977179
transform 1 0 17664 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_184
timestamp 1649977179
transform 1 0 18032 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_187
timestamp 1649977179
transform 1 0 18308 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_191
timestamp 1649977179
transform 1 0 18676 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1649977179
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_199
timestamp 1649977179
transform 1 0 19412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_203
timestamp 1649977179
transform 1 0 19780 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_38
timestamp 1649977179
transform 1 0 4600 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_49
timestamp 1649977179
transform 1 0 5612 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1649977179
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_66
timestamp 1649977179
transform 1 0 7176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_86
timestamp 1649977179
transform 1 0 9016 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_104
timestamp 1649977179
transform 1 0 10672 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1649977179
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_133
timestamp 1649977179
transform 1 0 13340 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_151
timestamp 1649977179
transform 1 0 14996 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_155
timestamp 1649977179
transform 1 0 15364 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_160
timestamp 1649977179
transform 1 0 15824 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_185
timestamp 1649977179
transform 1 0 18124 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_211
timestamp 1649977179
transform 1 0 20516 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1649977179
transform 1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_40
timestamp 1649977179
transform 1 0 4784 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_52
timestamp 1649977179
transform 1 0 5888 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_61
timestamp 1649977179
transform 1 0 6716 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1649977179
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_102
timestamp 1649977179
transform 1 0 10488 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_120
timestamp 1649977179
transform 1 0 12144 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_124
timestamp 1649977179
transform 1 0 12512 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_128
timestamp 1649977179
transform 1 0 12880 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_131
timestamp 1649977179
transform 1 0 13156 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_135
timestamp 1649977179
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_157
timestamp 1649977179
transform 1 0 15548 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_175
timestamp 1649977179
transform 1 0 17204 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1649977179
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_213
timestamp 1649977179
transform 1 0 20700 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1649977179
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_35
timestamp 1649977179
transform 1 0 4324 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_43
timestamp 1649977179
transform 1 0 5060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1649977179
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_80
timestamp 1649977179
transform 1 0 8464 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_84
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_102
timestamp 1649977179
transform 1 0 10488 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_106
timestamp 1649977179
transform 1 0 10856 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1649977179
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_115
timestamp 1649977179
transform 1 0 11684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_119
timestamp 1649977179
transform 1 0 12052 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_123
timestamp 1649977179
transform 1 0 12420 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_127
timestamp 1649977179
transform 1 0 12788 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_131
timestamp 1649977179
transform 1 0 13156 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_135
timestamp 1649977179
transform 1 0 13524 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_153
timestamp 1649977179
transform 1 0 15180 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_159
timestamp 1649977179
transform 1 0 15732 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_163
timestamp 1649977179
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_171
timestamp 1649977179
transform 1 0 16836 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_177
timestamp 1649977179
transform 1 0 17388 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_185
timestamp 1649977179
transform 1 0 18124 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_191
timestamp 1649977179
transform 1 0 18676 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_209
timestamp 1649977179
transform 1 0 20332 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_218
timestamp 1649977179
transform 1 0 21160 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_222
timestamp 1649977179
transform 1 0 21528 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_61
timestamp 1649977179
transform 1 0 6716 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_70
timestamp 1649977179
transform 1 0 7544 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1649977179
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_87
timestamp 1649977179
transform 1 0 9108 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_93
timestamp 1649977179
transform 1 0 9660 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_110
timestamp 1649977179
transform 1 0 11224 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_114
timestamp 1649977179
transform 1 0 11592 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_132
timestamp 1649977179
transform 1 0 13248 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1649977179
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_143
timestamp 1649977179
transform 1 0 14260 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_147
timestamp 1649977179
transform 1 0 14628 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_150
timestamp 1649977179
transform 1 0 14904 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_168
timestamp 1649977179
transform 1 0 16560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_172
timestamp 1649977179
transform 1 0 16928 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_190
timestamp 1649977179
transform 1 0 18584 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1649977179
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_203
timestamp 1649977179
transform 1 0 19780 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_63
timestamp 1649977179
transform 1 0 6900 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_67
timestamp 1649977179
transform 1 0 7268 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp 1649977179
transform 1 0 8280 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_82
timestamp 1649977179
transform 1 0 8648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_102
timestamp 1649977179
transform 1 0 10488 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_106
timestamp 1649977179
transform 1 0 10856 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1649977179
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1649977179
transform 1 0 11960 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_122
timestamp 1649977179
transform 1 0 12328 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_140
timestamp 1649977179
transform 1 0 13984 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_159
timestamp 1649977179
transform 1 0 15732 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1649977179
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_185
timestamp 1649977179
transform 1 0 18124 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_203
timestamp 1649977179
transform 1 0 19780 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1649977179
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_49
timestamp 1649977179
transform 1 0 5612 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_52
timestamp 1649977179
transform 1 0 5888 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_56
timestamp 1649977179
transform 1 0 6256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_64
timestamp 1649977179
transform 1 0 6992 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1649977179
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_101
timestamp 1649977179
transform 1 0 10396 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_105
timestamp 1649977179
transform 1 0 10764 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_128
timestamp 1649977179
transform 1 0 12880 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_132
timestamp 1649977179
transform 1 0 13248 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_143
timestamp 1649977179
transform 1 0 14260 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_161
timestamp 1649977179
transform 1 0 15916 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_169
timestamp 1649977179
transform 1 0 16652 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_187
timestamp 1649977179
transform 1 0 18308 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1649977179
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_213
timestamp 1649977179
transform 1 0 20700 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_43
timestamp 1649977179
transform 1 0 5060 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1649977179
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_66
timestamp 1649977179
transform 1 0 7176 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_74
timestamp 1649977179
transform 1 0 7912 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_92
timestamp 1649977179
transform 1 0 9568 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1649977179
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_115
timestamp 1649977179
transform 1 0 11684 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_119
timestamp 1649977179
transform 1 0 12052 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_123
timestamp 1649977179
transform 1 0 12420 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_127
timestamp 1649977179
transform 1 0 12788 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_145
timestamp 1649977179
transform 1 0 14444 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1649977179
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_171
timestamp 1649977179
transform 1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_189
timestamp 1649977179
transform 1 0 18492 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_207
timestamp 1649977179
transform 1 0 20148 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_35
timestamp 1649977179
transform 1 0 4324 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_40
timestamp 1649977179
transform 1 0 4784 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_44
timestamp 1649977179
transform 1 0 5152 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_48
timestamp 1649977179
transform 1 0 5520 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_51
timestamp 1649977179
transform 1 0 5796 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_57
timestamp 1649977179
transform 1 0 6348 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_70
timestamp 1649977179
transform 1 0 7544 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_76
timestamp 1649977179
transform 1 0 8096 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1649977179
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_104
timestamp 1649977179
transform 1 0 10672 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_122
timestamp 1649977179
transform 1 0 12328 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_126
timestamp 1649977179
transform 1 0 12696 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_130
timestamp 1649977179
transform 1 0 13064 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1649977179
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_157
timestamp 1649977179
transform 1 0 15548 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_167
timestamp 1649977179
transform 1 0 16468 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_175
timestamp 1649977179
transform 1 0 17204 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_181
timestamp 1649977179
transform 1 0 17756 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_187
timestamp 1649977179
transform 1 0 18308 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_193
timestamp 1649977179
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1649977179
transform 1 0 19780 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_29
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_41
timestamp 1649977179
transform 1 0 4876 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_47
timestamp 1649977179
transform 1 0 5428 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_50
timestamp 1649977179
transform 1 0 5704 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1649977179
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_64
timestamp 1649977179
transform 1 0 6992 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_70
timestamp 1649977179
transform 1 0 7544 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_76
timestamp 1649977179
transform 1 0 8096 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_82
timestamp 1649977179
transform 1 0 8648 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_94
timestamp 1649977179
transform 1 0 9752 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_103
timestamp 1649977179
transform 1 0 10580 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_107
timestamp 1649977179
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_115
timestamp 1649977179
transform 1 0 11684 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_119
timestamp 1649977179
transform 1 0 12052 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_122
timestamp 1649977179
transform 1 0 12328 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_126
timestamp 1649977179
transform 1 0 12696 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_130
timestamp 1649977179
transform 1 0 13064 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_134
timestamp 1649977179
transform 1 0 13432 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_138
timestamp 1649977179
transform 1 0 13800 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_145
timestamp 1649977179
transform 1 0 14444 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_155
timestamp 1649977179
transform 1 0 15364 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_162
timestamp 1649977179
transform 1 0 16008 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1649977179
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_173
timestamp 1649977179
transform 1 0 17020 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_187
timestamp 1649977179
transform 1 0 18308 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_201
timestamp 1649977179
transform 1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1649977179
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _033_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1649977179
transform -1 0 16744 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1649977179
transform -1 0 6256 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1649977179
transform -1 0 17848 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1649977179
transform -1 0 17020 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1649977179
transform -1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1649977179
transform -1 0 16376 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1649977179
transform 1 0 10856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1649977179
transform -1 0 12144 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1649977179
transform 1 0 11592 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1649977179
transform 1 0 5336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1649977179
transform -1 0 5980 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1649977179
transform 1 0 21160 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1649977179
transform -1 0 13340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1649977179
transform 1 0 18676 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1649977179
transform 1 0 7360 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1649977179
transform -1 0 6808 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1649977179
transform -1 0 13064 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1649977179
transform -1 0 21068 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1649977179
transform -1 0 15364 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1649977179
transform -1 0 14720 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1649977179
transform -1 0 12972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1649977179
transform -1 0 15180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1649977179
transform 1 0 9568 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1649977179
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1649977179
transform 1 0 6440 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1649977179
transform 1 0 10212 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _066_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20792 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1649977179
transform 1 0 18032 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1649977179
transform 1 0 18584 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1649977179
transform 1 0 20976 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1649977179
transform 1 0 20884 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1649977179
transform -1 0 17756 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1649977179
transform -1 0 19964 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1649977179
transform 1 0 20884 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1649977179
transform 1 0 20148 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1649977179
transform 1 0 19504 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1649977179
transform 1 0 19412 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1649977179
transform 1 0 20700 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1649977179
transform 1 0 20056 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1649977179
transform 1 0 20148 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1649977179
transform 1 0 20884 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1649977179
transform -1 0 18952 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1649977179
transform -1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1649977179
transform -1 0 18124 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1649977179
transform 1 0 18492 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1649977179
transform 1 0 19412 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1649977179
transform -1 0 11224 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1649977179
transform 1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1649977179
transform 1 0 12512 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1649977179
transform 1 0 13064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1649977179
transform 1 0 12696 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1649977179
transform 1 0 13248 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1649977179
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1649977179
transform -1 0 17020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1649977179
transform -1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1649977179
transform 1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1649977179
transform 1 0 18124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1649977179
transform 1 0 17480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1649977179
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1649977179
transform 1 0 20792 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1649977179
transform 1 0 18584 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1649977179
transform 1 0 7728 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1649977179
transform 1 0 6624 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1649977179
transform 1 0 7728 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1649977179
transform 1 0 8280 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1649977179
transform -1 0 6348 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1649977179
transform 1 0 7176 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1649977179
transform 1 0 4416 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1649977179
transform 1 0 8280 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1649977179
transform -1 0 18308 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1649977179
transform 1 0 15640 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1649977179
transform -1 0 18860 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1649977179
transform 1 0 13248 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1649977179
transform 1 0 14996 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1649977179
transform -1 0 18308 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1649977179
transform 1 0 18308 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7176 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9108 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10672 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6440 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16192 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20700 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15732 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16376 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15640 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13524 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 15824 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19780 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21436 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17940 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18308 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13800 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10948 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7176 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13432 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10488 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10672 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9752 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13340 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 9016 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8648 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9016 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11224 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10488 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10856 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13984 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 9568 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9752 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12880 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10396 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8648 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9752 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14444 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10672 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16100 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14260 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18492 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19688 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17020 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20700 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20148 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17204 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14812 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16468 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18860 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10672 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8096 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9752 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11224 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14352 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9016 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12144 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11776 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15088 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16008 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10672 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15180 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10672 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14444 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18584 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15732 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 20332 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18952 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18308 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 18308 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12328 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17664 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12880 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11684 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12788 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 10672 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12604 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform -1 0 16100 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16560 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 15548 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15180 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12236 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13800 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14904 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 15088 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12972 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12604 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11592 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1649977179
transform -1 0 15364 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1649977179
transform -1 0 16192 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 16192 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14168 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13340 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19320 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1649977179
transform -1 0 18952 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17848 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1649977179
transform 1 0 17296 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 17296 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16376 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 20608 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform -1 0 20332 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1649977179
transform 1 0 20516 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 20332 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18768 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16928 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15916 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15916 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 17112 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10580 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9476 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9476 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9568 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 10120 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10580 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20700 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5796 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform -1 0 6072 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1649977179
transform -1 0 9844 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1649977179
transform -1 0 7176 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7636 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10120 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10028 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15824 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4784 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6348 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6900 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1649977179
transform -1 0 5704 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5980 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 6900 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 7176 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6072 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1649977179
transform -1 0 6164 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9108 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_3_
timestamp 1649977179
transform -1 0 5888 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7176 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8188 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 16928 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5796 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5244 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5796 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 17204 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4784 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4600 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5060 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18400 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7176 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_1_
timestamp 1649977179
transform -1 0 6348 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l3_in_0_
timestamp 1649977179
transform -1 0 7360 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20240 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9200 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_1_
timestamp 1649977179
transform -1 0 9936 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10672 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 16836 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14168 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1649977179
transform -1 0 14904 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14996 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16560 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_1_
timestamp 1649977179
transform -1 0 17480 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18676 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_1_
timestamp 1649977179
transform -1 0 18676 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18032 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16376 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20240 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_1_
timestamp 1649977179
transform 1 0 20240 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1649977179
transform -1 0 20056 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20148 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14076 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13984 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19688 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17388 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13984 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14168 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19504 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11868 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10948 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20608 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12972 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13156 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20884 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10856 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10212 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15916 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12420 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17296 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6164 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 6624 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 7728 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7912 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1649977179
transform -1 0 12604 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11868 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6992 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7084 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12236 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1649977179
transform -1 0 6072 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12880 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7636 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6808 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6992 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14996 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8280 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14352 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8096 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7636 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7544 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18124 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17664 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18492 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1649977179
transform 1 0 20148 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1649977179
transform 1 0 17664 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17204 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15088 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14260 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12144 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10580 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20608 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20424 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1649977179
transform -1 0 18768 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 1142 592
<< labels >>
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 386 0 442 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_1_
port 2 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 ccff_head
port 3 nsew signal input
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal3 s 22200 4904 23000 5024 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 5 nsew signal input
flabel metal3 s 22200 8984 23000 9104 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 6 nsew signal input
flabel metal3 s 22200 9392 23000 9512 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 7 nsew signal input
flabel metal3 s 22200 9800 23000 9920 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 8 nsew signal input
flabel metal3 s 22200 10208 23000 10328 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 9 nsew signal input
flabel metal3 s 22200 10616 23000 10736 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 10 nsew signal input
flabel metal3 s 22200 11024 23000 11144 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 11 nsew signal input
flabel metal3 s 22200 11432 23000 11552 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 12 nsew signal input
flabel metal3 s 22200 11840 23000 11960 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 13 nsew signal input
flabel metal3 s 22200 12248 23000 12368 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 14 nsew signal input
flabel metal3 s 22200 12656 23000 12776 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 15 nsew signal input
flabel metal3 s 22200 5312 23000 5432 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 16 nsew signal input
flabel metal3 s 22200 5720 23000 5840 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 17 nsew signal input
flabel metal3 s 22200 6128 23000 6248 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 18 nsew signal input
flabel metal3 s 22200 6536 23000 6656 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 19 nsew signal input
flabel metal3 s 22200 6944 23000 7064 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 20 nsew signal input
flabel metal3 s 22200 7352 23000 7472 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 21 nsew signal input
flabel metal3 s 22200 7760 23000 7880 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 22 nsew signal input
flabel metal3 s 22200 8168 23000 8288 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 23 nsew signal input
flabel metal3 s 22200 8576 23000 8696 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 24 nsew signal input
flabel metal3 s 22200 13064 23000 13184 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 25 nsew signal tristate
flabel metal3 s 22200 17144 23000 17264 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 26 nsew signal tristate
flabel metal3 s 22200 17552 23000 17672 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 27 nsew signal tristate
flabel metal3 s 22200 17960 23000 18080 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 28 nsew signal tristate
flabel metal3 s 22200 18368 23000 18488 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 29 nsew signal tristate
flabel metal3 s 22200 18776 23000 18896 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 30 nsew signal tristate
flabel metal3 s 22200 19184 23000 19304 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 31 nsew signal tristate
flabel metal3 s 22200 19592 23000 19712 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 32 nsew signal tristate
flabel metal3 s 22200 20000 23000 20120 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 33 nsew signal tristate
flabel metal3 s 22200 20408 23000 20528 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 34 nsew signal tristate
flabel metal3 s 22200 20816 23000 20936 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 35 nsew signal tristate
flabel metal3 s 22200 13472 23000 13592 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 36 nsew signal tristate
flabel metal3 s 22200 13880 23000 14000 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 37 nsew signal tristate
flabel metal3 s 22200 14288 23000 14408 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 38 nsew signal tristate
flabel metal3 s 22200 14696 23000 14816 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 39 nsew signal tristate
flabel metal3 s 22200 15104 23000 15224 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 40 nsew signal tristate
flabel metal3 s 22200 15512 23000 15632 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 41 nsew signal tristate
flabel metal3 s 22200 15920 23000 16040 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 42 nsew signal tristate
flabel metal3 s 22200 16328 23000 16448 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 43 nsew signal tristate
flabel metal3 s 22200 16736 23000 16856 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 44 nsew signal tristate
flabel metal2 s 938 0 994 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 45 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 46 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 47 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 48 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 49 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 50 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 51 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 52 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 53 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 54 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 55 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 56 nsew signal input
flabel metal2 s 2042 0 2098 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 57 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 58 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 59 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 60 nsew signal input
flabel metal2 s 4250 0 4306 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 61 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 62 nsew signal input
flabel metal2 s 5354 0 5410 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 63 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 64 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 65 nsew signal tristate
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 66 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 67 nsew signal tristate
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 68 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 69 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 70 nsew signal tristate
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 71 nsew signal tristate
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 72 nsew signal tristate
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 73 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 74 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 75 nsew signal tristate
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 76 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 77 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 78 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 79 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 80 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 81 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 82 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 83 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 84 nsew signal tristate
flabel metal2 s 938 22200 994 23000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 85 nsew signal input
flabel metal2 s 6458 22200 6514 23000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 86 nsew signal input
flabel metal2 s 7010 22200 7066 23000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 87 nsew signal input
flabel metal2 s 7562 22200 7618 23000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 88 nsew signal input
flabel metal2 s 8114 22200 8170 23000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 89 nsew signal input
flabel metal2 s 8666 22200 8722 23000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 90 nsew signal input
flabel metal2 s 9218 22200 9274 23000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 91 nsew signal input
flabel metal2 s 9770 22200 9826 23000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 92 nsew signal input
flabel metal2 s 10322 22200 10378 23000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 93 nsew signal input
flabel metal2 s 10874 22200 10930 23000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 94 nsew signal input
flabel metal2 s 11426 22200 11482 23000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 95 nsew signal input
flabel metal2 s 1490 22200 1546 23000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 96 nsew signal input
flabel metal2 s 2042 22200 2098 23000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 97 nsew signal input
flabel metal2 s 2594 22200 2650 23000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 98 nsew signal input
flabel metal2 s 3146 22200 3202 23000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 99 nsew signal input
flabel metal2 s 3698 22200 3754 23000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 100 nsew signal input
flabel metal2 s 4250 22200 4306 23000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 101 nsew signal input
flabel metal2 s 4802 22200 4858 23000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 102 nsew signal input
flabel metal2 s 5354 22200 5410 23000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 103 nsew signal input
flabel metal2 s 5906 22200 5962 23000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 104 nsew signal input
flabel metal2 s 11978 22200 12034 23000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 105 nsew signal tristate
flabel metal2 s 17498 22200 17554 23000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 106 nsew signal tristate
flabel metal2 s 18050 22200 18106 23000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 107 nsew signal tristate
flabel metal2 s 18602 22200 18658 23000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 108 nsew signal tristate
flabel metal2 s 19154 22200 19210 23000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 109 nsew signal tristate
flabel metal2 s 19706 22200 19762 23000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 110 nsew signal tristate
flabel metal2 s 20258 22200 20314 23000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 111 nsew signal tristate
flabel metal2 s 20810 22200 20866 23000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 112 nsew signal tristate
flabel metal2 s 21362 22200 21418 23000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 113 nsew signal tristate
flabel metal2 s 21914 22200 21970 23000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 114 nsew signal tristate
flabel metal2 s 22466 22200 22522 23000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 115 nsew signal tristate
flabel metal2 s 12530 22200 12586 23000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 116 nsew signal tristate
flabel metal2 s 13082 22200 13138 23000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 117 nsew signal tristate
flabel metal2 s 13634 22200 13690 23000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 118 nsew signal tristate
flabel metal2 s 14186 22200 14242 23000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 119 nsew signal tristate
flabel metal2 s 14738 22200 14794 23000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 120 nsew signal tristate
flabel metal2 s 15290 22200 15346 23000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 121 nsew signal tristate
flabel metal2 s 15842 22200 15898 23000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 122 nsew signal tristate
flabel metal2 s 16394 22200 16450 23000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 123 nsew signal tristate
flabel metal2 s 16946 22200 17002 23000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 124 nsew signal tristate
flabel metal3 s 22200 21224 23000 21344 0 FreeSans 480 0 0 0 prog_clk_0_E_in
port 125 nsew signal input
flabel metal3 s 22200 1640 23000 1760 0 FreeSans 480 0 0 0 right_bottom_grid_pin_34_
port 126 nsew signal input
flabel metal3 s 22200 2048 23000 2168 0 FreeSans 480 0 0 0 right_bottom_grid_pin_35_
port 127 nsew signal input
flabel metal3 s 22200 2456 23000 2576 0 FreeSans 480 0 0 0 right_bottom_grid_pin_36_
port 128 nsew signal input
flabel metal3 s 22200 2864 23000 2984 0 FreeSans 480 0 0 0 right_bottom_grid_pin_37_
port 129 nsew signal input
flabel metal3 s 22200 3272 23000 3392 0 FreeSans 480 0 0 0 right_bottom_grid_pin_38_
port 130 nsew signal input
flabel metal3 s 22200 3680 23000 3800 0 FreeSans 480 0 0 0 right_bottom_grid_pin_39_
port 131 nsew signal input
flabel metal3 s 22200 4088 23000 4208 0 FreeSans 480 0 0 0 right_bottom_grid_pin_40_
port 132 nsew signal input
flabel metal3 s 22200 4496 23000 4616 0 FreeSans 480 0 0 0 right_bottom_grid_pin_41_
port 133 nsew signal input
flabel metal2 s 386 22200 442 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_1_
port 134 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
