magic
tech sky130A
magscale 1 2
timestamp 1679321272
<< viali >>
rect 22569 54281 22603 54315
rect 23213 54281 23247 54315
rect 26157 54281 26191 54315
rect 27813 54281 27847 54315
rect 28917 54281 28951 54315
rect 32781 54281 32815 54315
rect 3249 54213 3283 54247
rect 8401 54213 8435 54247
rect 10701 54213 10735 54247
rect 13553 54213 13587 54247
rect 15853 54213 15887 54247
rect 18705 54213 18739 54247
rect 28825 54213 28859 54247
rect 29837 54213 29871 54247
rect 32689 54213 32723 54247
rect 33425 54213 33459 54247
rect 34161 54213 34195 54247
rect 34989 54213 35023 54247
rect 37841 54213 37875 54247
rect 42625 54213 42659 54247
rect 2237 54145 2271 54179
rect 4813 54145 4847 54179
rect 7389 54145 7423 54179
rect 9965 54145 9999 54179
rect 12541 54145 12575 54179
rect 14933 54145 14967 54179
rect 17693 54145 17727 54179
rect 20085 54145 20119 54179
rect 22753 54145 22787 54179
rect 23397 54145 23431 54179
rect 24041 54145 24075 54179
rect 25053 54145 25087 54179
rect 25697 54145 25731 54179
rect 26341 54145 26375 54179
rect 27353 54145 27387 54179
rect 27997 54145 28031 54179
rect 30665 54145 30699 54179
rect 31309 54145 31343 54179
rect 35817 54145 35851 54179
rect 36461 54145 36495 54179
rect 38669 54145 38703 54179
rect 40049 54145 40083 54179
rect 45201 54145 45235 54179
rect 45937 54145 45971 54179
rect 46673 54145 46707 54179
rect 47777 54145 47811 54179
rect 48513 54145 48547 54179
rect 5457 54077 5491 54111
rect 20545 54077 20579 54111
rect 33609 54077 33643 54111
rect 38945 54077 38979 54111
rect 40325 54077 40359 54111
rect 23857 54009 23891 54043
rect 25513 54009 25547 54043
rect 35633 54009 35667 54043
rect 36277 54009 36311 54043
rect 24869 53941 24903 53975
rect 27169 53941 27203 53975
rect 29929 53941 29963 53975
rect 30481 53941 30515 53975
rect 31125 53941 31159 53975
rect 34253 53941 34287 53975
rect 35081 53941 35115 53975
rect 37933 53941 37967 53975
rect 43913 53941 43947 53975
rect 45385 53941 45419 53975
rect 46121 53941 46155 53975
rect 46857 53941 46891 53975
rect 47961 53941 47995 53975
rect 48697 53941 48731 53975
rect 36461 53737 36495 53771
rect 31309 53669 31343 53703
rect 37105 53669 37139 53703
rect 2881 53601 2915 53635
rect 6101 53601 6135 53635
rect 7849 53601 7883 53635
rect 11253 53601 11287 53635
rect 13369 53601 13403 53635
rect 16405 53601 16439 53635
rect 18337 53601 18371 53635
rect 21465 53601 21499 53635
rect 2237 53533 2271 53567
rect 5457 53533 5491 53567
rect 7389 53533 7423 53567
rect 10701 53533 10735 53567
rect 12357 53533 12391 53567
rect 15669 53533 15703 53567
rect 17693 53533 17727 53567
rect 21005 53533 21039 53567
rect 23029 53533 23063 53567
rect 28273 53533 28307 53567
rect 31493 53533 31527 53567
rect 32137 53533 32171 53567
rect 36645 53533 36679 53567
rect 37289 53533 37323 53567
rect 38485 53533 38519 53567
rect 40509 53533 40543 53567
rect 44189 53533 44223 53567
rect 46765 53533 46799 53567
rect 48237 53533 48271 53567
rect 48697 53533 48731 53567
rect 38669 53465 38703 53499
rect 22845 53397 22879 53431
rect 28089 53397 28123 53431
rect 31953 53397 31987 53431
rect 40325 53397 40359 53431
rect 44373 53397 44407 53431
rect 46949 53397 46983 53431
rect 48053 53397 48087 53431
rect 48881 53397 48915 53431
rect 2513 53057 2547 53091
rect 4721 53057 4755 53091
rect 7665 53057 7699 53091
rect 9965 53057 9999 53091
rect 12633 53057 12667 53091
rect 15117 53057 15151 53091
rect 17785 53057 17819 53091
rect 19901 53057 19935 53091
rect 22201 53057 22235 53091
rect 49065 53057 49099 53091
rect 2789 52989 2823 53023
rect 5089 52989 5123 53023
rect 7941 52989 7975 53023
rect 10241 52989 10275 53023
rect 13093 52989 13127 53023
rect 15393 52989 15427 53023
rect 18245 52989 18279 53023
rect 20177 52989 20211 53023
rect 22017 52853 22051 52887
rect 49249 52853 49283 52887
rect 21005 52649 21039 52683
rect 49249 52581 49283 52615
rect 2145 52513 2179 52547
rect 4721 52513 4755 52547
rect 7297 52513 7331 52547
rect 9873 52513 9907 52547
rect 12449 52513 12483 52547
rect 15025 52513 15059 52547
rect 17601 52513 17635 52547
rect 1869 52445 1903 52479
rect 4261 52445 4295 52479
rect 7021 52445 7055 52479
rect 9597 52445 9631 52479
rect 11989 52445 12023 52479
rect 14565 52445 14599 52479
rect 17141 52445 17175 52479
rect 21189 52445 21223 52479
rect 49065 52445 49099 52479
rect 7757 52105 7791 52139
rect 9689 52105 9723 52139
rect 10333 52105 10367 52139
rect 15577 52105 15611 52139
rect 17601 52105 17635 52139
rect 18889 52105 18923 52139
rect 8677 52037 8711 52071
rect 7941 51969 7975 52003
rect 8493 51969 8527 52003
rect 9873 51969 9907 52003
rect 10517 51969 10551 52003
rect 15761 51969 15795 52003
rect 17785 51969 17819 52003
rect 19073 51969 19107 52003
rect 17049 51765 17083 51799
rect 7665 51561 7699 51595
rect 9229 51561 9263 51595
rect 10885 51561 10919 51595
rect 13553 51561 13587 51595
rect 8585 51493 8619 51527
rect 17601 51493 17635 51527
rect 2053 51425 2087 51459
rect 14933 51425 14967 51459
rect 18613 51425 18647 51459
rect 19993 51425 20027 51459
rect 20085 51425 20119 51459
rect 1777 51357 1811 51391
rect 7849 51357 7883 51391
rect 9413 51357 9447 51391
rect 11069 51357 11103 51391
rect 13737 51357 13771 51391
rect 15853 51357 15887 51391
rect 18521 51357 18555 51391
rect 8401 51289 8435 51323
rect 16129 51289 16163 51323
rect 18061 51221 18095 51255
rect 18429 51221 18463 51255
rect 19533 51221 19567 51255
rect 19901 51221 19935 51255
rect 8401 51017 8435 51051
rect 9045 51017 9079 51051
rect 12173 51017 12207 51051
rect 12817 51017 12851 51051
rect 21005 51017 21039 51051
rect 23489 51017 23523 51051
rect 13553 50949 13587 50983
rect 17325 50949 17359 50983
rect 20269 50949 20303 50983
rect 1777 50881 1811 50915
rect 8585 50881 8619 50915
rect 9229 50881 9263 50915
rect 12357 50881 12391 50915
rect 13001 50881 13035 50915
rect 17049 50881 17083 50915
rect 20177 50881 20211 50915
rect 21189 50881 21223 50915
rect 23397 50881 23431 50915
rect 2053 50813 2087 50847
rect 14565 50813 14599 50847
rect 14841 50813 14875 50847
rect 20361 50813 20395 50847
rect 23581 50813 23615 50847
rect 37565 50813 37599 50847
rect 37841 50813 37875 50847
rect 13645 50677 13679 50711
rect 16313 50677 16347 50711
rect 18797 50677 18831 50711
rect 19809 50677 19843 50711
rect 23029 50677 23063 50711
rect 39313 50677 39347 50711
rect 11713 50473 11747 50507
rect 13553 50473 13587 50507
rect 16129 50473 16163 50507
rect 23305 50473 23339 50507
rect 17417 50337 17451 50371
rect 20269 50337 20303 50371
rect 23857 50337 23891 50371
rect 11897 50269 11931 50303
rect 14381 50269 14415 50303
rect 17141 50269 17175 50303
rect 20913 50269 20947 50303
rect 23765 50269 23799 50303
rect 49065 50269 49099 50303
rect 13461 50201 13495 50235
rect 14657 50201 14691 50235
rect 20085 50201 20119 50235
rect 21189 50201 21223 50235
rect 18889 50133 18923 50167
rect 19717 50133 19751 50167
rect 20177 50133 20211 50167
rect 22661 50133 22695 50167
rect 23673 50133 23707 50167
rect 49249 50133 49283 50167
rect 15853 49929 15887 49963
rect 17141 49929 17175 49963
rect 17601 49929 17635 49963
rect 23397 49929 23431 49963
rect 23857 49929 23891 49963
rect 12173 49861 12207 49895
rect 12725 49861 12759 49895
rect 13645 49861 13679 49895
rect 19073 49861 19107 49895
rect 22017 49861 22051 49895
rect 22845 49861 22879 49895
rect 1777 49793 1811 49827
rect 11989 49793 12023 49827
rect 13461 49793 13495 49827
rect 17509 49793 17543 49827
rect 18337 49793 18371 49827
rect 19717 49793 19751 49827
rect 23765 49793 23799 49827
rect 2053 49725 2087 49759
rect 12909 49725 12943 49759
rect 14105 49725 14139 49759
rect 17693 49725 17727 49759
rect 21465 49725 21499 49759
rect 23949 49725 23983 49759
rect 14368 49589 14402 49623
rect 19980 49589 20014 49623
rect 13001 49385 13035 49419
rect 11805 49317 11839 49351
rect 12541 49317 12575 49351
rect 15945 49317 15979 49351
rect 19717 49317 19751 49351
rect 2053 49249 2087 49283
rect 13645 49249 13679 49283
rect 15301 49249 15335 49283
rect 16405 49249 16439 49283
rect 16497 49249 16531 49283
rect 17141 49249 17175 49283
rect 17417 49249 17451 49283
rect 18889 49249 18923 49283
rect 20821 49249 20855 49283
rect 20913 49249 20947 49283
rect 21557 49249 21591 49283
rect 21833 49249 21867 49283
rect 24961 49249 24995 49283
rect 26065 49249 26099 49283
rect 1777 49181 1811 49215
rect 13369 49181 13403 49215
rect 15117 49181 15151 49215
rect 15209 49181 15243 49215
rect 24869 49181 24903 49215
rect 11621 49113 11655 49147
rect 12357 49113 12391 49147
rect 13461 49113 13495 49147
rect 19533 49113 19567 49147
rect 20729 49113 20763 49147
rect 24777 49113 24811 49147
rect 14749 49045 14783 49079
rect 16313 49045 16347 49079
rect 20361 49045 20395 49079
rect 23305 49045 23339 49079
rect 24409 49045 24443 49079
rect 25513 49045 25547 49079
rect 25881 49045 25915 49079
rect 25973 49045 26007 49079
rect 9597 48841 9631 48875
rect 15945 48841 15979 48875
rect 17785 48841 17819 48875
rect 20177 48841 20211 48875
rect 23765 48841 23799 48875
rect 25053 48841 25087 48875
rect 25973 48841 26007 48875
rect 16037 48773 16071 48807
rect 9781 48705 9815 48739
rect 13001 48705 13035 48739
rect 17693 48705 17727 48739
rect 19257 48705 19291 48739
rect 20361 48705 20395 48739
rect 22017 48705 22051 48739
rect 25881 48705 25915 48739
rect 13277 48637 13311 48671
rect 16221 48637 16255 48671
rect 17877 48637 17911 48671
rect 19349 48637 19383 48671
rect 19533 48637 19567 48671
rect 22293 48637 22327 48671
rect 26065 48637 26099 48671
rect 12541 48501 12575 48535
rect 14749 48501 14783 48535
rect 15577 48501 15611 48535
rect 17325 48501 17359 48535
rect 18889 48501 18923 48535
rect 21005 48501 21039 48535
rect 25513 48501 25547 48535
rect 16405 48297 16439 48331
rect 24041 48229 24075 48263
rect 2053 48161 2087 48195
rect 13645 48161 13679 48195
rect 14657 48161 14691 48195
rect 17141 48161 17175 48195
rect 17417 48161 17451 48195
rect 20269 48161 20303 48195
rect 22569 48161 22603 48195
rect 26341 48161 26375 48195
rect 1777 48093 1811 48127
rect 12541 48093 12575 48127
rect 13369 48093 13403 48127
rect 13461 48093 13495 48127
rect 19993 48093 20027 48127
rect 21281 48093 21315 48127
rect 22293 48093 22327 48127
rect 26157 48093 26191 48127
rect 14933 48025 14967 48059
rect 20085 48025 20119 48059
rect 25329 48025 25363 48059
rect 26249 48025 26283 48059
rect 48973 48025 49007 48059
rect 13001 47957 13035 47991
rect 18889 47957 18923 47991
rect 19625 47957 19659 47991
rect 21097 47957 21131 47991
rect 25789 47957 25823 47991
rect 49065 47957 49099 47991
rect 9689 47753 9723 47787
rect 10333 47753 10367 47787
rect 11713 47753 11747 47787
rect 15945 47753 15979 47787
rect 16037 47753 16071 47787
rect 25329 47753 25363 47787
rect 26249 47753 26283 47787
rect 1777 47617 1811 47651
rect 9873 47617 9907 47651
rect 10517 47617 10551 47651
rect 11161 47617 11195 47651
rect 11897 47617 11931 47651
rect 19717 47617 19751 47651
rect 23029 47617 23063 47651
rect 26157 47617 26191 47651
rect 2053 47549 2087 47583
rect 13369 47549 13403 47583
rect 13645 47549 13679 47583
rect 15117 47549 15151 47583
rect 16221 47549 16255 47583
rect 17417 47549 17451 47583
rect 17693 47549 17727 47583
rect 19993 47549 20027 47583
rect 22201 47549 22235 47583
rect 23305 47549 23339 47583
rect 24777 47549 24811 47583
rect 26341 47549 26375 47583
rect 10977 47481 11011 47515
rect 15577 47413 15611 47447
rect 19165 47413 19199 47447
rect 21465 47413 21499 47447
rect 25789 47413 25823 47447
rect 11161 47209 11195 47243
rect 18889 47209 18923 47243
rect 21373 47209 21407 47243
rect 24041 47209 24075 47243
rect 11805 47141 11839 47175
rect 13001 47141 13035 47175
rect 16037 47141 16071 47175
rect 12265 47073 12299 47107
rect 12357 47073 12391 47107
rect 13645 47073 13679 47107
rect 14289 47073 14323 47107
rect 17141 47073 17175 47107
rect 17417 47073 17451 47107
rect 22569 47073 22603 47107
rect 11345 47005 11379 47039
rect 13461 47005 13495 47039
rect 16681 47005 16715 47039
rect 19625 47005 19659 47039
rect 22293 47005 22327 47039
rect 12173 46937 12207 46971
rect 14565 46937 14599 46971
rect 19901 46937 19935 46971
rect 13369 46869 13403 46903
rect 4261 46665 4295 46699
rect 5181 46665 5215 46699
rect 10977 46665 11011 46699
rect 13829 46665 13863 46699
rect 16313 46665 16347 46699
rect 21465 46665 21499 46699
rect 24133 46665 24167 46699
rect 1777 46529 1811 46563
rect 4169 46529 4203 46563
rect 5089 46529 5123 46563
rect 11161 46529 11195 46563
rect 12909 46529 12943 46563
rect 13737 46529 13771 46563
rect 17509 46529 17543 46563
rect 25513 46529 25547 46563
rect 25605 46529 25639 46563
rect 2053 46461 2087 46495
rect 14013 46461 14047 46495
rect 14565 46461 14599 46495
rect 14841 46461 14875 46495
rect 17785 46461 17819 46495
rect 19717 46461 19751 46495
rect 19993 46461 20027 46495
rect 22385 46461 22419 46495
rect 22661 46461 22695 46495
rect 24685 46461 24719 46495
rect 25697 46461 25731 46495
rect 13369 46393 13403 46427
rect 17049 46325 17083 46359
rect 19257 46325 19291 46359
rect 25145 46325 25179 46359
rect 4169 46121 4203 46155
rect 8033 46121 8067 46155
rect 11253 46121 11287 46155
rect 13737 46121 13771 46155
rect 16313 46121 16347 46155
rect 18889 46121 18923 46155
rect 20348 46121 20382 46155
rect 2053 45985 2087 46019
rect 14841 45985 14875 46019
rect 17141 45985 17175 46019
rect 17417 45985 17451 46019
rect 20085 45985 20119 46019
rect 22569 45985 22603 46019
rect 1777 45917 1811 45951
rect 8217 45917 8251 45951
rect 11437 45917 11471 45951
rect 14565 45917 14599 45951
rect 19625 45917 19659 45951
rect 22293 45917 22327 45951
rect 47961 45917 47995 45951
rect 49157 45917 49191 45951
rect 4077 45849 4111 45883
rect 21833 45781 21867 45815
rect 24041 45781 24075 45815
rect 19349 45577 19383 45611
rect 2697 45509 2731 45543
rect 3893 45509 3927 45543
rect 4629 45509 4663 45543
rect 15945 45509 15979 45543
rect 20085 45509 20119 45543
rect 2513 45441 2547 45475
rect 3709 45441 3743 45475
rect 4445 45441 4479 45475
rect 8125 45441 8159 45475
rect 9229 45441 9263 45475
rect 11897 45441 11931 45475
rect 12725 45441 12759 45475
rect 14473 45441 14507 45475
rect 15117 45441 15151 45475
rect 17417 45441 17451 45475
rect 19257 45441 19291 45475
rect 22201 45441 22235 45475
rect 16037 45373 16071 45407
rect 16129 45373 16163 45407
rect 18245 45373 18279 45407
rect 19441 45373 19475 45407
rect 20913 45373 20947 45407
rect 22845 45373 22879 45407
rect 23121 45373 23155 45407
rect 7941 45305 7975 45339
rect 9045 45305 9079 45339
rect 12541 45305 12575 45339
rect 15577 45305 15611 45339
rect 11713 45237 11747 45271
rect 14289 45237 14323 45271
rect 14933 45237 14967 45271
rect 18889 45237 18923 45271
rect 24593 45237 24627 45271
rect 4169 45033 4203 45067
rect 4905 45033 4939 45067
rect 9137 45033 9171 45067
rect 11069 45033 11103 45067
rect 15117 45033 15151 45067
rect 13093 44965 13127 44999
rect 16957 44965 16991 44999
rect 18153 44965 18187 44999
rect 2053 44897 2087 44931
rect 16405 44897 16439 44931
rect 17601 44897 17635 44931
rect 18613 44897 18647 44931
rect 18797 44897 18831 44931
rect 19441 44897 19475 44931
rect 22293 44897 22327 44931
rect 27445 44897 27479 44931
rect 1777 44829 1811 44863
rect 9321 44829 9355 44863
rect 9965 44829 9999 44863
rect 10609 44829 10643 44863
rect 11253 44829 11287 44863
rect 11897 44829 11931 44863
rect 12541 44829 12575 44863
rect 13277 44829 13311 44863
rect 14473 44829 14507 44863
rect 15301 44829 15335 44863
rect 17325 44829 17359 44863
rect 17417 44829 17451 44863
rect 18521 44829 18555 44863
rect 22109 44829 22143 44863
rect 26341 44829 26375 44863
rect 27169 44829 27203 44863
rect 4077 44761 4111 44795
rect 4813 44761 4847 44795
rect 19717 44761 19751 44795
rect 9781 44693 9815 44727
rect 10425 44693 10459 44727
rect 14289 44693 14323 44727
rect 15761 44693 15795 44727
rect 16129 44693 16163 44727
rect 16221 44693 16255 44727
rect 21189 44693 21223 44727
rect 21649 44693 21683 44727
rect 22017 44693 22051 44727
rect 26801 44693 26835 44727
rect 27261 44693 27295 44727
rect 27997 44693 28031 44727
rect 4537 44489 4571 44523
rect 8585 44489 8619 44523
rect 12817 44489 12851 44523
rect 17509 44489 17543 44523
rect 20269 44489 20303 44523
rect 3801 44421 3835 44455
rect 4445 44421 4479 44455
rect 9321 44421 9355 44455
rect 20729 44421 20763 44455
rect 1777 44353 1811 44387
rect 3617 44353 3651 44387
rect 8769 44353 8803 44387
rect 13001 44353 13035 44387
rect 17049 44353 17083 44387
rect 17693 44353 17727 44387
rect 18337 44353 18371 44387
rect 19165 44353 19199 44387
rect 19257 44353 19291 44387
rect 20637 44353 20671 44387
rect 22201 44353 22235 44387
rect 24869 44353 24903 44387
rect 2053 44285 2087 44319
rect 19441 44285 19475 44319
rect 20821 44285 20855 44319
rect 25145 44285 25179 44319
rect 18797 44217 18831 44251
rect 9413 44149 9447 44183
rect 11069 44149 11103 44183
rect 12357 44149 12391 44183
rect 18153 44149 18187 44183
rect 26617 44149 26651 44183
rect 5089 43945 5123 43979
rect 10701 43945 10735 43979
rect 11253 43945 11287 43979
rect 13461 43945 13495 43979
rect 17693 43945 17727 43979
rect 18889 43945 18923 43979
rect 20913 43945 20947 43979
rect 24041 43945 24075 43979
rect 26801 43945 26835 43979
rect 14289 43877 14323 43911
rect 11805 43809 11839 43843
rect 20085 43809 20119 43843
rect 22569 43809 22603 43843
rect 25237 43809 25271 43843
rect 27813 43809 27847 43843
rect 4997 43741 5031 43775
rect 10609 43741 10643 43775
rect 11621 43741 11655 43775
rect 13001 43741 13035 43775
rect 13645 43741 13679 43775
rect 14473 43741 14507 43775
rect 15485 43741 15519 43775
rect 17877 43741 17911 43775
rect 19901 43741 19935 43775
rect 21833 43741 21867 43775
rect 22293 43741 22327 43775
rect 25053 43741 25087 43775
rect 27721 43741 27755 43775
rect 11713 43673 11747 43707
rect 15761 43673 15795 43707
rect 24961 43673 24995 43707
rect 27629 43673 27663 43707
rect 28457 43673 28491 43707
rect 12817 43605 12851 43639
rect 17233 43605 17267 43639
rect 19533 43605 19567 43639
rect 19993 43605 20027 43639
rect 24593 43605 24627 43639
rect 27261 43605 27295 43639
rect 9781 43401 9815 43435
rect 10425 43401 10459 43435
rect 10793 43401 10827 43435
rect 11713 43401 11747 43435
rect 12081 43401 12115 43435
rect 13461 43401 13495 43435
rect 14841 43401 14875 43435
rect 15301 43401 15335 43435
rect 19901 43401 19935 43435
rect 20729 43401 20763 43435
rect 22385 43401 22419 43435
rect 22477 43401 22511 43435
rect 10885 43333 10919 43367
rect 14197 43333 14231 43367
rect 21189 43333 21223 43367
rect 1777 43265 1811 43299
rect 9137 43265 9171 43299
rect 9965 43265 9999 43299
rect 13645 43265 13679 43299
rect 15209 43265 15243 43299
rect 16313 43265 16347 43299
rect 17049 43265 17083 43299
rect 17693 43265 17727 43299
rect 21097 43265 21131 43299
rect 2053 43197 2087 43231
rect 10977 43197 11011 43231
rect 12173 43197 12207 43231
rect 12265 43197 12299 43231
rect 15393 43197 15427 43231
rect 18153 43197 18187 43231
rect 18429 43197 18463 43231
rect 21373 43197 21407 43231
rect 22661 43197 22695 43231
rect 14381 43129 14415 43163
rect 9229 43061 9263 43095
rect 16129 43061 16163 43095
rect 17509 43061 17543 43095
rect 22017 43061 22051 43095
rect 7008 42857 7042 42891
rect 11529 42857 11563 42891
rect 12246 42857 12280 42891
rect 16110 42857 16144 42891
rect 21084 42857 21118 42891
rect 2053 42721 2087 42755
rect 4813 42721 4847 42755
rect 6745 42721 6779 42755
rect 11989 42721 12023 42755
rect 15025 42721 15059 42755
rect 17601 42721 17635 42755
rect 19993 42721 20027 42755
rect 20821 42721 20855 42755
rect 1593 42653 1627 42687
rect 4629 42653 4663 42687
rect 9321 42653 9355 42687
rect 9781 42653 9815 42687
rect 15853 42653 15887 42687
rect 10057 42585 10091 42619
rect 14749 42585 14783 42619
rect 18153 42585 18187 42619
rect 18705 42585 18739 42619
rect 8493 42517 8527 42551
rect 9137 42517 9171 42551
rect 13737 42517 13771 42551
rect 14381 42517 14415 42551
rect 14841 42517 14875 42551
rect 18797 42517 18831 42551
rect 19441 42517 19475 42551
rect 19809 42517 19843 42551
rect 19901 42517 19935 42551
rect 22569 42517 22603 42551
rect 4997 42313 5031 42347
rect 13461 42313 13495 42347
rect 16313 42313 16347 42347
rect 17233 42313 17267 42347
rect 20729 42313 20763 42347
rect 21097 42313 21131 42347
rect 24133 42313 24167 42347
rect 4905 42177 4939 42211
rect 8769 42177 8803 42211
rect 11161 42177 11195 42211
rect 11713 42177 11747 42211
rect 17417 42177 17451 42211
rect 18061 42177 18095 42211
rect 19349 42177 19383 42211
rect 19901 42177 19935 42211
rect 19993 42177 20027 42211
rect 22385 42177 22419 42211
rect 9045 42109 9079 42143
rect 12449 42109 12483 42143
rect 13553 42109 13587 42143
rect 13645 42109 13679 42143
rect 14565 42109 14599 42143
rect 14841 42109 14875 42143
rect 18981 42109 19015 42143
rect 20085 42109 20119 42143
rect 21189 42109 21223 42143
rect 21281 42109 21315 42143
rect 22661 42109 22695 42143
rect 10517 42041 10551 42075
rect 13093 42041 13127 42075
rect 19533 42041 19567 42075
rect 10977 41973 11011 42007
rect 17877 41973 17911 42007
rect 22293 41973 22327 42007
rect 4813 41769 4847 41803
rect 13001 41769 13035 41803
rect 18061 41769 18095 41803
rect 21005 41769 21039 41803
rect 9965 41701 9999 41735
rect 14289 41701 14323 41735
rect 17233 41701 17267 41735
rect 17785 41701 17819 41735
rect 2053 41633 2087 41667
rect 10425 41633 10459 41667
rect 10701 41633 10735 41667
rect 13461 41633 13495 41667
rect 13645 41633 13679 41667
rect 14749 41633 14783 41667
rect 14933 41633 14967 41667
rect 15761 41633 15795 41667
rect 18521 41633 18555 41667
rect 18705 41633 18739 41667
rect 21557 41633 21591 41667
rect 22569 41633 22603 41667
rect 23857 41633 23891 41667
rect 1777 41565 1811 41599
rect 4721 41565 4755 41599
rect 8585 41565 8619 41599
rect 9781 41565 9815 41599
rect 15485 41565 15519 41599
rect 17969 41565 18003 41599
rect 18429 41565 18463 41599
rect 19073 41565 19107 41599
rect 20177 41565 20211 41599
rect 20729 41565 20763 41599
rect 20913 41565 20947 41599
rect 23673 41565 23707 41599
rect 6469 41497 6503 41531
rect 14657 41497 14691 41531
rect 21465 41497 21499 41531
rect 22385 41497 22419 41531
rect 6561 41429 6595 41463
rect 12173 41429 12207 41463
rect 13369 41429 13403 41463
rect 21373 41429 21407 41463
rect 22017 41429 22051 41463
rect 22477 41429 22511 41463
rect 23305 41429 23339 41463
rect 23765 41429 23799 41463
rect 16313 41225 16347 41259
rect 16865 41225 16899 41259
rect 19257 41225 19291 41259
rect 19625 41225 19659 41259
rect 20545 41225 20579 41259
rect 24501 41225 24535 41259
rect 24869 41225 24903 41259
rect 24961 41225 24995 41259
rect 6745 41157 6779 41191
rect 23489 41157 23523 41191
rect 23581 41157 23615 41191
rect 1777 41089 1811 41123
rect 8033 41089 8067 41123
rect 9413 41089 9447 41123
rect 12357 41089 12391 41123
rect 14565 41089 14599 41123
rect 17233 41089 17267 41123
rect 19717 41089 19751 41123
rect 22661 41089 22695 41123
rect 2053 41021 2087 41055
rect 8769 41021 8803 41055
rect 9689 41021 9723 41055
rect 12633 41021 12667 41055
rect 14105 41021 14139 41055
rect 14841 41021 14875 41055
rect 17325 41021 17359 41055
rect 17509 41021 17543 41055
rect 19901 41021 19935 41055
rect 23673 41021 23707 41055
rect 25053 41021 25087 41055
rect 6929 40953 6963 40987
rect 11161 40885 11195 40919
rect 11897 40885 11931 40919
rect 18705 40885 18739 40919
rect 23121 40885 23155 40919
rect 24409 40885 24443 40919
rect 7849 40681 7883 40715
rect 9137 40681 9171 40715
rect 11989 40681 12023 40715
rect 13001 40681 13035 40715
rect 17128 40681 17162 40715
rect 7389 40613 7423 40647
rect 8401 40545 8435 40579
rect 9689 40545 9723 40579
rect 13553 40545 13587 40579
rect 14289 40545 14323 40579
rect 16865 40545 16899 40579
rect 20913 40545 20947 40579
rect 21833 40545 21867 40579
rect 25145 40545 25179 40579
rect 8217 40477 8251 40511
rect 10241 40477 10275 40511
rect 13369 40477 13403 40511
rect 13461 40477 13495 40511
rect 21557 40477 21591 40511
rect 23857 40477 23891 40511
rect 25053 40477 25087 40511
rect 9597 40409 9631 40443
rect 10517 40409 10551 40443
rect 14565 40409 14599 40443
rect 18889 40409 18923 40443
rect 20729 40409 20763 40443
rect 24961 40409 24995 40443
rect 8309 40341 8343 40375
rect 9505 40341 9539 40375
rect 12541 40341 12575 40375
rect 16037 40341 16071 40375
rect 19809 40341 19843 40375
rect 20361 40341 20395 40375
rect 20821 40341 20855 40375
rect 23305 40341 23339 40375
rect 24593 40341 24627 40375
rect 25881 40341 25915 40375
rect 10241 40137 10275 40171
rect 7849 40069 7883 40103
rect 10977 40069 11011 40103
rect 15485 40069 15519 40103
rect 17601 40069 17635 40103
rect 19993 40069 20027 40103
rect 22017 40069 22051 40103
rect 1777 40001 1811 40035
rect 8493 40001 8527 40035
rect 11713 40001 11747 40035
rect 19717 40001 19751 40035
rect 24685 40001 24719 40035
rect 2053 39933 2087 39967
rect 7297 39933 7331 39967
rect 8769 39933 8803 39967
rect 11989 39933 12023 39967
rect 13461 39933 13495 39967
rect 15577 39933 15611 39967
rect 15669 39933 15703 39967
rect 18337 39933 18371 39967
rect 22753 39933 22787 39967
rect 24777 39933 24811 39967
rect 24869 39933 24903 39967
rect 14657 39865 14691 39899
rect 7941 39797 7975 39831
rect 11069 39797 11103 39831
rect 15117 39797 15151 39831
rect 21465 39797 21499 39831
rect 23857 39797 23891 39831
rect 24317 39797 24351 39831
rect 8585 39593 8619 39627
rect 10609 39593 10643 39627
rect 11805 39593 11839 39627
rect 13185 39593 13219 39627
rect 14841 39593 14875 39627
rect 16497 39593 16531 39627
rect 16957 39593 16991 39627
rect 18153 39593 18187 39627
rect 23213 39525 23247 39559
rect 2053 39457 2087 39491
rect 5549 39457 5583 39491
rect 5733 39457 5767 39491
rect 6837 39457 6871 39491
rect 9689 39457 9723 39491
rect 11069 39457 11103 39491
rect 11253 39457 11287 39491
rect 12449 39457 12483 39491
rect 13829 39457 13863 39491
rect 15485 39457 15519 39491
rect 17601 39457 17635 39491
rect 18797 39457 18831 39491
rect 20361 39457 20395 39491
rect 20637 39457 20671 39491
rect 22109 39457 22143 39491
rect 22753 39457 22787 39491
rect 23765 39457 23799 39491
rect 1777 39389 1811 39423
rect 5457 39389 5491 39423
rect 12173 39389 12207 39423
rect 12265 39389 12299 39423
rect 22569 39389 22603 39423
rect 7113 39321 7147 39355
rect 9597 39321 9631 39355
rect 10977 39321 11011 39355
rect 13645 39321 13679 39355
rect 17417 39321 17451 39355
rect 22661 39321 22695 39355
rect 5089 39253 5123 39287
rect 9137 39253 9171 39287
rect 9505 39253 9539 39287
rect 13553 39253 13587 39287
rect 15209 39253 15243 39287
rect 15301 39253 15335 39287
rect 17325 39253 17359 39287
rect 18521 39253 18555 39287
rect 18613 39253 18647 39287
rect 22201 39253 22235 39287
rect 23581 39253 23615 39287
rect 23673 39253 23707 39287
rect 5641 39049 5675 39083
rect 12173 39049 12207 39083
rect 13001 39049 13035 39083
rect 13369 39049 13403 39083
rect 14197 39049 14231 39083
rect 16865 39049 16899 39083
rect 17325 39049 17359 39083
rect 18061 39049 18095 39083
rect 20637 39049 20671 39083
rect 22845 39049 22879 39083
rect 23857 39049 23891 39083
rect 6653 38981 6687 39015
rect 10977 38981 11011 39015
rect 14565 38981 14599 39015
rect 7665 38913 7699 38947
rect 8493 38913 8527 38947
rect 12541 38913 12575 38947
rect 12633 38913 12667 38947
rect 14013 38913 14047 38947
rect 14657 38913 14691 38947
rect 15577 38913 15611 38947
rect 16221 38913 16255 38947
rect 17233 38913 17267 38947
rect 18429 38913 18463 38947
rect 23765 38913 23799 38947
rect 5733 38845 5767 38879
rect 5917 38845 5951 38879
rect 7757 38845 7791 38879
rect 7941 38845 7975 38879
rect 8769 38845 8803 38879
rect 12817 38845 12851 38879
rect 13461 38845 13495 38879
rect 13645 38845 13679 38879
rect 14749 38845 14783 38879
rect 17417 38845 17451 38879
rect 18889 38845 18923 38879
rect 19165 38845 19199 38879
rect 23949 38845 23983 38879
rect 7297 38777 7331 38811
rect 11161 38777 11195 38811
rect 23397 38777 23431 38811
rect 5273 38709 5307 38743
rect 6745 38709 6779 38743
rect 10241 38709 10275 38743
rect 15393 38709 15427 38743
rect 4629 38505 4663 38539
rect 5273 38505 5307 38539
rect 9229 38505 9263 38539
rect 13737 38505 13771 38539
rect 22293 38505 22327 38539
rect 8585 38437 8619 38471
rect 18245 38437 18279 38471
rect 2053 38369 2087 38403
rect 5825 38369 5859 38403
rect 7113 38369 7147 38403
rect 9781 38369 9815 38403
rect 10977 38369 11011 38403
rect 16497 38369 16531 38403
rect 20821 38369 20855 38403
rect 23765 38369 23799 38403
rect 1777 38301 1811 38335
rect 4813 38301 4847 38335
rect 5641 38301 5675 38335
rect 6837 38301 6871 38335
rect 9597 38301 9631 38335
rect 11989 38301 12023 38335
rect 14289 38301 14323 38335
rect 20545 38301 20579 38335
rect 23489 38301 23523 38335
rect 23581 38301 23615 38335
rect 10793 38233 10827 38267
rect 12265 38233 12299 38267
rect 14565 38233 14599 38267
rect 16773 38233 16807 38267
rect 5733 38165 5767 38199
rect 9689 38165 9723 38199
rect 10425 38165 10459 38199
rect 10885 38165 10919 38199
rect 16037 38165 16071 38199
rect 23121 38165 23155 38199
rect 4353 37961 4387 37995
rect 5641 37961 5675 37995
rect 8585 37961 8619 37995
rect 9597 37961 9631 37995
rect 9689 37961 9723 37995
rect 10425 37961 10459 37995
rect 12541 37961 12575 37995
rect 23121 37961 23155 37995
rect 23213 37961 23247 37995
rect 13829 37893 13863 37927
rect 14841 37893 14875 37927
rect 20085 37893 20119 37927
rect 1777 37825 1811 37859
rect 4261 37825 4295 37859
rect 10793 37825 10827 37859
rect 11897 37825 11931 37859
rect 12909 37825 12943 37859
rect 14565 37825 14599 37859
rect 16957 37825 16991 37859
rect 2053 37757 2087 37791
rect 5733 37757 5767 37791
rect 5917 37757 5951 37791
rect 6837 37757 6871 37791
rect 7113 37757 7147 37791
rect 9873 37757 9907 37791
rect 10885 37757 10919 37791
rect 10977 37757 11011 37791
rect 13001 37757 13035 37791
rect 13093 37757 13127 37791
rect 17233 37757 17267 37791
rect 20821 37757 20855 37791
rect 23305 37757 23339 37791
rect 14013 37689 14047 37723
rect 5273 37621 5307 37655
rect 9229 37621 9263 37655
rect 16313 37621 16347 37655
rect 18705 37621 18739 37655
rect 22753 37621 22787 37655
rect 13737 37417 13771 37451
rect 18797 37417 18831 37451
rect 22293 37417 22327 37451
rect 5641 37281 5675 37315
rect 5825 37281 5859 37315
rect 6837 37281 6871 37315
rect 7021 37281 7055 37315
rect 8217 37281 8251 37315
rect 11253 37281 11287 37315
rect 12265 37281 12299 37315
rect 14657 37281 14691 37315
rect 14933 37281 14967 37315
rect 17325 37281 17359 37315
rect 23305 37281 23339 37315
rect 7941 37213 7975 37247
rect 10333 37213 10367 37247
rect 11069 37213 11103 37247
rect 11989 37213 12023 37247
rect 17049 37213 17083 37247
rect 20545 37213 20579 37247
rect 23121 37213 23155 37247
rect 23213 37213 23247 37247
rect 9597 37145 9631 37179
rect 20821 37145 20855 37179
rect 5181 37077 5215 37111
rect 5549 37077 5583 37111
rect 6377 37077 6411 37111
rect 6745 37077 6779 37111
rect 7573 37077 7607 37111
rect 8033 37077 8067 37111
rect 16405 37077 16439 37111
rect 22753 37077 22787 37111
rect 5641 36873 5675 36907
rect 7021 36873 7055 36907
rect 8401 36873 8435 36907
rect 8493 36873 8527 36907
rect 9597 36873 9631 36907
rect 10425 36873 10459 36907
rect 14749 36873 14783 36907
rect 15485 36873 15519 36907
rect 15945 36873 15979 36907
rect 22017 36873 22051 36907
rect 22385 36873 22419 36907
rect 22477 36873 22511 36907
rect 4629 36805 4663 36839
rect 10885 36805 10919 36839
rect 13001 36805 13035 36839
rect 18153 36805 18187 36839
rect 19257 36805 19291 36839
rect 1777 36737 1811 36771
rect 10793 36737 10827 36771
rect 12173 36737 12207 36771
rect 13737 36737 13771 36771
rect 14657 36737 14691 36771
rect 15853 36737 15887 36771
rect 16865 36737 16899 36771
rect 17325 36737 17359 36771
rect 18245 36737 18279 36771
rect 18981 36737 19015 36771
rect 2053 36669 2087 36703
rect 5733 36669 5767 36703
rect 5917 36669 5951 36703
rect 7113 36669 7147 36703
rect 7297 36669 7331 36703
rect 8677 36669 8711 36703
rect 9689 36669 9723 36703
rect 9781 36669 9815 36703
rect 10977 36669 11011 36703
rect 14841 36669 14875 36703
rect 16037 36669 16071 36703
rect 17417 36669 17451 36703
rect 17601 36669 17635 36703
rect 18429 36669 18463 36703
rect 22569 36669 22603 36703
rect 8033 36601 8067 36635
rect 14289 36601 14323 36635
rect 4721 36533 4755 36567
rect 5273 36533 5307 36567
rect 6653 36533 6687 36567
rect 9229 36533 9263 36567
rect 13553 36533 13587 36567
rect 16957 36533 16991 36567
rect 17785 36533 17819 36567
rect 20729 36533 20763 36567
rect 7849 36329 7883 36363
rect 11805 36329 11839 36363
rect 12449 36329 12483 36363
rect 16129 36329 16163 36363
rect 21925 36261 21959 36295
rect 6101 36193 6135 36227
rect 7205 36193 7239 36227
rect 8309 36193 8343 36227
rect 8493 36193 8527 36227
rect 11161 36193 11195 36227
rect 13093 36193 13127 36227
rect 14657 36193 14691 36227
rect 18705 36193 18739 36227
rect 20177 36193 20211 36227
rect 1777 36125 1811 36159
rect 5825 36125 5859 36159
rect 9137 36125 9171 36159
rect 14381 36125 14415 36159
rect 18521 36125 18555 36159
rect 2789 36057 2823 36091
rect 5917 36057 5951 36091
rect 7021 36057 7055 36091
rect 7113 36057 7147 36091
rect 9413 36057 9447 36091
rect 17601 36057 17635 36091
rect 18613 36057 18647 36091
rect 20453 36057 20487 36091
rect 5457 35989 5491 36023
rect 6653 35989 6687 36023
rect 8217 35989 8251 36023
rect 12817 35989 12851 36023
rect 12909 35989 12943 36023
rect 18153 35989 18187 36023
rect 7205 35785 7239 35819
rect 8033 35785 8067 35819
rect 9597 35785 9631 35819
rect 10425 35785 10459 35819
rect 14289 35785 14323 35819
rect 16037 35785 16071 35819
rect 17417 35785 17451 35819
rect 18889 35785 18923 35819
rect 5641 35717 5675 35751
rect 8401 35717 8435 35751
rect 10885 35717 10919 35751
rect 17325 35717 17359 35751
rect 18981 35717 19015 35751
rect 19993 35717 20027 35751
rect 22017 35717 22051 35751
rect 7297 35649 7331 35683
rect 9689 35649 9723 35683
rect 10793 35649 10827 35683
rect 11989 35649 12023 35683
rect 15945 35649 15979 35683
rect 5733 35581 5767 35615
rect 5917 35581 5951 35615
rect 7481 35581 7515 35615
rect 8493 35581 8527 35615
rect 8585 35581 8619 35615
rect 9781 35581 9815 35615
rect 11069 35581 11103 35615
rect 12541 35581 12575 35615
rect 12817 35581 12851 35615
rect 16221 35581 16255 35615
rect 17601 35581 17635 35615
rect 19073 35581 19107 35615
rect 19717 35581 19751 35615
rect 22845 35581 22879 35615
rect 16957 35513 16991 35547
rect 5273 35445 5307 35479
rect 6837 35445 6871 35479
rect 9229 35445 9263 35479
rect 15577 35445 15611 35479
rect 18521 35445 18555 35479
rect 21465 35445 21499 35479
rect 7849 35241 7883 35275
rect 11437 35241 11471 35275
rect 12541 35241 12575 35275
rect 13001 35241 13035 35275
rect 15577 35241 15611 35275
rect 18889 35241 18923 35275
rect 5457 35173 5491 35207
rect 2053 35105 2087 35139
rect 5917 35105 5951 35139
rect 6101 35105 6135 35139
rect 7113 35105 7147 35139
rect 7205 35105 7239 35139
rect 8401 35105 8435 35139
rect 9689 35105 9723 35139
rect 13553 35105 13587 35139
rect 14933 35105 14967 35139
rect 16129 35105 16163 35139
rect 17141 35105 17175 35139
rect 20637 35105 20671 35139
rect 21741 35105 21775 35139
rect 21833 35105 21867 35139
rect 1777 35037 1811 35071
rect 5825 35037 5859 35071
rect 7021 35037 7055 35071
rect 13369 35037 13403 35071
rect 13461 35037 13495 35071
rect 14841 35037 14875 35071
rect 20453 35037 20487 35071
rect 21649 35037 21683 35071
rect 9965 34969 9999 35003
rect 14749 34969 14783 35003
rect 17417 34969 17451 35003
rect 20545 34969 20579 35003
rect 6653 34901 6687 34935
rect 8217 34901 8251 34935
rect 8309 34901 8343 34935
rect 14381 34901 14415 34935
rect 15945 34901 15979 34935
rect 16037 34901 16071 34935
rect 20085 34901 20119 34935
rect 21281 34901 21315 34935
rect 8769 34697 8803 34731
rect 9229 34697 9263 34731
rect 16313 34697 16347 34731
rect 21465 34697 21499 34731
rect 10425 34629 10459 34663
rect 12357 34629 12391 34663
rect 17693 34629 17727 34663
rect 1777 34561 1811 34595
rect 7941 34561 7975 34595
rect 8033 34561 8067 34595
rect 9137 34561 9171 34595
rect 10333 34561 10367 34595
rect 12081 34561 12115 34595
rect 19717 34561 19751 34595
rect 2053 34493 2087 34527
rect 8125 34493 8159 34527
rect 9321 34493 9355 34527
rect 10517 34493 10551 34527
rect 13829 34493 13863 34527
rect 14565 34493 14599 34527
rect 14841 34493 14875 34527
rect 17417 34493 17451 34527
rect 7573 34357 7607 34391
rect 9965 34357 9999 34391
rect 19165 34357 19199 34391
rect 19980 34357 20014 34391
rect 8125 34153 8159 34187
rect 21281 34153 21315 34187
rect 6377 34017 6411 34051
rect 10885 34017 10919 34051
rect 11989 34017 12023 34051
rect 13185 34017 13219 34051
rect 14565 34017 14599 34051
rect 19809 34017 19843 34051
rect 10609 33949 10643 33983
rect 11805 33949 11839 33983
rect 14289 33949 14323 33983
rect 16681 33949 16715 33983
rect 19533 33949 19567 33983
rect 6653 33881 6687 33915
rect 11897 33881 11931 33915
rect 13001 33881 13035 33915
rect 13093 33881 13127 33915
rect 16957 33881 16991 33915
rect 10241 33813 10275 33847
rect 10701 33813 10735 33847
rect 11437 33813 11471 33847
rect 12633 33813 12667 33847
rect 16037 33813 16071 33847
rect 18429 33813 18463 33847
rect 8217 33609 8251 33643
rect 17233 33609 17267 33643
rect 17693 33609 17727 33643
rect 18429 33609 18463 33643
rect 18889 33609 18923 33643
rect 6653 33541 6687 33575
rect 8309 33541 8343 33575
rect 13461 33541 13495 33575
rect 16129 33541 16163 33575
rect 1777 33473 1811 33507
rect 9045 33473 9079 33507
rect 11069 33473 11103 33507
rect 13369 33473 13403 33507
rect 14565 33473 14599 33507
rect 15393 33473 15427 33507
rect 17601 33473 17635 33507
rect 18797 33473 18831 33507
rect 2053 33405 2087 33439
rect 8401 33405 8435 33439
rect 9321 33405 9355 33439
rect 13553 33405 13587 33439
rect 14657 33405 14691 33439
rect 14841 33405 14875 33439
rect 17877 33405 17911 33439
rect 19073 33405 19107 33439
rect 14197 33337 14231 33371
rect 6745 33269 6779 33303
rect 7849 33269 7883 33303
rect 13001 33269 13035 33303
rect 10517 33065 10551 33099
rect 13461 33065 13495 33099
rect 14565 33065 14599 33099
rect 15025 33065 15059 33099
rect 20821 33065 20855 33099
rect 7481 32997 7515 33031
rect 2053 32929 2087 32963
rect 8033 32929 8067 32963
rect 9965 32929 9999 32963
rect 11069 32929 11103 32963
rect 15669 32929 15703 32963
rect 1777 32861 1811 32895
rect 7849 32861 7883 32895
rect 9689 32861 9723 32895
rect 9781 32861 9815 32895
rect 11713 32861 11747 32895
rect 15393 32861 15427 32895
rect 16405 32861 16439 32895
rect 16957 32861 16991 32895
rect 5457 32793 5491 32827
rect 7941 32793 7975 32827
rect 10885 32793 10919 32827
rect 11989 32793 12023 32827
rect 17785 32793 17819 32827
rect 19533 32793 19567 32827
rect 5549 32725 5583 32759
rect 9321 32725 9355 32759
rect 10977 32725 11011 32759
rect 15485 32725 15519 32759
rect 8861 32521 8895 32555
rect 9229 32521 9263 32555
rect 9321 32521 9355 32555
rect 10425 32521 10459 32555
rect 16313 32521 16347 32555
rect 18889 32521 18923 32555
rect 21097 32521 21131 32555
rect 7205 32385 7239 32419
rect 8033 32385 8067 32419
rect 8125 32385 8159 32419
rect 10517 32385 10551 32419
rect 11897 32385 11931 32419
rect 12357 32385 12391 32419
rect 14565 32385 14599 32419
rect 8217 32317 8251 32351
rect 9413 32317 9447 32351
rect 10701 32317 10735 32351
rect 12633 32317 12667 32351
rect 14105 32317 14139 32351
rect 14841 32317 14875 32351
rect 17141 32317 17175 32351
rect 17417 32317 17451 32351
rect 19349 32317 19383 32351
rect 19625 32317 19659 32351
rect 7665 32181 7699 32215
rect 10057 32181 10091 32215
rect 10885 31977 10919 32011
rect 12252 31977 12286 32011
rect 14933 31977 14967 32011
rect 17877 31977 17911 32011
rect 2053 31841 2087 31875
rect 6653 31841 6687 31875
rect 6929 31841 6963 31875
rect 9137 31841 9171 31875
rect 13737 31841 13771 31875
rect 15393 31841 15427 31875
rect 15577 31841 15611 31875
rect 16129 31841 16163 31875
rect 16405 31841 16439 31875
rect 1777 31773 1811 31807
rect 11989 31773 12023 31807
rect 14473 31773 14507 31807
rect 9413 31705 9447 31739
rect 15301 31705 15335 31739
rect 8401 31637 8435 31671
rect 16313 31433 16347 31467
rect 19441 31433 19475 31467
rect 11161 31365 11195 31399
rect 13737 31365 13771 31399
rect 1777 31297 1811 31331
rect 17693 31297 17727 31331
rect 2053 31229 2087 31263
rect 9137 31229 9171 31263
rect 9413 31229 9447 31263
rect 11713 31229 11747 31263
rect 11989 31229 12023 31263
rect 14565 31229 14599 31263
rect 14841 31229 14875 31263
rect 17969 31229 18003 31263
rect 7849 30889 7883 30923
rect 16681 30889 16715 30923
rect 8309 30753 8343 30787
rect 8401 30753 8435 30787
rect 10241 30753 10275 30787
rect 10885 30753 10919 30787
rect 14933 30753 14967 30787
rect 8217 30685 8251 30719
rect 9505 30685 9539 30719
rect 14473 30685 14507 30719
rect 11161 30617 11195 30651
rect 15209 30617 15243 30651
rect 12633 30549 12667 30583
rect 10057 30277 10091 30311
rect 1777 30209 1811 30243
rect 11805 30209 11839 30243
rect 14381 30209 14415 30243
rect 15393 30209 15427 30243
rect 2053 30141 2087 30175
rect 8033 30141 8067 30175
rect 8309 30141 8343 30175
rect 12081 30141 12115 30175
rect 13553 30141 13587 30175
rect 14473 30141 14507 30175
rect 14657 30141 14691 30175
rect 14013 30073 14047 30107
rect 11437 29801 11471 29835
rect 14289 29801 14323 29835
rect 9689 29665 9723 29699
rect 12633 29665 12667 29699
rect 14933 29665 14967 29699
rect 1777 29597 1811 29631
rect 11897 29597 11931 29631
rect 14657 29597 14691 29631
rect 2513 29529 2547 29563
rect 9965 29529 9999 29563
rect 14749 29461 14783 29495
rect 10609 29257 10643 29291
rect 13277 29257 13311 29291
rect 7757 29189 7791 29223
rect 7481 29121 7515 29155
rect 9229 29053 9263 29087
rect 10701 29053 10735 29087
rect 10793 29053 10827 29087
rect 13369 29053 13403 29087
rect 13461 29053 13495 29087
rect 10241 28985 10275 29019
rect 12909 28917 12943 28951
rect 7849 28713 7883 28747
rect 9873 28713 9907 28747
rect 11161 28713 11195 28747
rect 12357 28645 12391 28679
rect 2053 28577 2087 28611
rect 8309 28577 8343 28611
rect 8401 28577 8435 28611
rect 10425 28577 10459 28611
rect 11713 28577 11747 28611
rect 12909 28577 12943 28611
rect 1777 28509 1811 28543
rect 8217 28509 8251 28543
rect 10333 28509 10367 28543
rect 11529 28509 11563 28543
rect 11621 28509 11655 28543
rect 10241 28441 10275 28475
rect 12725 28373 12759 28407
rect 12817 28373 12851 28407
rect 9781 28169 9815 28203
rect 9873 28169 9907 28203
rect 13001 28169 13035 28203
rect 13093 28101 13127 28135
rect 1777 28033 1811 28067
rect 2053 27965 2087 27999
rect 9965 27965 9999 27999
rect 13277 27965 13311 27999
rect 9413 27829 9447 27863
rect 12633 27829 12667 27863
rect 11713 27557 11747 27591
rect 12357 27489 12391 27523
rect 13185 27421 13219 27455
rect 12081 27353 12115 27387
rect 12173 27353 12207 27387
rect 13001 27285 13035 27319
rect 12081 27081 12115 27115
rect 1869 27013 1903 27047
rect 12173 27013 12207 27047
rect 1685 26945 1719 26979
rect 12265 26877 12299 26911
rect 11713 26741 11747 26775
rect 1869 26401 1903 26435
rect 1593 26333 1627 26367
rect 10241 25449 10275 25483
rect 1869 25313 1903 25347
rect 10885 25313 10919 25347
rect 1593 25245 1627 25279
rect 10609 25245 10643 25279
rect 11621 25245 11655 25279
rect 10701 25109 10735 25143
rect 1685 24769 1719 24803
rect 1869 24769 1903 24803
rect 32321 24701 32355 24735
rect 32597 24701 32631 24735
rect 34345 24701 34379 24735
rect 10977 24565 11011 24599
rect 10425 24361 10459 24395
rect 10977 24225 11011 24259
rect 10793 24157 10827 24191
rect 12449 24157 12483 24191
rect 10885 24021 10919 24055
rect 12081 23817 12115 23851
rect 1869 23681 1903 23715
rect 12449 23681 12483 23715
rect 13461 23681 13495 23715
rect 1593 23613 1627 23647
rect 12541 23613 12575 23647
rect 12725 23613 12759 23647
rect 11897 23273 11931 23307
rect 1869 23137 1903 23171
rect 12541 23137 12575 23171
rect 1593 23069 1627 23103
rect 12265 23069 12299 23103
rect 12357 22933 12391 22967
rect 1869 22049 1903 22083
rect 1593 21981 1627 22015
rect 1869 21505 1903 21539
rect 1593 21437 1627 21471
rect 14289 21029 14323 21063
rect 14473 20893 14507 20927
rect 15853 20893 15887 20927
rect 15669 20757 15703 20791
rect 1869 20417 1903 20451
rect 16221 20417 16255 20451
rect 30113 20417 30147 20451
rect 1593 20349 1627 20383
rect 30573 20281 30607 20315
rect 16037 20213 16071 20247
rect 30389 20213 30423 20247
rect 1869 19941 1903 19975
rect 1685 19737 1719 19771
rect 1593 18921 1627 18955
rect 1777 18717 1811 18751
rect 1593 18377 1627 18411
rect 1777 18241 1811 18275
rect 25421 17697 25455 17731
rect 27721 17697 27755 17731
rect 24961 17629 24995 17663
rect 27261 17629 27295 17663
rect 25145 17561 25179 17595
rect 27445 17561 27479 17595
rect 26433 17289 26467 17323
rect 30757 17221 30791 17255
rect 1685 17153 1719 17187
rect 17141 17153 17175 17187
rect 17325 17153 17359 17187
rect 24685 17153 24719 17187
rect 1869 17085 1903 17119
rect 24961 17085 24995 17119
rect 28917 17085 28951 17119
rect 29101 17085 29135 17119
rect 17785 16949 17819 16983
rect 1869 16677 1903 16711
rect 31033 16609 31067 16643
rect 23616 16541 23650 16575
rect 23719 16541 23753 16575
rect 32873 16541 32907 16575
rect 1685 16473 1719 16507
rect 31217 16473 31251 16507
rect 26157 15657 26191 15691
rect 1869 15589 1903 15623
rect 25881 15453 25915 15487
rect 1685 15385 1719 15419
rect 26341 15317 26375 15351
rect 24455 15113 24489 15147
rect 1869 14977 1903 15011
rect 24352 14977 24386 15011
rect 1593 14909 1627 14943
rect 25272 14365 25306 14399
rect 25375 14229 25409 14263
rect 1593 14025 1627 14059
rect 19257 14025 19291 14059
rect 21465 14025 21499 14059
rect 27307 14025 27341 14059
rect 1777 13889 1811 13923
rect 18613 13889 18647 13923
rect 19717 13889 19751 13923
rect 27204 13889 27238 13923
rect 18797 13821 18831 13855
rect 19980 13685 20014 13719
rect 24685 13481 24719 13515
rect 1777 13277 1811 13311
rect 24593 13277 24627 13311
rect 25513 13277 25547 13311
rect 1593 13141 1627 13175
rect 25053 13141 25087 13175
rect 19165 12801 19199 12835
rect 20821 12801 20855 12835
rect 19349 12733 19383 12767
rect 21005 12733 21039 12767
rect 19809 12665 19843 12699
rect 21465 12597 21499 12631
rect 1685 12121 1719 12155
rect 1777 12053 1811 12087
rect 1685 11713 1719 11747
rect 1777 11509 1811 11543
rect 22109 11305 22143 11339
rect 22477 11169 22511 11203
rect 21557 11101 21591 11135
rect 22017 11101 22051 11135
rect 1685 10625 1719 10659
rect 1777 10421 1811 10455
rect 1685 9945 1719 9979
rect 1777 9877 1811 9911
rect 1593 9129 1627 9163
rect 1777 8925 1811 8959
rect 18337 8925 18371 8959
rect 18521 8857 18555 8891
rect 1777 8449 1811 8483
rect 1593 8313 1627 8347
rect 13369 8041 13403 8075
rect 10425 7905 10459 7939
rect 13277 7837 13311 7871
rect 10701 7769 10735 7803
rect 12173 7701 12207 7735
rect 1685 7361 1719 7395
rect 1777 7157 1811 7191
rect 1869 6817 1903 6851
rect 15025 6749 15059 6783
rect 20913 6749 20947 6783
rect 22661 6749 22695 6783
rect 1685 6681 1719 6715
rect 15209 6681 15243 6715
rect 21097 6681 21131 6715
rect 22845 6681 22879 6715
rect 16957 6341 16991 6375
rect 25145 6341 25179 6375
rect 25329 6137 25363 6171
rect 17049 6069 17083 6103
rect 19533 5661 19567 5695
rect 1685 5593 1719 5627
rect 1777 5525 1811 5559
rect 19625 5525 19659 5559
rect 1869 5253 1903 5287
rect 1685 5185 1719 5219
rect 1593 4029 1627 4063
rect 1869 4029 1903 4063
rect 1593 3485 1627 3519
rect 1869 3485 1903 3519
rect 28825 3009 28859 3043
rect 46673 3009 46707 3043
rect 29285 2941 29319 2975
rect 46857 2805 46891 2839
rect 45569 2601 45603 2635
rect 7021 2465 7055 2499
rect 9689 2465 9723 2499
rect 12725 2465 12759 2499
rect 15485 2465 15519 2499
rect 19901 2465 19935 2499
rect 22661 2465 22695 2499
rect 25697 2465 25731 2499
rect 32597 2465 32631 2499
rect 38945 2465 38979 2499
rect 42901 2465 42935 2499
rect 2513 2397 2547 2431
rect 6745 2397 6779 2431
rect 9321 2397 9355 2431
rect 12357 2397 12391 2431
rect 15117 2397 15151 2431
rect 19441 2397 19475 2431
rect 22201 2397 22235 2431
rect 25237 2397 25271 2431
rect 32321 2397 32355 2431
rect 35449 2397 35483 2431
rect 35725 2397 35759 2431
rect 38669 2397 38703 2431
rect 42625 2397 42659 2431
rect 45477 2329 45511 2363
rect 2329 2261 2363 2295
<< metal1 >>
rect 10410 54680 10416 54732
rect 10468 54720 10474 54732
rect 28902 54720 28908 54732
rect 10468 54692 28908 54720
rect 10468 54680 10474 54692
rect 28902 54680 28908 54692
rect 28960 54680 28966 54732
rect 12710 54612 12716 54664
rect 12768 54652 12774 54664
rect 27706 54652 27712 54664
rect 12768 54624 27712 54652
rect 12768 54612 12774 54624
rect 27706 54612 27712 54624
rect 27764 54612 27770 54664
rect 11606 54544 11612 54596
rect 11664 54584 11670 54596
rect 32766 54584 32772 54596
rect 11664 54556 32772 54584
rect 11664 54544 11670 54556
rect 32766 54544 32772 54556
rect 32824 54544 32830 54596
rect 18690 54476 18696 54528
rect 18748 54516 18754 54528
rect 22554 54516 22560 54528
rect 18748 54488 22560 54516
rect 18748 54476 18754 54488
rect 22554 54476 22560 54488
rect 22612 54476 22618 54528
rect 1104 54426 49864 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 27950 54426
rect 28002 54374 28014 54426
rect 28066 54374 28078 54426
rect 28130 54374 28142 54426
rect 28194 54374 28206 54426
rect 28258 54374 37950 54426
rect 38002 54374 38014 54426
rect 38066 54374 38078 54426
rect 38130 54374 38142 54426
rect 38194 54374 38206 54426
rect 38258 54374 47950 54426
rect 48002 54374 48014 54426
rect 48066 54374 48078 54426
rect 48130 54374 48142 54426
rect 48194 54374 48206 54426
rect 48258 54374 49864 54426
rect 1104 54352 49864 54374
rect 19978 54272 19984 54324
rect 20036 54312 20042 54324
rect 22462 54312 22468 54324
rect 20036 54284 22468 54312
rect 20036 54272 20042 54284
rect 22462 54272 22468 54284
rect 22520 54272 22526 54324
rect 22554 54272 22560 54324
rect 22612 54272 22618 54324
rect 22646 54272 22652 54324
rect 22704 54312 22710 54324
rect 23201 54315 23259 54321
rect 23201 54312 23213 54315
rect 22704 54284 23213 54312
rect 22704 54272 22710 54284
rect 23201 54281 23213 54284
rect 23247 54281 23259 54315
rect 23201 54275 23259 54281
rect 23566 54272 23572 54324
rect 23624 54312 23630 54324
rect 26145 54315 26203 54321
rect 26145 54312 26157 54315
rect 23624 54284 26157 54312
rect 23624 54272 23630 54284
rect 26145 54281 26157 54284
rect 26191 54281 26203 54315
rect 26145 54275 26203 54281
rect 27706 54272 27712 54324
rect 27764 54312 27770 54324
rect 27801 54315 27859 54321
rect 27801 54312 27813 54315
rect 27764 54284 27813 54312
rect 27764 54272 27770 54284
rect 27801 54281 27813 54284
rect 27847 54281 27859 54315
rect 27801 54275 27859 54281
rect 28902 54272 28908 54324
rect 28960 54272 28966 54324
rect 32766 54272 32772 54324
rect 32824 54272 32830 54324
rect 3237 54247 3295 54253
rect 3237 54213 3249 54247
rect 3283 54244 3295 54247
rect 3510 54244 3516 54256
rect 3283 54216 3516 54244
rect 3283 54213 3295 54216
rect 3237 54207 3295 54213
rect 3510 54204 3516 54216
rect 3568 54204 3574 54256
rect 8389 54247 8447 54253
rect 8389 54213 8401 54247
rect 8435 54244 8447 54247
rect 8662 54244 8668 54256
rect 8435 54216 8668 54244
rect 8435 54213 8447 54216
rect 8389 54207 8447 54213
rect 8662 54204 8668 54216
rect 8720 54204 8726 54256
rect 10594 54204 10600 54256
rect 10652 54244 10658 54256
rect 10689 54247 10747 54253
rect 10689 54244 10701 54247
rect 10652 54216 10701 54244
rect 10652 54204 10658 54216
rect 10689 54213 10701 54216
rect 10735 54213 10747 54247
rect 10689 54207 10747 54213
rect 13541 54247 13599 54253
rect 13541 54213 13553 54247
rect 13587 54244 13599 54247
rect 13814 54244 13820 54256
rect 13587 54216 13820 54244
rect 13587 54213 13599 54216
rect 13541 54207 13599 54213
rect 13814 54204 13820 54216
rect 13872 54204 13878 54256
rect 15746 54204 15752 54256
rect 15804 54244 15810 54256
rect 15841 54247 15899 54253
rect 15841 54244 15853 54247
rect 15804 54216 15853 54244
rect 15804 54204 15810 54216
rect 15841 54213 15853 54216
rect 15887 54213 15899 54247
rect 15841 54207 15899 54213
rect 18693 54247 18751 54253
rect 18693 54213 18705 54247
rect 18739 54244 18751 54247
rect 18966 54244 18972 54256
rect 18739 54216 18972 54244
rect 18739 54213 18751 54216
rect 18693 54207 18751 54213
rect 18966 54204 18972 54216
rect 19024 54204 19030 54256
rect 20530 54204 20536 54256
rect 20588 54244 20594 54256
rect 20588 54216 28120 54244
rect 20588 54204 20594 54216
rect 2225 54179 2283 54185
rect 2225 54145 2237 54179
rect 2271 54176 2283 54179
rect 2314 54176 2320 54188
rect 2271 54148 2320 54176
rect 2271 54145 2283 54148
rect 2225 54139 2283 54145
rect 2314 54136 2320 54148
rect 2372 54136 2378 54188
rect 4801 54179 4859 54185
rect 4801 54145 4813 54179
rect 4847 54176 4859 54179
rect 4890 54176 4896 54188
rect 4847 54148 4896 54176
rect 4847 54145 4859 54148
rect 4801 54139 4859 54145
rect 4890 54136 4896 54148
rect 4948 54136 4954 54188
rect 7377 54179 7435 54185
rect 7377 54145 7389 54179
rect 7423 54176 7435 54179
rect 7742 54176 7748 54188
rect 7423 54148 7748 54176
rect 7423 54145 7435 54148
rect 7377 54139 7435 54145
rect 7742 54136 7748 54148
rect 7800 54136 7806 54188
rect 9953 54179 10011 54185
rect 9953 54145 9965 54179
rect 9999 54176 10011 54179
rect 10870 54176 10876 54188
rect 9999 54148 10876 54176
rect 9999 54145 10011 54148
rect 9953 54139 10011 54145
rect 10870 54136 10876 54148
rect 10928 54136 10934 54188
rect 12526 54136 12532 54188
rect 12584 54136 12590 54188
rect 12618 54136 12624 54188
rect 12676 54176 12682 54188
rect 14921 54179 14979 54185
rect 14921 54176 14933 54179
rect 12676 54148 14933 54176
rect 12676 54136 12682 54148
rect 14921 54145 14933 54148
rect 14967 54145 14979 54179
rect 14921 54139 14979 54145
rect 17681 54179 17739 54185
rect 17681 54145 17693 54179
rect 17727 54176 17739 54179
rect 17862 54176 17868 54188
rect 17727 54148 17868 54176
rect 17727 54145 17739 54148
rect 17681 54139 17739 54145
rect 17862 54136 17868 54148
rect 17920 54136 17926 54188
rect 19702 54136 19708 54188
rect 19760 54176 19766 54188
rect 20073 54179 20131 54185
rect 20346 54180 20352 54188
rect 20073 54176 20085 54179
rect 19760 54148 20085 54176
rect 19760 54136 19766 54148
rect 20073 54145 20085 54148
rect 20119 54145 20131 54179
rect 20073 54139 20131 54145
rect 20180 54152 20352 54180
rect 5442 54068 5448 54120
rect 5500 54068 5506 54120
rect 10594 54068 10600 54120
rect 10652 54108 10658 54120
rect 20180 54108 20208 54152
rect 20346 54136 20352 54152
rect 20404 54136 20410 54188
rect 22741 54179 22799 54185
rect 22741 54145 22753 54179
rect 22787 54176 22799 54179
rect 22830 54176 22836 54188
rect 22787 54148 22836 54176
rect 22787 54145 22799 54148
rect 22741 54139 22799 54145
rect 22830 54136 22836 54148
rect 22888 54136 22894 54188
rect 23385 54179 23443 54185
rect 23385 54145 23397 54179
rect 23431 54176 23443 54179
rect 23474 54176 23480 54188
rect 23431 54148 23480 54176
rect 23431 54145 23443 54148
rect 23385 54139 23443 54145
rect 23474 54136 23480 54148
rect 23532 54136 23538 54188
rect 24029 54179 24087 54185
rect 24029 54145 24041 54179
rect 24075 54176 24087 54179
rect 24118 54176 24124 54188
rect 24075 54148 24124 54176
rect 24075 54145 24087 54148
rect 24029 54139 24087 54145
rect 24118 54136 24124 54148
rect 24176 54136 24182 54188
rect 24854 54136 24860 54188
rect 24912 54176 24918 54188
rect 25041 54179 25099 54185
rect 25041 54176 25053 54179
rect 24912 54148 25053 54176
rect 24912 54136 24918 54148
rect 25041 54145 25053 54148
rect 25087 54145 25099 54179
rect 25041 54139 25099 54145
rect 25406 54136 25412 54188
rect 25464 54176 25470 54188
rect 25685 54179 25743 54185
rect 25685 54176 25697 54179
rect 25464 54148 25697 54176
rect 25464 54136 25470 54148
rect 25685 54145 25697 54148
rect 25731 54145 25743 54179
rect 25685 54139 25743 54145
rect 26234 54136 26240 54188
rect 26292 54176 26298 54188
rect 26329 54179 26387 54185
rect 26329 54176 26341 54179
rect 26292 54148 26341 54176
rect 26292 54136 26298 54148
rect 26329 54145 26341 54148
rect 26375 54145 26387 54179
rect 26329 54139 26387 54145
rect 26694 54136 26700 54188
rect 26752 54176 26758 54188
rect 27341 54179 27399 54185
rect 27341 54176 27353 54179
rect 26752 54148 27353 54176
rect 26752 54136 26758 54148
rect 27341 54145 27353 54148
rect 27387 54145 27399 54179
rect 27341 54139 27399 54145
rect 27614 54136 27620 54188
rect 27672 54176 27678 54188
rect 27985 54179 28043 54185
rect 27985 54176 27997 54179
rect 27672 54148 27997 54176
rect 27672 54136 27678 54148
rect 27985 54145 27997 54148
rect 28031 54145 28043 54179
rect 28092 54176 28120 54216
rect 28626 54204 28632 54256
rect 28684 54244 28690 54256
rect 28813 54247 28871 54253
rect 28813 54244 28825 54247
rect 28684 54216 28825 54244
rect 28684 54204 28690 54216
rect 28813 54213 28825 54216
rect 28859 54213 28871 54247
rect 28813 54207 28871 54213
rect 29270 54204 29276 54256
rect 29328 54244 29334 54256
rect 29825 54247 29883 54253
rect 29825 54244 29837 54247
rect 29328 54216 29837 54244
rect 29328 54204 29334 54216
rect 29825 54213 29837 54216
rect 29871 54213 29883 54247
rect 29825 54207 29883 54213
rect 30558 54204 30564 54256
rect 30616 54244 30622 54256
rect 30616 54216 31340 54244
rect 30616 54204 30622 54216
rect 28092 54148 29040 54176
rect 27985 54139 28043 54145
rect 10652 54080 20208 54108
rect 10652 54068 10658 54080
rect 20254 54068 20260 54120
rect 20312 54108 20318 54120
rect 20533 54111 20591 54117
rect 20533 54108 20545 54111
rect 20312 54080 20545 54108
rect 20312 54068 20318 54080
rect 20533 54077 20545 54080
rect 20579 54077 20591 54111
rect 22554 54108 22560 54120
rect 20533 54071 20591 54077
rect 20640 54080 22560 54108
rect 16482 54000 16488 54052
rect 16540 54040 16546 54052
rect 20640 54040 20668 54080
rect 22554 54068 22560 54080
rect 22612 54068 22618 54120
rect 22646 54068 22652 54120
rect 22704 54108 22710 54120
rect 22704 54080 25544 54108
rect 22704 54068 22710 54080
rect 25516 54049 25544 54080
rect 28902 54068 28908 54120
rect 28960 54068 28966 54120
rect 29012 54108 29040 54148
rect 30374 54136 30380 54188
rect 30432 54176 30438 54188
rect 31312 54185 31340 54216
rect 32490 54204 32496 54256
rect 32548 54244 32554 54256
rect 32677 54247 32735 54253
rect 32677 54244 32689 54247
rect 32548 54216 32689 54244
rect 32548 54204 32554 54216
rect 32677 54213 32689 54216
rect 32723 54213 32735 54247
rect 32677 54207 32735 54213
rect 33134 54204 33140 54256
rect 33192 54244 33198 54256
rect 33413 54247 33471 54253
rect 33413 54244 33425 54247
rect 33192 54216 33425 54244
rect 33192 54204 33198 54216
rect 33413 54213 33425 54216
rect 33459 54213 33471 54247
rect 33413 54207 33471 54213
rect 33778 54204 33784 54256
rect 33836 54244 33842 54256
rect 34149 54247 34207 54253
rect 34149 54244 34161 54247
rect 33836 54216 34161 54244
rect 33836 54204 33842 54216
rect 34149 54213 34161 54216
rect 34195 54213 34207 54247
rect 34149 54207 34207 54213
rect 34422 54204 34428 54256
rect 34480 54244 34486 54256
rect 34977 54247 35035 54253
rect 34977 54244 34989 54247
rect 34480 54216 34989 54244
rect 34480 54204 34486 54216
rect 34977 54213 34989 54216
rect 35023 54213 35035 54247
rect 34977 54207 35035 54213
rect 37642 54204 37648 54256
rect 37700 54244 37706 54256
rect 37829 54247 37887 54253
rect 37829 54244 37841 54247
rect 37700 54216 37841 54244
rect 37700 54204 37706 54216
rect 37829 54213 37841 54216
rect 37875 54213 37887 54247
rect 37829 54207 37887 54213
rect 38930 54204 38936 54256
rect 38988 54204 38994 54256
rect 42150 54204 42156 54256
rect 42208 54244 42214 54256
rect 42613 54247 42671 54253
rect 42613 54244 42625 54247
rect 42208 54216 42625 54244
rect 42208 54204 42214 54216
rect 42613 54213 42625 54216
rect 42659 54213 42671 54247
rect 42613 54207 42671 54213
rect 30653 54179 30711 54185
rect 30653 54176 30665 54179
rect 30432 54148 30665 54176
rect 30432 54136 30438 54148
rect 30653 54145 30665 54148
rect 30699 54145 30711 54179
rect 30653 54139 30711 54145
rect 31297 54179 31355 54185
rect 31297 54145 31309 54179
rect 31343 54145 31355 54179
rect 31297 54139 31355 54145
rect 35066 54136 35072 54188
rect 35124 54176 35130 54188
rect 35805 54179 35863 54185
rect 35805 54176 35817 54179
rect 35124 54148 35817 54176
rect 35124 54136 35130 54148
rect 35805 54145 35817 54148
rect 35851 54145 35863 54179
rect 35805 54139 35863 54145
rect 35894 54136 35900 54188
rect 35952 54176 35958 54188
rect 36449 54179 36507 54185
rect 36449 54176 36461 54179
rect 35952 54148 36461 54176
rect 35952 54136 35958 54148
rect 36449 54145 36461 54148
rect 36495 54145 36507 54179
rect 36449 54139 36507 54145
rect 38657 54179 38715 54185
rect 38657 54145 38669 54179
rect 38703 54176 38715 54179
rect 38948 54176 38976 54204
rect 38703 54148 38976 54176
rect 38703 54145 38715 54148
rect 38657 54139 38715 54145
rect 39574 54136 39580 54188
rect 39632 54176 39638 54188
rect 40037 54179 40095 54185
rect 40037 54176 40049 54179
rect 39632 54148 40049 54176
rect 39632 54136 39638 54148
rect 40037 54145 40049 54148
rect 40083 54145 40095 54179
rect 40037 54139 40095 54145
rect 44726 54136 44732 54188
rect 44784 54176 44790 54188
rect 45189 54179 45247 54185
rect 45189 54176 45201 54179
rect 44784 54148 45201 54176
rect 44784 54136 44790 54148
rect 45189 54145 45201 54148
rect 45235 54145 45247 54179
rect 45189 54139 45247 54145
rect 45554 54136 45560 54188
rect 45612 54176 45618 54188
rect 45925 54179 45983 54185
rect 45925 54176 45937 54179
rect 45612 54148 45937 54176
rect 45612 54136 45618 54148
rect 45925 54145 45937 54148
rect 45971 54145 45983 54179
rect 45925 54139 45983 54145
rect 46014 54136 46020 54188
rect 46072 54176 46078 54188
rect 46661 54179 46719 54185
rect 46661 54176 46673 54179
rect 46072 54148 46673 54176
rect 46072 54136 46078 54148
rect 46661 54145 46673 54148
rect 46707 54145 46719 54179
rect 46661 54139 46719 54145
rect 47302 54136 47308 54188
rect 47360 54176 47366 54188
rect 47765 54179 47823 54185
rect 47765 54176 47777 54179
rect 47360 54148 47777 54176
rect 47360 54136 47366 54148
rect 47765 54145 47777 54148
rect 47811 54145 47823 54179
rect 47765 54139 47823 54145
rect 47854 54136 47860 54188
rect 47912 54176 47918 54188
rect 48501 54179 48559 54185
rect 48501 54176 48513 54179
rect 47912 54148 48513 54176
rect 47912 54136 47918 54148
rect 48501 54145 48513 54148
rect 48547 54145 48559 54179
rect 48501 54139 48559 54145
rect 33597 54111 33655 54117
rect 33597 54108 33609 54111
rect 29012 54080 33609 54108
rect 33597 54077 33609 54080
rect 33643 54077 33655 54111
rect 33597 54071 33655 54077
rect 33704 54080 35894 54108
rect 23845 54043 23903 54049
rect 23845 54040 23857 54043
rect 16540 54012 20668 54040
rect 22066 54012 23857 54040
rect 16540 54000 16546 54012
rect 18506 53932 18512 53984
rect 18564 53972 18570 53984
rect 22066 53972 22094 54012
rect 23845 54009 23857 54012
rect 23891 54009 23903 54043
rect 23845 54003 23903 54009
rect 25501 54043 25559 54049
rect 25501 54009 25513 54043
rect 25547 54009 25559 54043
rect 28920 54040 28948 54068
rect 28920 54012 31754 54040
rect 25501 54003 25559 54009
rect 18564 53944 22094 53972
rect 18564 53932 18570 53944
rect 22462 53932 22468 53984
rect 22520 53972 22526 53984
rect 24857 53975 24915 53981
rect 24857 53972 24869 53975
rect 22520 53944 24869 53972
rect 22520 53932 22526 53944
rect 24857 53941 24869 53944
rect 24903 53941 24915 53975
rect 24857 53935 24915 53941
rect 27154 53932 27160 53984
rect 27212 53932 27218 53984
rect 29822 53932 29828 53984
rect 29880 53972 29886 53984
rect 29917 53975 29975 53981
rect 29917 53972 29929 53975
rect 29880 53944 29929 53972
rect 29880 53932 29886 53944
rect 29917 53941 29929 53944
rect 29963 53941 29975 53975
rect 29917 53935 29975 53941
rect 30466 53932 30472 53984
rect 30524 53932 30530 53984
rect 31110 53932 31116 53984
rect 31168 53932 31174 53984
rect 31726 53972 31754 54012
rect 33704 53972 33732 54080
rect 33778 54000 33784 54052
rect 33836 54040 33842 54052
rect 35621 54043 35679 54049
rect 35621 54040 35633 54043
rect 33836 54012 35633 54040
rect 33836 54000 33842 54012
rect 35621 54009 35633 54012
rect 35667 54009 35679 54043
rect 35866 54040 35894 54080
rect 38838 54068 38844 54120
rect 38896 54108 38902 54120
rect 38933 54111 38991 54117
rect 38933 54108 38945 54111
rect 38896 54080 38945 54108
rect 38896 54068 38902 54080
rect 38933 54077 38945 54080
rect 38979 54077 38991 54111
rect 38933 54071 38991 54077
rect 40310 54068 40316 54120
rect 40368 54068 40374 54120
rect 36265 54043 36323 54049
rect 36265 54040 36277 54043
rect 35866 54012 36277 54040
rect 35621 54003 35679 54009
rect 36265 54009 36277 54012
rect 36311 54009 36323 54043
rect 36265 54003 36323 54009
rect 31726 53944 33732 53972
rect 34238 53932 34244 53984
rect 34296 53932 34302 53984
rect 35066 53932 35072 53984
rect 35124 53932 35130 53984
rect 37826 53932 37832 53984
rect 37884 53972 37890 53984
rect 37921 53975 37979 53981
rect 37921 53972 37933 53975
rect 37884 53944 37933 53972
rect 37884 53932 37890 53944
rect 37921 53941 37933 53944
rect 37967 53941 37979 53975
rect 37921 53935 37979 53941
rect 43898 53932 43904 53984
rect 43956 53932 43962 53984
rect 45278 53932 45284 53984
rect 45336 53972 45342 53984
rect 45373 53975 45431 53981
rect 45373 53972 45385 53975
rect 45336 53944 45385 53972
rect 45336 53932 45342 53944
rect 45373 53941 45385 53944
rect 45419 53941 45431 53975
rect 45373 53935 45431 53941
rect 46106 53932 46112 53984
rect 46164 53932 46170 53984
rect 46842 53932 46848 53984
rect 46900 53932 46906 53984
rect 47762 53932 47768 53984
rect 47820 53972 47826 53984
rect 47949 53975 48007 53981
rect 47949 53972 47961 53975
rect 47820 53944 47961 53972
rect 47820 53932 47826 53944
rect 47949 53941 47961 53944
rect 47995 53941 48007 53975
rect 47949 53935 48007 53941
rect 48682 53932 48688 53984
rect 48740 53932 48746 53984
rect 1104 53882 49864 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 32950 53882
rect 33002 53830 33014 53882
rect 33066 53830 33078 53882
rect 33130 53830 33142 53882
rect 33194 53830 33206 53882
rect 33258 53830 42950 53882
rect 43002 53830 43014 53882
rect 43066 53830 43078 53882
rect 43130 53830 43142 53882
rect 43194 53830 43206 53882
rect 43258 53830 49864 53882
rect 1104 53808 49864 53830
rect 30374 53728 30380 53780
rect 30432 53768 30438 53780
rect 36449 53771 36507 53777
rect 36449 53768 36461 53771
rect 30432 53740 36461 53768
rect 30432 53728 30438 53740
rect 36449 53737 36461 53740
rect 36495 53737 36507 53771
rect 36449 53731 36507 53737
rect 23474 53660 23480 53712
rect 23532 53700 23538 53712
rect 31297 53703 31355 53709
rect 31297 53700 31309 53703
rect 23532 53672 31309 53700
rect 23532 53660 23538 53672
rect 31297 53669 31309 53672
rect 31343 53669 31355 53703
rect 31297 53663 31355 53669
rect 33502 53660 33508 53712
rect 33560 53700 33566 53712
rect 37093 53703 37151 53709
rect 37093 53700 37105 53703
rect 33560 53672 37105 53700
rect 33560 53660 33566 53672
rect 37093 53669 37105 53672
rect 37139 53669 37151 53703
rect 37093 53663 37151 53669
rect 2866 53592 2872 53644
rect 2924 53592 2930 53644
rect 6086 53592 6092 53644
rect 6144 53592 6150 53644
rect 7834 53592 7840 53644
rect 7892 53592 7898 53644
rect 11238 53592 11244 53644
rect 11296 53592 11302 53644
rect 13354 53592 13360 53644
rect 13412 53592 13418 53644
rect 16390 53592 16396 53644
rect 16448 53592 16454 53644
rect 18322 53592 18328 53644
rect 18380 53592 18386 53644
rect 20898 53592 20904 53644
rect 20956 53632 20962 53644
rect 21453 53635 21511 53641
rect 21453 53632 21465 53635
rect 20956 53604 21465 53632
rect 20956 53592 20962 53604
rect 21453 53601 21465 53604
rect 21499 53601 21511 53635
rect 49234 53632 49240 53644
rect 21453 53595 21511 53601
rect 48240 53604 49240 53632
rect 2225 53567 2283 53573
rect 2225 53533 2237 53567
rect 2271 53564 2283 53567
rect 4706 53564 4712 53576
rect 2271 53536 4712 53564
rect 2271 53533 2283 53536
rect 2225 53527 2283 53533
rect 4706 53524 4712 53536
rect 4764 53524 4770 53576
rect 5445 53567 5503 53573
rect 5445 53533 5457 53567
rect 5491 53564 5503 53567
rect 5534 53564 5540 53576
rect 5491 53536 5540 53564
rect 5491 53533 5503 53536
rect 5445 53527 5503 53533
rect 5534 53524 5540 53536
rect 5592 53524 5598 53576
rect 7374 53524 7380 53576
rect 7432 53524 7438 53576
rect 10689 53567 10747 53573
rect 10689 53533 10701 53567
rect 10735 53564 10747 53567
rect 11698 53564 11704 53576
rect 10735 53536 11704 53564
rect 10735 53533 10747 53536
rect 10689 53527 10747 53533
rect 11698 53524 11704 53536
rect 11756 53524 11762 53576
rect 12342 53524 12348 53576
rect 12400 53524 12406 53576
rect 13814 53524 13820 53576
rect 13872 53564 13878 53576
rect 15657 53567 15715 53573
rect 15657 53564 15669 53567
rect 13872 53536 15669 53564
rect 13872 53524 13878 53536
rect 15657 53533 15669 53536
rect 15703 53533 15715 53567
rect 15657 53527 15715 53533
rect 17681 53567 17739 53573
rect 17681 53533 17693 53567
rect 17727 53564 17739 53567
rect 20806 53564 20812 53576
rect 17727 53536 20812 53564
rect 17727 53533 17739 53536
rect 17681 53527 17739 53533
rect 20806 53524 20812 53536
rect 20864 53524 20870 53576
rect 20990 53524 20996 53576
rect 21048 53524 21054 53576
rect 22186 53524 22192 53576
rect 22244 53564 22250 53576
rect 23017 53567 23075 53573
rect 23017 53564 23029 53567
rect 22244 53536 23029 53564
rect 22244 53524 22250 53536
rect 23017 53533 23029 53536
rect 23063 53533 23075 53567
rect 23017 53527 23075 53533
rect 27798 53524 27804 53576
rect 27856 53564 27862 53576
rect 28261 53567 28319 53573
rect 28261 53564 28273 53567
rect 27856 53536 28273 53564
rect 27856 53524 27862 53536
rect 28261 53533 28273 53536
rect 28307 53533 28319 53567
rect 28261 53527 28319 53533
rect 31202 53524 31208 53576
rect 31260 53564 31266 53576
rect 31481 53567 31539 53573
rect 31481 53564 31493 53567
rect 31260 53536 31493 53564
rect 31260 53524 31266 53536
rect 31481 53533 31493 53536
rect 31527 53533 31539 53567
rect 31481 53527 31539 53533
rect 31846 53524 31852 53576
rect 31904 53564 31910 53576
rect 32125 53567 32183 53573
rect 32125 53564 32137 53567
rect 31904 53536 32137 53564
rect 31904 53524 31910 53536
rect 32125 53533 32137 53536
rect 32171 53533 32183 53567
rect 32125 53527 32183 53533
rect 36354 53524 36360 53576
rect 36412 53564 36418 53576
rect 36633 53567 36691 53573
rect 36633 53564 36645 53567
rect 36412 53536 36645 53564
rect 36412 53524 36418 53536
rect 36633 53533 36645 53536
rect 36679 53533 36691 53567
rect 36633 53527 36691 53533
rect 36998 53524 37004 53576
rect 37056 53564 37062 53576
rect 37277 53567 37335 53573
rect 37277 53564 37289 53567
rect 37056 53536 37289 53564
rect 37056 53524 37062 53536
rect 37277 53533 37289 53536
rect 37323 53533 37335 53567
rect 37277 53527 37335 53533
rect 38286 53524 38292 53576
rect 38344 53564 38350 53576
rect 38473 53567 38531 53573
rect 38473 53564 38485 53567
rect 38344 53536 38485 53564
rect 38344 53524 38350 53536
rect 38473 53533 38485 53536
rect 38519 53533 38531 53567
rect 38473 53527 38531 53533
rect 40218 53524 40224 53576
rect 40276 53564 40282 53576
rect 40497 53567 40555 53573
rect 40497 53564 40509 53567
rect 40276 53536 40509 53564
rect 40276 53524 40282 53536
rect 40497 53533 40509 53536
rect 40543 53533 40555 53567
rect 40497 53527 40555 53533
rect 44082 53524 44088 53576
rect 44140 53564 44146 53576
rect 44177 53567 44235 53573
rect 44177 53564 44189 53567
rect 44140 53536 44189 53564
rect 44140 53524 44146 53536
rect 44177 53533 44189 53536
rect 44223 53533 44235 53567
rect 44177 53527 44235 53533
rect 46658 53524 46664 53576
rect 46716 53564 46722 53576
rect 48240 53573 48268 53604
rect 49234 53592 49240 53604
rect 49292 53592 49298 53644
rect 46753 53567 46811 53573
rect 46753 53564 46765 53567
rect 46716 53536 46765 53564
rect 46716 53524 46722 53536
rect 46753 53533 46765 53536
rect 46799 53533 46811 53567
rect 46753 53527 46811 53533
rect 48225 53567 48283 53573
rect 48225 53533 48237 53567
rect 48271 53533 48283 53567
rect 48225 53527 48283 53533
rect 48590 53524 48596 53576
rect 48648 53564 48654 53576
rect 48685 53567 48743 53573
rect 48685 53564 48697 53567
rect 48648 53536 48697 53564
rect 48648 53524 48654 53536
rect 48685 53533 48697 53536
rect 48731 53533 48743 53567
rect 48685 53527 48743 53533
rect 24854 53456 24860 53508
rect 24912 53496 24918 53508
rect 24912 53468 31984 53496
rect 24912 53456 24918 53468
rect 18414 53388 18420 53440
rect 18472 53428 18478 53440
rect 22833 53431 22891 53437
rect 22833 53428 22845 53431
rect 18472 53400 22845 53428
rect 18472 53388 18478 53400
rect 22833 53397 22845 53400
rect 22879 53397 22891 53431
rect 22833 53391 22891 53397
rect 25038 53388 25044 53440
rect 25096 53428 25102 53440
rect 31956 53437 31984 53468
rect 38654 53456 38660 53508
rect 38712 53456 38718 53508
rect 28077 53431 28135 53437
rect 28077 53428 28089 53431
rect 25096 53400 28089 53428
rect 25096 53388 25102 53400
rect 28077 53397 28089 53400
rect 28123 53397 28135 53431
rect 28077 53391 28135 53397
rect 31941 53431 31999 53437
rect 31941 53397 31953 53431
rect 31987 53397 31999 53431
rect 31941 53391 31999 53397
rect 40034 53388 40040 53440
rect 40092 53428 40098 53440
rect 40313 53431 40371 53437
rect 40313 53428 40325 53431
rect 40092 53400 40325 53428
rect 40092 53388 40098 53400
rect 40313 53397 40325 53400
rect 40359 53397 40371 53431
rect 40313 53391 40371 53397
rect 44358 53388 44364 53440
rect 44416 53388 44422 53440
rect 46934 53388 46940 53440
rect 46992 53388 46998 53440
rect 47026 53388 47032 53440
rect 47084 53428 47090 53440
rect 48041 53431 48099 53437
rect 48041 53428 48053 53431
rect 47084 53400 48053 53428
rect 47084 53388 47090 53400
rect 48041 53397 48053 53400
rect 48087 53397 48099 53431
rect 48041 53391 48099 53397
rect 48866 53388 48872 53440
rect 48924 53388 48930 53440
rect 1104 53338 49864 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 27950 53338
rect 28002 53286 28014 53338
rect 28066 53286 28078 53338
rect 28130 53286 28142 53338
rect 28194 53286 28206 53338
rect 28258 53286 37950 53338
rect 38002 53286 38014 53338
rect 38066 53286 38078 53338
rect 38130 53286 38142 53338
rect 38194 53286 38206 53338
rect 38258 53286 47950 53338
rect 48002 53286 48014 53338
rect 48066 53286 48078 53338
rect 48130 53286 48142 53338
rect 48194 53286 48206 53338
rect 48258 53286 49864 53338
rect 1104 53264 49864 53286
rect 14366 53116 14372 53168
rect 14424 53156 14430 53168
rect 25038 53156 25044 53168
rect 14424 53128 25044 53156
rect 14424 53116 14430 53128
rect 25038 53116 25044 53128
rect 25096 53116 25102 53168
rect 2501 53091 2559 53097
rect 2501 53057 2513 53091
rect 2547 53088 2559 53091
rect 2682 53088 2688 53100
rect 2547 53060 2688 53088
rect 2547 53057 2559 53060
rect 2501 53051 2559 53057
rect 2682 53048 2688 53060
rect 2740 53048 2746 53100
rect 4709 53091 4767 53097
rect 4709 53057 4721 53091
rect 4755 53088 4767 53091
rect 5810 53088 5816 53100
rect 4755 53060 5816 53088
rect 4755 53057 4767 53060
rect 4709 53051 4767 53057
rect 5810 53048 5816 53060
rect 5868 53048 5874 53100
rect 7653 53091 7711 53097
rect 7653 53057 7665 53091
rect 7699 53088 7711 53091
rect 9030 53088 9036 53100
rect 7699 53060 9036 53088
rect 7699 53057 7711 53060
rect 7653 53051 7711 53057
rect 9030 53048 9036 53060
rect 9088 53048 9094 53100
rect 9950 53048 9956 53100
rect 10008 53048 10014 53100
rect 12158 53048 12164 53100
rect 12216 53088 12222 53100
rect 12621 53091 12679 53097
rect 12621 53088 12633 53091
rect 12216 53060 12633 53088
rect 12216 53048 12222 53060
rect 12621 53057 12633 53060
rect 12667 53057 12679 53091
rect 12621 53051 12679 53057
rect 15105 53091 15163 53097
rect 15105 53057 15117 53091
rect 15151 53088 15163 53091
rect 15562 53088 15568 53100
rect 15151 53060 15568 53088
rect 15151 53057 15163 53060
rect 15105 53051 15163 53057
rect 15562 53048 15568 53060
rect 15620 53048 15626 53100
rect 17770 53048 17776 53100
rect 17828 53048 17834 53100
rect 19886 53048 19892 53100
rect 19944 53048 19950 53100
rect 21542 53048 21548 53100
rect 21600 53088 21606 53100
rect 22189 53091 22247 53097
rect 22189 53088 22201 53091
rect 21600 53060 22201 53088
rect 21600 53048 21606 53060
rect 22189 53057 22201 53060
rect 22235 53057 22247 53091
rect 22189 53051 22247 53057
rect 49050 53048 49056 53100
rect 49108 53048 49114 53100
rect 2222 52980 2228 53032
rect 2280 53020 2286 53032
rect 2777 53023 2835 53029
rect 2777 53020 2789 53023
rect 2280 52992 2789 53020
rect 2280 52980 2286 52992
rect 2777 52989 2789 52992
rect 2823 52989 2835 53023
rect 2777 52983 2835 52989
rect 4798 52980 4804 53032
rect 4856 53020 4862 53032
rect 5077 53023 5135 53029
rect 5077 53020 5089 53023
rect 4856 52992 5089 53020
rect 4856 52980 4862 52992
rect 5077 52989 5089 52992
rect 5123 52989 5135 53023
rect 5077 52983 5135 52989
rect 7558 52980 7564 53032
rect 7616 53020 7622 53032
rect 7929 53023 7987 53029
rect 7929 53020 7941 53023
rect 7616 52992 7941 53020
rect 7616 52980 7622 52992
rect 7929 52989 7941 52992
rect 7975 52989 7987 53023
rect 7929 52983 7987 52989
rect 10042 52980 10048 53032
rect 10100 53020 10106 53032
rect 10229 53023 10287 53029
rect 10229 53020 10241 53023
rect 10100 52992 10241 53020
rect 10100 52980 10106 52992
rect 10229 52989 10241 52992
rect 10275 52989 10287 53023
rect 10229 52983 10287 52989
rect 12434 52980 12440 53032
rect 12492 53020 12498 53032
rect 13081 53023 13139 53029
rect 13081 53020 13093 53023
rect 12492 52992 13093 53020
rect 12492 52980 12498 52992
rect 13081 52989 13093 52992
rect 13127 52989 13139 53023
rect 15381 53023 15439 53029
rect 15381 53020 15393 53023
rect 13081 52983 13139 52989
rect 15120 52992 15393 53020
rect 15120 52964 15148 52992
rect 15381 52989 15393 52992
rect 15427 52989 15439 53023
rect 15381 52983 15439 52989
rect 17678 52980 17684 53032
rect 17736 53020 17742 53032
rect 18233 53023 18291 53029
rect 18233 53020 18245 53023
rect 17736 52992 18245 53020
rect 17736 52980 17742 52992
rect 18233 52989 18245 52992
rect 18279 52989 18291 53023
rect 18233 52983 18291 52989
rect 19610 52980 19616 53032
rect 19668 53020 19674 53032
rect 20165 53023 20223 53029
rect 20165 53020 20177 53023
rect 19668 52992 20177 53020
rect 19668 52980 19674 52992
rect 20165 52989 20177 52992
rect 20211 52989 20223 53023
rect 20165 52983 20223 52989
rect 15102 52912 15108 52964
rect 15160 52912 15166 52964
rect 21266 52844 21272 52896
rect 21324 52884 21330 52896
rect 22005 52887 22063 52893
rect 22005 52884 22017 52887
rect 21324 52856 22017 52884
rect 21324 52844 21330 52856
rect 22005 52853 22017 52856
rect 22051 52853 22063 52887
rect 22005 52847 22063 52853
rect 48774 52844 48780 52896
rect 48832 52884 48838 52896
rect 49237 52887 49295 52893
rect 49237 52884 49249 52887
rect 48832 52856 49249 52884
rect 48832 52844 48838 52856
rect 49237 52853 49249 52856
rect 49283 52853 49295 52887
rect 49237 52847 49295 52853
rect 1104 52794 49864 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 32950 52794
rect 33002 52742 33014 52794
rect 33066 52742 33078 52794
rect 33130 52742 33142 52794
rect 33194 52742 33206 52794
rect 33258 52742 42950 52794
rect 43002 52742 43014 52794
rect 43066 52742 43078 52794
rect 43130 52742 43142 52794
rect 43194 52742 43206 52794
rect 43258 52742 49864 52794
rect 1104 52720 49864 52742
rect 2774 52640 2780 52692
rect 2832 52680 2838 52692
rect 14642 52680 14648 52692
rect 2832 52652 14648 52680
rect 2832 52640 2838 52652
rect 14642 52640 14648 52652
rect 14700 52640 14706 52692
rect 20990 52640 20996 52692
rect 21048 52640 21054 52692
rect 8478 52612 8484 52624
rect 4080 52584 8484 52612
rect 1578 52504 1584 52556
rect 1636 52544 1642 52556
rect 2133 52547 2191 52553
rect 2133 52544 2145 52547
rect 1636 52516 2145 52544
rect 1636 52504 1642 52516
rect 2133 52513 2145 52516
rect 2179 52513 2191 52547
rect 2133 52507 2191 52513
rect 1857 52479 1915 52485
rect 1857 52445 1869 52479
rect 1903 52476 1915 52479
rect 4080 52476 4108 52584
rect 8478 52572 8484 52584
rect 8536 52572 8542 52624
rect 49142 52572 49148 52624
rect 49200 52612 49206 52624
rect 49237 52615 49295 52621
rect 49237 52612 49249 52615
rect 49200 52584 49249 52612
rect 49200 52572 49206 52584
rect 49237 52581 49249 52584
rect 49283 52581 49295 52615
rect 49237 52575 49295 52581
rect 4154 52504 4160 52556
rect 4212 52544 4218 52556
rect 4709 52547 4767 52553
rect 4709 52544 4721 52547
rect 4212 52516 4721 52544
rect 4212 52504 4218 52516
rect 4709 52513 4721 52516
rect 4755 52513 4767 52547
rect 4709 52507 4767 52513
rect 6730 52504 6736 52556
rect 6788 52544 6794 52556
rect 7285 52547 7343 52553
rect 7285 52544 7297 52547
rect 6788 52516 7297 52544
rect 6788 52504 6794 52516
rect 7285 52513 7297 52516
rect 7331 52513 7343 52547
rect 7285 52507 7343 52513
rect 9306 52504 9312 52556
rect 9364 52544 9370 52556
rect 9861 52547 9919 52553
rect 9861 52544 9873 52547
rect 9364 52516 9873 52544
rect 9364 52504 9370 52516
rect 9861 52513 9873 52516
rect 9907 52513 9919 52547
rect 9861 52507 9919 52513
rect 11882 52504 11888 52556
rect 11940 52544 11946 52556
rect 12437 52547 12495 52553
rect 12437 52544 12449 52547
rect 11940 52516 12449 52544
rect 11940 52504 11946 52516
rect 12437 52513 12449 52516
rect 12483 52513 12495 52547
rect 12437 52507 12495 52513
rect 14458 52504 14464 52556
rect 14516 52544 14522 52556
rect 15013 52547 15071 52553
rect 15013 52544 15025 52547
rect 14516 52516 15025 52544
rect 14516 52504 14522 52516
rect 15013 52513 15025 52516
rect 15059 52513 15071 52547
rect 15013 52507 15071 52513
rect 17034 52504 17040 52556
rect 17092 52544 17098 52556
rect 17589 52547 17647 52553
rect 17589 52544 17601 52547
rect 17092 52516 17601 52544
rect 17092 52504 17098 52516
rect 17589 52513 17601 52516
rect 17635 52513 17647 52547
rect 17589 52507 17647 52513
rect 1903 52448 4108 52476
rect 1903 52445 1915 52448
rect 1857 52439 1915 52445
rect 4246 52436 4252 52488
rect 4304 52436 4310 52488
rect 7009 52479 7067 52485
rect 7009 52445 7021 52479
rect 7055 52476 7067 52479
rect 9214 52476 9220 52488
rect 7055 52448 9220 52476
rect 7055 52445 7067 52448
rect 7009 52439 7067 52445
rect 9214 52436 9220 52448
rect 9272 52436 9278 52488
rect 9585 52479 9643 52485
rect 9585 52445 9597 52479
rect 9631 52476 9643 52479
rect 9674 52476 9680 52488
rect 9631 52448 9680 52476
rect 9631 52445 9643 52448
rect 9585 52439 9643 52445
rect 9674 52436 9680 52448
rect 9732 52436 9738 52488
rect 11790 52436 11796 52488
rect 11848 52476 11854 52488
rect 11977 52479 12035 52485
rect 11977 52476 11989 52479
rect 11848 52448 11989 52476
rect 11848 52436 11854 52448
rect 11977 52445 11989 52448
rect 12023 52445 12035 52479
rect 11977 52439 12035 52445
rect 14550 52436 14556 52488
rect 14608 52436 14614 52488
rect 16850 52436 16856 52488
rect 16908 52476 16914 52488
rect 17129 52479 17187 52485
rect 17129 52476 17141 52479
rect 16908 52448 17141 52476
rect 16908 52436 16914 52448
rect 17129 52445 17141 52448
rect 17175 52445 17187 52479
rect 17129 52439 17187 52445
rect 21174 52436 21180 52488
rect 21232 52436 21238 52488
rect 49050 52436 49056 52488
rect 49108 52436 49114 52488
rect 1104 52250 49864 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 27950 52250
rect 28002 52198 28014 52250
rect 28066 52198 28078 52250
rect 28130 52198 28142 52250
rect 28194 52198 28206 52250
rect 28258 52198 37950 52250
rect 38002 52198 38014 52250
rect 38066 52198 38078 52250
rect 38130 52198 38142 52250
rect 38194 52198 38206 52250
rect 38258 52198 47950 52250
rect 48002 52198 48014 52250
rect 48066 52198 48078 52250
rect 48130 52198 48142 52250
rect 48194 52198 48206 52250
rect 48258 52198 49864 52250
rect 1104 52176 49864 52198
rect 5810 52096 5816 52148
rect 5868 52136 5874 52148
rect 7745 52139 7803 52145
rect 7745 52136 7757 52139
rect 5868 52108 7757 52136
rect 5868 52096 5874 52108
rect 7745 52105 7757 52108
rect 7791 52105 7803 52139
rect 7745 52099 7803 52105
rect 9674 52096 9680 52148
rect 9732 52096 9738 52148
rect 9950 52096 9956 52148
rect 10008 52136 10014 52148
rect 10321 52139 10379 52145
rect 10321 52136 10333 52139
rect 10008 52108 10333 52136
rect 10008 52096 10014 52108
rect 10321 52105 10333 52108
rect 10367 52105 10379 52139
rect 10321 52099 10379 52105
rect 15562 52096 15568 52148
rect 15620 52096 15626 52148
rect 17589 52139 17647 52145
rect 17589 52105 17601 52139
rect 17635 52136 17647 52139
rect 17770 52136 17776 52148
rect 17635 52108 17776 52136
rect 17635 52105 17647 52108
rect 17589 52099 17647 52105
rect 17770 52096 17776 52108
rect 17828 52096 17834 52148
rect 17862 52096 17868 52148
rect 17920 52136 17926 52148
rect 18877 52139 18935 52145
rect 18877 52136 18889 52139
rect 17920 52108 18889 52136
rect 17920 52096 17926 52108
rect 18877 52105 18889 52108
rect 18923 52105 18935 52139
rect 18877 52099 18935 52105
rect 4890 52028 4896 52080
rect 4948 52068 4954 52080
rect 8665 52071 8723 52077
rect 8665 52068 8677 52071
rect 4948 52040 8677 52068
rect 4948 52028 4954 52040
rect 8665 52037 8677 52040
rect 8711 52037 8723 52071
rect 8665 52031 8723 52037
rect 7929 52003 7987 52009
rect 7929 51969 7941 52003
rect 7975 52000 7987 52003
rect 8386 52000 8392 52012
rect 7975 51972 8392 52000
rect 7975 51969 7987 51972
rect 7929 51963 7987 51969
rect 8386 51960 8392 51972
rect 8444 51960 8450 52012
rect 8481 52003 8539 52009
rect 8481 51969 8493 52003
rect 8527 51969 8539 52003
rect 8481 51963 8539 51969
rect 8496 51932 8524 51963
rect 9858 51960 9864 52012
rect 9916 51960 9922 52012
rect 10502 51960 10508 52012
rect 10560 51960 10566 52012
rect 14458 51960 14464 52012
rect 14516 52000 14522 52012
rect 15749 52003 15807 52009
rect 15749 52000 15761 52003
rect 14516 51972 15761 52000
rect 14516 51960 14522 51972
rect 15749 51969 15761 51972
rect 15795 51969 15807 52003
rect 15749 51963 15807 51969
rect 17678 51960 17684 52012
rect 17736 52000 17742 52012
rect 17773 52003 17831 52009
rect 17773 52000 17785 52003
rect 17736 51972 17785 52000
rect 17736 51960 17742 51972
rect 17773 51969 17785 51972
rect 17819 51969 17831 52003
rect 17773 51963 17831 51969
rect 18966 51960 18972 52012
rect 19024 52000 19030 52012
rect 19061 52003 19119 52009
rect 19061 52000 19073 52003
rect 19024 51972 19073 52000
rect 19024 51960 19030 51972
rect 19061 51969 19073 51972
rect 19107 51969 19119 52003
rect 19061 51963 19119 51969
rect 10686 51932 10692 51944
rect 8496 51904 10692 51932
rect 10686 51892 10692 51904
rect 10744 51892 10750 51944
rect 16298 51756 16304 51808
rect 16356 51796 16362 51808
rect 17037 51799 17095 51805
rect 17037 51796 17049 51799
rect 16356 51768 17049 51796
rect 16356 51756 16362 51768
rect 17037 51765 17049 51768
rect 17083 51765 17095 51799
rect 17037 51759 17095 51765
rect 1104 51706 49864 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 32950 51706
rect 33002 51654 33014 51706
rect 33066 51654 33078 51706
rect 33130 51654 33142 51706
rect 33194 51654 33206 51706
rect 33258 51654 42950 51706
rect 43002 51654 43014 51706
rect 43066 51654 43078 51706
rect 43130 51654 43142 51706
rect 43194 51654 43206 51706
rect 43258 51654 49864 51706
rect 1104 51632 49864 51654
rect 7374 51552 7380 51604
rect 7432 51592 7438 51604
rect 7653 51595 7711 51601
rect 7653 51592 7665 51595
rect 7432 51564 7665 51592
rect 7432 51552 7438 51564
rect 7653 51561 7665 51564
rect 7699 51561 7711 51595
rect 7653 51555 7711 51561
rect 9214 51552 9220 51604
rect 9272 51552 9278 51604
rect 10870 51552 10876 51604
rect 10928 51552 10934 51604
rect 13541 51595 13599 51601
rect 13541 51561 13553 51595
rect 13587 51592 13599 51595
rect 14550 51592 14556 51604
rect 13587 51564 14556 51592
rect 13587 51561 13599 51564
rect 13541 51555 13599 51561
rect 14550 51552 14556 51564
rect 14608 51552 14614 51604
rect 14642 51552 14648 51604
rect 14700 51592 14706 51604
rect 18598 51592 18604 51604
rect 14700 51564 18604 51592
rect 14700 51552 14706 51564
rect 18598 51552 18604 51564
rect 18656 51552 18662 51604
rect 5534 51484 5540 51536
rect 5592 51524 5598 51536
rect 8573 51527 8631 51533
rect 8573 51524 8585 51527
rect 5592 51496 8585 51524
rect 5592 51484 5598 51496
rect 8573 51493 8585 51496
rect 8619 51493 8631 51527
rect 8573 51487 8631 51493
rect 17310 51484 17316 51536
rect 17368 51524 17374 51536
rect 17589 51527 17647 51533
rect 17589 51524 17601 51527
rect 17368 51496 17601 51524
rect 17368 51484 17374 51496
rect 17589 51493 17601 51496
rect 17635 51524 17647 51527
rect 17635 51496 20116 51524
rect 17635 51493 17647 51496
rect 17589 51487 17647 51493
rect 1302 51416 1308 51468
rect 1360 51456 1366 51468
rect 2041 51459 2099 51465
rect 2041 51456 2053 51459
rect 1360 51428 2053 51456
rect 1360 51416 1366 51428
rect 2041 51425 2053 51428
rect 2087 51425 2099 51459
rect 2041 51419 2099 51425
rect 3326 51416 3332 51468
rect 3384 51456 3390 51468
rect 3384 51428 11744 51456
rect 3384 51416 3390 51428
rect 1765 51391 1823 51397
rect 1765 51357 1777 51391
rect 1811 51388 1823 51391
rect 5166 51388 5172 51400
rect 1811 51360 5172 51388
rect 1811 51357 1823 51360
rect 1765 51351 1823 51357
rect 5166 51348 5172 51360
rect 5224 51348 5230 51400
rect 7834 51348 7840 51400
rect 7892 51348 7898 51400
rect 9401 51391 9459 51397
rect 9401 51357 9413 51391
rect 9447 51388 9459 51391
rect 10962 51388 10968 51400
rect 9447 51360 10968 51388
rect 9447 51357 9459 51360
rect 9401 51351 9459 51357
rect 10962 51348 10968 51360
rect 11020 51348 11026 51400
rect 11054 51348 11060 51400
rect 11112 51348 11118 51400
rect 8389 51323 8447 51329
rect 8389 51289 8401 51323
rect 8435 51320 8447 51323
rect 10778 51320 10784 51332
rect 8435 51292 10784 51320
rect 8435 51289 8447 51292
rect 8389 51283 8447 51289
rect 10778 51280 10784 51292
rect 10836 51280 10842 51332
rect 11716 51320 11744 51428
rect 13354 51416 13360 51468
rect 13412 51456 13418 51468
rect 14921 51459 14979 51465
rect 14921 51456 14933 51459
rect 13412 51428 14933 51456
rect 13412 51416 13418 51428
rect 14921 51425 14933 51428
rect 14967 51425 14979 51459
rect 14921 51419 14979 51425
rect 16114 51416 16120 51468
rect 16172 51456 16178 51468
rect 18601 51459 18659 51465
rect 18601 51456 18613 51459
rect 16172 51428 18613 51456
rect 16172 51416 16178 51428
rect 18601 51425 18613 51428
rect 18647 51425 18659 51459
rect 18601 51419 18659 51425
rect 19978 51416 19984 51468
rect 20036 51416 20042 51468
rect 20088 51465 20116 51496
rect 20073 51459 20131 51465
rect 20073 51425 20085 51459
rect 20119 51425 20131 51459
rect 20073 51419 20131 51425
rect 13725 51391 13783 51397
rect 13725 51357 13737 51391
rect 13771 51388 13783 51391
rect 14182 51388 14188 51400
rect 13771 51360 14188 51388
rect 13771 51357 13783 51360
rect 13725 51351 13783 51357
rect 14182 51348 14188 51360
rect 14240 51348 14246 51400
rect 15838 51348 15844 51400
rect 15896 51348 15902 51400
rect 18506 51348 18512 51400
rect 18564 51348 18570 51400
rect 15654 51320 15660 51332
rect 11716 51292 15660 51320
rect 15654 51280 15660 51292
rect 15712 51280 15718 51332
rect 16022 51280 16028 51332
rect 16080 51320 16086 51332
rect 16117 51323 16175 51329
rect 16117 51320 16129 51323
rect 16080 51292 16129 51320
rect 16080 51280 16086 51292
rect 16117 51289 16129 51292
rect 16163 51289 16175 51323
rect 17402 51320 17408 51332
rect 17342 51292 17408 51320
rect 16117 51283 16175 51289
rect 17402 51280 17408 51292
rect 17460 51280 17466 51332
rect 17494 51212 17500 51264
rect 17552 51252 17558 51264
rect 18049 51255 18107 51261
rect 18049 51252 18061 51255
rect 17552 51224 18061 51252
rect 17552 51212 17558 51224
rect 18049 51221 18061 51224
rect 18095 51221 18107 51255
rect 18049 51215 18107 51221
rect 18417 51255 18475 51261
rect 18417 51221 18429 51255
rect 18463 51252 18475 51255
rect 18598 51252 18604 51264
rect 18463 51224 18604 51252
rect 18463 51221 18475 51224
rect 18417 51215 18475 51221
rect 18598 51212 18604 51224
rect 18656 51212 18662 51264
rect 19518 51212 19524 51264
rect 19576 51212 19582 51264
rect 19610 51212 19616 51264
rect 19668 51252 19674 51264
rect 19889 51255 19947 51261
rect 19889 51252 19901 51255
rect 19668 51224 19901 51252
rect 19668 51212 19674 51224
rect 19889 51221 19901 51224
rect 19935 51252 19947 51255
rect 20438 51252 20444 51264
rect 19935 51224 20444 51252
rect 19935 51221 19947 51224
rect 19889 51215 19947 51221
rect 20438 51212 20444 51224
rect 20496 51212 20502 51264
rect 1104 51162 49864 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 27950 51162
rect 28002 51110 28014 51162
rect 28066 51110 28078 51162
rect 28130 51110 28142 51162
rect 28194 51110 28206 51162
rect 28258 51110 37950 51162
rect 38002 51110 38014 51162
rect 38066 51110 38078 51162
rect 38130 51110 38142 51162
rect 38194 51110 38206 51162
rect 38258 51110 47950 51162
rect 48002 51110 48014 51162
rect 48066 51110 48078 51162
rect 48130 51110 48142 51162
rect 48194 51110 48206 51162
rect 48258 51110 49864 51162
rect 1104 51088 49864 51110
rect 7742 51008 7748 51060
rect 7800 51048 7806 51060
rect 8389 51051 8447 51057
rect 8389 51048 8401 51051
rect 7800 51020 8401 51048
rect 7800 51008 7806 51020
rect 8389 51017 8401 51020
rect 8435 51017 8447 51051
rect 8389 51011 8447 51017
rect 9030 51008 9036 51060
rect 9088 51008 9094 51060
rect 12161 51051 12219 51057
rect 12161 51017 12173 51051
rect 12207 51048 12219 51051
rect 12342 51048 12348 51060
rect 12207 51020 12348 51048
rect 12207 51017 12219 51020
rect 12161 51011 12219 51017
rect 12342 51008 12348 51020
rect 12400 51008 12406 51060
rect 12526 51008 12532 51060
rect 12584 51048 12590 51060
rect 12805 51051 12863 51057
rect 12805 51048 12817 51051
rect 12584 51020 12817 51048
rect 12584 51008 12590 51020
rect 12805 51017 12817 51020
rect 12851 51017 12863 51051
rect 15838 51048 15844 51060
rect 12805 51011 12863 51017
rect 14568 51020 15844 51048
rect 13541 50983 13599 50989
rect 13541 50949 13553 50983
rect 13587 50980 13599 50983
rect 14366 50980 14372 50992
rect 13587 50952 14372 50980
rect 13587 50949 13599 50952
rect 13541 50943 13599 50949
rect 14366 50940 14372 50952
rect 14424 50940 14430 50992
rect 1765 50915 1823 50921
rect 1765 50881 1777 50915
rect 1811 50912 1823 50915
rect 3326 50912 3332 50924
rect 1811 50884 3332 50912
rect 1811 50881 1823 50884
rect 1765 50875 1823 50881
rect 3326 50872 3332 50884
rect 3384 50872 3390 50924
rect 7650 50872 7656 50924
rect 7708 50912 7714 50924
rect 8573 50915 8631 50921
rect 8573 50912 8585 50915
rect 7708 50884 8585 50912
rect 7708 50872 7714 50884
rect 8573 50881 8585 50884
rect 8619 50881 8631 50915
rect 8573 50875 8631 50881
rect 9214 50872 9220 50924
rect 9272 50872 9278 50924
rect 12342 50872 12348 50924
rect 12400 50872 12406 50924
rect 12802 50872 12808 50924
rect 12860 50912 12866 50924
rect 12989 50915 13047 50921
rect 12989 50912 13001 50915
rect 12860 50884 13001 50912
rect 12860 50872 12866 50884
rect 12989 50881 13001 50884
rect 13035 50881 13047 50915
rect 12989 50875 13047 50881
rect 1302 50804 1308 50856
rect 1360 50844 1366 50856
rect 2041 50847 2099 50853
rect 2041 50844 2053 50847
rect 1360 50816 2053 50844
rect 1360 50804 1366 50816
rect 2041 50813 2053 50816
rect 2087 50813 2099 50847
rect 2041 50807 2099 50813
rect 14090 50804 14096 50856
rect 14148 50844 14154 50856
rect 14568 50853 14596 51020
rect 15838 51008 15844 51020
rect 15896 51048 15902 51060
rect 15896 51020 17080 51048
rect 15896 51008 15902 51020
rect 15286 50940 15292 50992
rect 15344 50940 15350 50992
rect 17052 50924 17080 51020
rect 17402 51008 17408 51060
rect 17460 51048 17466 51060
rect 17460 51020 18460 51048
rect 17460 51008 17466 51020
rect 17310 50940 17316 50992
rect 17368 50940 17374 50992
rect 18432 50924 18460 51020
rect 20806 51008 20812 51060
rect 20864 51048 20870 51060
rect 20993 51051 21051 51057
rect 20993 51048 21005 51051
rect 20864 51020 21005 51048
rect 20864 51008 20870 51020
rect 20993 51017 21005 51020
rect 21039 51017 21051 51051
rect 20993 51011 21051 51017
rect 23474 51008 23480 51060
rect 23532 51008 23538 51060
rect 33410 51008 33416 51060
rect 33468 51048 33474 51060
rect 33468 51020 39160 51048
rect 33468 51008 33474 51020
rect 20257 50983 20315 50989
rect 20257 50949 20269 50983
rect 20303 50980 20315 50983
rect 22646 50980 22652 50992
rect 20303 50952 22652 50980
rect 20303 50949 20315 50952
rect 20257 50943 20315 50949
rect 22646 50940 22652 50952
rect 22704 50940 22710 50992
rect 39132 50980 39160 51020
rect 43898 50980 43904 50992
rect 39054 50952 43904 50980
rect 43898 50940 43904 50952
rect 43956 50940 43962 50992
rect 17034 50872 17040 50924
rect 17092 50872 17098 50924
rect 18414 50872 18420 50924
rect 18472 50872 18478 50924
rect 19426 50872 19432 50924
rect 19484 50912 19490 50924
rect 20162 50912 20168 50924
rect 19484 50884 20168 50912
rect 19484 50872 19490 50884
rect 20162 50872 20168 50884
rect 20220 50872 20226 50924
rect 21177 50915 21235 50921
rect 21177 50881 21189 50915
rect 21223 50912 21235 50915
rect 21450 50912 21456 50924
rect 21223 50884 21456 50912
rect 21223 50881 21235 50884
rect 21177 50875 21235 50881
rect 21450 50872 21456 50884
rect 21508 50872 21514 50924
rect 21542 50872 21548 50924
rect 21600 50912 21606 50924
rect 23385 50915 23443 50921
rect 23385 50912 23397 50915
rect 21600 50884 23397 50912
rect 21600 50872 21606 50884
rect 23385 50881 23397 50884
rect 23431 50912 23443 50915
rect 26142 50912 26148 50924
rect 23431 50884 26148 50912
rect 23431 50881 23443 50884
rect 23385 50875 23443 50881
rect 26142 50872 26148 50884
rect 26200 50872 26206 50924
rect 14553 50847 14611 50853
rect 14553 50844 14565 50847
rect 14148 50816 14565 50844
rect 14148 50804 14154 50816
rect 14553 50813 14565 50816
rect 14599 50813 14611 50847
rect 14553 50807 14611 50813
rect 14829 50847 14887 50853
rect 14829 50813 14841 50847
rect 14875 50844 14887 50847
rect 16114 50844 16120 50856
rect 14875 50816 16120 50844
rect 14875 50813 14887 50816
rect 14829 50807 14887 50813
rect 16114 50804 16120 50816
rect 16172 50804 16178 50856
rect 17770 50804 17776 50856
rect 17828 50844 17834 50856
rect 20349 50847 20407 50853
rect 20349 50844 20361 50847
rect 17828 50816 20361 50844
rect 17828 50804 17834 50816
rect 20349 50813 20361 50816
rect 20395 50813 20407 50847
rect 20349 50807 20407 50813
rect 20438 50804 20444 50856
rect 20496 50844 20502 50856
rect 20496 50816 23244 50844
rect 20496 50804 20502 50816
rect 20162 50736 20168 50788
rect 20220 50776 20226 50788
rect 23216 50776 23244 50816
rect 23290 50804 23296 50856
rect 23348 50844 23354 50856
rect 23569 50847 23627 50853
rect 23569 50844 23581 50847
rect 23348 50816 23581 50844
rect 23348 50804 23354 50816
rect 23569 50813 23581 50816
rect 23615 50813 23627 50847
rect 23569 50807 23627 50813
rect 37550 50804 37556 50856
rect 37608 50804 37614 50856
rect 37829 50847 37887 50853
rect 37829 50813 37841 50847
rect 37875 50844 37887 50847
rect 47026 50844 47032 50856
rect 37875 50816 47032 50844
rect 37875 50813 37887 50816
rect 37829 50807 37887 50813
rect 47026 50804 47032 50816
rect 47084 50804 47090 50856
rect 24762 50776 24768 50788
rect 20220 50748 23152 50776
rect 23216 50748 24768 50776
rect 20220 50736 20226 50748
rect 13630 50668 13636 50720
rect 13688 50668 13694 50720
rect 15838 50668 15844 50720
rect 15896 50708 15902 50720
rect 16022 50708 16028 50720
rect 15896 50680 16028 50708
rect 15896 50668 15902 50680
rect 16022 50668 16028 50680
rect 16080 50708 16086 50720
rect 16301 50711 16359 50717
rect 16301 50708 16313 50711
rect 16080 50680 16313 50708
rect 16080 50668 16086 50680
rect 16301 50677 16313 50680
rect 16347 50677 16359 50711
rect 16301 50671 16359 50677
rect 17402 50668 17408 50720
rect 17460 50708 17466 50720
rect 18785 50711 18843 50717
rect 18785 50708 18797 50711
rect 17460 50680 18797 50708
rect 17460 50668 17466 50680
rect 18785 50677 18797 50680
rect 18831 50677 18843 50711
rect 18785 50671 18843 50677
rect 19518 50668 19524 50720
rect 19576 50708 19582 50720
rect 19797 50711 19855 50717
rect 19797 50708 19809 50711
rect 19576 50680 19809 50708
rect 19576 50668 19582 50680
rect 19797 50677 19809 50680
rect 19843 50677 19855 50711
rect 19797 50671 19855 50677
rect 22462 50668 22468 50720
rect 22520 50708 22526 50720
rect 23017 50711 23075 50717
rect 23017 50708 23029 50711
rect 22520 50680 23029 50708
rect 22520 50668 22526 50680
rect 23017 50677 23029 50680
rect 23063 50677 23075 50711
rect 23124 50708 23152 50748
rect 24762 50736 24768 50748
rect 24820 50736 24826 50788
rect 24946 50708 24952 50720
rect 23124 50680 24952 50708
rect 23017 50671 23075 50677
rect 24946 50668 24952 50680
rect 25004 50668 25010 50720
rect 27614 50668 27620 50720
rect 27672 50708 27678 50720
rect 39301 50711 39359 50717
rect 39301 50708 39313 50711
rect 27672 50680 39313 50708
rect 27672 50668 27678 50680
rect 39301 50677 39313 50680
rect 39347 50677 39359 50711
rect 39301 50671 39359 50677
rect 1104 50618 49864 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 32950 50618
rect 33002 50566 33014 50618
rect 33066 50566 33078 50618
rect 33130 50566 33142 50618
rect 33194 50566 33206 50618
rect 33258 50566 42950 50618
rect 43002 50566 43014 50618
rect 43066 50566 43078 50618
rect 43130 50566 43142 50618
rect 43194 50566 43206 50618
rect 43258 50566 49864 50618
rect 1104 50544 49864 50566
rect 11698 50464 11704 50516
rect 11756 50464 11762 50516
rect 13541 50507 13599 50513
rect 13541 50473 13553 50507
rect 13587 50504 13599 50507
rect 13587 50476 15700 50504
rect 13587 50473 13599 50476
rect 13541 50467 13599 50473
rect 1578 50396 1584 50448
rect 1636 50436 1642 50448
rect 13630 50436 13636 50448
rect 1636 50408 13636 50436
rect 1636 50396 1642 50408
rect 13630 50396 13636 50408
rect 13688 50396 13694 50448
rect 15672 50436 15700 50476
rect 16114 50464 16120 50516
rect 16172 50464 16178 50516
rect 17586 50464 17592 50516
rect 17644 50504 17650 50516
rect 19610 50504 19616 50516
rect 17644 50476 19616 50504
rect 17644 50464 17650 50476
rect 19610 50464 19616 50476
rect 19668 50464 19674 50516
rect 20070 50464 20076 50516
rect 20128 50504 20134 50516
rect 21542 50504 21548 50516
rect 20128 50476 21548 50504
rect 20128 50464 20134 50476
rect 21542 50464 21548 50476
rect 21600 50464 21606 50516
rect 21726 50464 21732 50516
rect 21784 50504 21790 50516
rect 23293 50507 23351 50513
rect 23293 50504 23305 50507
rect 21784 50476 23305 50504
rect 21784 50464 21790 50476
rect 23293 50473 23305 50476
rect 23339 50473 23351 50507
rect 23293 50467 23351 50473
rect 16850 50436 16856 50448
rect 15672 50408 16856 50436
rect 16850 50396 16856 50408
rect 16908 50396 16914 50448
rect 16206 50328 16212 50380
rect 16264 50368 16270 50380
rect 17402 50368 17408 50380
rect 16264 50340 17408 50368
rect 16264 50328 16270 50340
rect 17402 50328 17408 50340
rect 17460 50328 17466 50380
rect 18598 50328 18604 50380
rect 18656 50368 18662 50380
rect 20070 50368 20076 50380
rect 18656 50340 20076 50368
rect 18656 50328 18662 50340
rect 20070 50328 20076 50340
rect 20128 50328 20134 50380
rect 20257 50371 20315 50377
rect 20257 50337 20269 50371
rect 20303 50337 20315 50371
rect 20257 50331 20315 50337
rect 11882 50260 11888 50312
rect 11940 50260 11946 50312
rect 14090 50260 14096 50312
rect 14148 50300 14154 50312
rect 14369 50303 14427 50309
rect 14369 50300 14381 50303
rect 14148 50272 14381 50300
rect 14148 50260 14154 50272
rect 14369 50269 14381 50272
rect 14415 50269 14427 50303
rect 14369 50263 14427 50269
rect 17034 50260 17040 50312
rect 17092 50300 17098 50312
rect 17129 50303 17187 50309
rect 17129 50300 17141 50303
rect 17092 50272 17141 50300
rect 17092 50260 17098 50272
rect 17129 50269 17141 50272
rect 17175 50269 17187 50303
rect 17129 50263 17187 50269
rect 18966 50260 18972 50312
rect 19024 50300 19030 50312
rect 20272 50300 20300 50331
rect 21542 50328 21548 50380
rect 21600 50368 21606 50380
rect 21600 50340 22324 50368
rect 21600 50328 21606 50340
rect 19024 50272 20300 50300
rect 19024 50260 19030 50272
rect 20898 50260 20904 50312
rect 20956 50260 20962 50312
rect 22296 50300 22324 50340
rect 22646 50328 22652 50380
rect 22704 50368 22710 50380
rect 23845 50371 23903 50377
rect 23845 50368 23857 50371
rect 22704 50340 23857 50368
rect 22704 50328 22710 50340
rect 23845 50337 23857 50340
rect 23891 50337 23903 50371
rect 23845 50331 23903 50337
rect 23382 50300 23388 50312
rect 22296 50286 23388 50300
rect 22310 50272 23388 50286
rect 23382 50260 23388 50272
rect 23440 50300 23446 50312
rect 23753 50303 23811 50309
rect 23440 50272 23704 50300
rect 23440 50260 23446 50272
rect 13449 50235 13507 50241
rect 13449 50201 13461 50235
rect 13495 50201 13507 50235
rect 13449 50195 13507 50201
rect 13464 50164 13492 50195
rect 13630 50192 13636 50244
rect 13688 50232 13694 50244
rect 14645 50235 14703 50241
rect 14645 50232 14657 50235
rect 13688 50204 14657 50232
rect 13688 50192 13694 50204
rect 14645 50201 14657 50204
rect 14691 50201 14703 50235
rect 14645 50195 14703 50201
rect 15194 50192 15200 50244
rect 15252 50192 15258 50244
rect 18414 50192 18420 50244
rect 18472 50192 18478 50244
rect 20070 50192 20076 50244
rect 20128 50192 20134 50244
rect 20254 50192 20260 50244
rect 20312 50232 20318 50244
rect 21177 50235 21235 50241
rect 21177 50232 21189 50235
rect 20312 50204 21189 50232
rect 20312 50192 20318 50204
rect 21177 50201 21189 50204
rect 21223 50232 21235 50235
rect 21450 50232 21456 50244
rect 21223 50204 21456 50232
rect 21223 50201 21235 50204
rect 21177 50195 21235 50201
rect 21450 50192 21456 50204
rect 21508 50192 21514 50244
rect 23566 50232 23572 50244
rect 22572 50204 23572 50232
rect 15562 50164 15568 50176
rect 13464 50136 15568 50164
rect 15562 50124 15568 50136
rect 15620 50124 15626 50176
rect 17770 50124 17776 50176
rect 17828 50164 17834 50176
rect 18877 50167 18935 50173
rect 18877 50164 18889 50167
rect 17828 50136 18889 50164
rect 17828 50124 17834 50136
rect 18877 50133 18889 50136
rect 18923 50133 18935 50167
rect 18877 50127 18935 50133
rect 19610 50124 19616 50176
rect 19668 50164 19674 50176
rect 19705 50167 19763 50173
rect 19705 50164 19717 50167
rect 19668 50136 19717 50164
rect 19668 50124 19674 50136
rect 19705 50133 19717 50136
rect 19751 50133 19763 50167
rect 19705 50127 19763 50133
rect 20165 50167 20223 50173
rect 20165 50133 20177 50167
rect 20211 50164 20223 50167
rect 22572 50164 22600 50204
rect 23566 50192 23572 50204
rect 23624 50192 23630 50244
rect 23676 50232 23704 50272
rect 23753 50269 23765 50303
rect 23799 50300 23811 50303
rect 24854 50300 24860 50312
rect 23799 50272 24860 50300
rect 23799 50269 23811 50272
rect 23753 50263 23811 50269
rect 24854 50260 24860 50272
rect 24912 50260 24918 50312
rect 49050 50260 49056 50312
rect 49108 50260 49114 50312
rect 31202 50232 31208 50244
rect 23676 50204 31208 50232
rect 31202 50192 31208 50204
rect 31260 50192 31266 50244
rect 20211 50136 22600 50164
rect 20211 50133 20223 50136
rect 20165 50127 20223 50133
rect 22646 50124 22652 50176
rect 22704 50124 22710 50176
rect 23658 50124 23664 50176
rect 23716 50124 23722 50176
rect 49234 50124 49240 50176
rect 49292 50124 49298 50176
rect 1104 50074 49864 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 27950 50074
rect 28002 50022 28014 50074
rect 28066 50022 28078 50074
rect 28130 50022 28142 50074
rect 28194 50022 28206 50074
rect 28258 50022 37950 50074
rect 38002 50022 38014 50074
rect 38066 50022 38078 50074
rect 38130 50022 38142 50074
rect 38194 50022 38206 50074
rect 38258 50022 47950 50074
rect 48002 50022 48014 50074
rect 48066 50022 48078 50074
rect 48130 50022 48142 50074
rect 48194 50022 48206 50074
rect 48258 50022 49864 50074
rect 1104 50000 49864 50022
rect 13722 49920 13728 49972
rect 13780 49960 13786 49972
rect 15841 49963 15899 49969
rect 15841 49960 15853 49963
rect 13780 49932 15853 49960
rect 13780 49920 13786 49932
rect 15841 49929 15853 49932
rect 15887 49929 15899 49963
rect 15841 49923 15899 49929
rect 16574 49920 16580 49972
rect 16632 49960 16638 49972
rect 17129 49963 17187 49969
rect 17129 49960 17141 49963
rect 16632 49932 17141 49960
rect 16632 49920 16638 49932
rect 17129 49929 17141 49932
rect 17175 49929 17187 49963
rect 17129 49923 17187 49929
rect 17589 49963 17647 49969
rect 17589 49929 17601 49963
rect 17635 49960 17647 49963
rect 18690 49960 18696 49972
rect 17635 49932 18696 49960
rect 17635 49929 17647 49932
rect 17589 49923 17647 49929
rect 18690 49920 18696 49932
rect 18748 49920 18754 49972
rect 20990 49960 20996 49972
rect 19904 49932 20996 49960
rect 12158 49852 12164 49904
rect 12216 49852 12222 49904
rect 12710 49852 12716 49904
rect 12768 49852 12774 49904
rect 13633 49895 13691 49901
rect 13633 49861 13645 49895
rect 13679 49892 13691 49895
rect 13814 49892 13820 49904
rect 13679 49864 13820 49892
rect 13679 49861 13691 49864
rect 13633 49855 13691 49861
rect 13814 49852 13820 49864
rect 13872 49852 13878 49904
rect 14826 49852 14832 49904
rect 14884 49852 14890 49904
rect 17034 49852 17040 49904
rect 17092 49892 17098 49904
rect 19061 49895 19119 49901
rect 19061 49892 19073 49895
rect 17092 49864 19073 49892
rect 17092 49852 17098 49864
rect 19061 49861 19073 49864
rect 19107 49861 19119 49895
rect 19904 49892 19932 49932
rect 20990 49920 20996 49932
rect 21048 49920 21054 49972
rect 22738 49920 22744 49972
rect 22796 49960 22802 49972
rect 23385 49963 23443 49969
rect 23385 49960 23397 49963
rect 22796 49932 23397 49960
rect 22796 49920 22802 49932
rect 23385 49929 23397 49932
rect 23431 49929 23443 49963
rect 23385 49923 23443 49929
rect 23845 49963 23903 49969
rect 23845 49929 23857 49963
rect 23891 49960 23903 49963
rect 31110 49960 31116 49972
rect 23891 49932 31116 49960
rect 23891 49929 23903 49932
rect 23845 49923 23903 49929
rect 31110 49920 31116 49932
rect 31168 49920 31174 49972
rect 31202 49920 31208 49972
rect 31260 49960 31266 49972
rect 33410 49960 33416 49972
rect 31260 49932 33416 49960
rect 31260 49920 31266 49932
rect 33410 49920 33416 49932
rect 33468 49960 33474 49972
rect 33686 49960 33692 49972
rect 33468 49932 33692 49960
rect 33468 49920 33474 49932
rect 33686 49920 33692 49932
rect 33744 49920 33750 49972
rect 21542 49892 21548 49904
rect 19061 49855 19119 49861
rect 19720 49864 19932 49892
rect 21206 49864 21548 49892
rect 1765 49827 1823 49833
rect 1765 49793 1777 49827
rect 1811 49824 1823 49827
rect 4614 49824 4620 49836
rect 1811 49796 4620 49824
rect 1811 49793 1823 49796
rect 1765 49787 1823 49793
rect 4614 49784 4620 49796
rect 4672 49784 4678 49836
rect 11974 49784 11980 49836
rect 12032 49784 12038 49836
rect 13449 49827 13507 49833
rect 13449 49793 13461 49827
rect 13495 49824 13507 49827
rect 13495 49796 14044 49824
rect 13495 49793 13507 49796
rect 13449 49787 13507 49793
rect 1302 49716 1308 49768
rect 1360 49756 1366 49768
rect 2041 49759 2099 49765
rect 2041 49756 2053 49759
rect 1360 49728 2053 49756
rect 1360 49716 1366 49728
rect 2041 49725 2053 49728
rect 2087 49725 2099 49759
rect 2041 49719 2099 49725
rect 5350 49716 5356 49768
rect 5408 49756 5414 49768
rect 12897 49759 12955 49765
rect 12897 49756 12909 49759
rect 5408 49728 12909 49756
rect 5408 49716 5414 49728
rect 12897 49725 12909 49728
rect 12943 49725 12955 49759
rect 12897 49719 12955 49725
rect 14016 49688 14044 49796
rect 15654 49784 15660 49836
rect 15712 49824 15718 49836
rect 17497 49827 17555 49833
rect 17497 49824 17509 49827
rect 15712 49796 17509 49824
rect 15712 49784 15718 49796
rect 17497 49793 17509 49796
rect 17543 49824 17555 49827
rect 17586 49824 17592 49836
rect 17543 49796 17592 49824
rect 17543 49793 17555 49796
rect 17497 49787 17555 49793
rect 17586 49784 17592 49796
rect 17644 49784 17650 49836
rect 18322 49784 18328 49836
rect 18380 49824 18386 49836
rect 19720 49833 19748 49864
rect 21542 49852 21548 49864
rect 21600 49852 21606 49904
rect 22005 49895 22063 49901
rect 22005 49892 22017 49895
rect 21652 49864 22017 49892
rect 19705 49827 19763 49833
rect 18380 49796 19334 49824
rect 18380 49784 18386 49796
rect 14090 49716 14096 49768
rect 14148 49716 14154 49768
rect 14200 49728 15700 49756
rect 14200 49688 14228 49728
rect 15672 49700 15700 49728
rect 16022 49716 16028 49768
rect 16080 49756 16086 49768
rect 17681 49759 17739 49765
rect 17681 49756 17693 49759
rect 16080 49728 17693 49756
rect 16080 49716 16086 49728
rect 17681 49725 17693 49728
rect 17727 49725 17739 49759
rect 19306 49756 19334 49796
rect 19705 49793 19717 49827
rect 19751 49793 19763 49827
rect 21652 49824 21680 49864
rect 22005 49861 22017 49864
rect 22051 49861 22063 49895
rect 22005 49855 22063 49861
rect 22833 49895 22891 49901
rect 22833 49861 22845 49895
rect 22879 49892 22891 49895
rect 22879 49864 31754 49892
rect 22879 49861 22891 49864
rect 22833 49855 22891 49861
rect 22848 49824 22876 49855
rect 19705 49787 19763 49793
rect 21192 49796 21680 49824
rect 21744 49796 22876 49824
rect 23753 49827 23811 49833
rect 21192 49756 21220 49796
rect 19306 49728 21220 49756
rect 17681 49719 17739 49725
rect 21450 49716 21456 49768
rect 21508 49716 21514 49768
rect 14016 49660 14228 49688
rect 15654 49648 15660 49700
rect 15712 49648 15718 49700
rect 20990 49648 20996 49700
rect 21048 49688 21054 49700
rect 21744 49688 21772 49796
rect 23753 49793 23765 49827
rect 23799 49824 23811 49827
rect 24854 49824 24860 49836
rect 23799 49796 24860 49824
rect 23799 49793 23811 49796
rect 23753 49787 23811 49793
rect 24854 49784 24860 49796
rect 24912 49784 24918 49836
rect 21818 49716 21824 49768
rect 21876 49756 21882 49768
rect 23937 49759 23995 49765
rect 21876 49728 23796 49756
rect 21876 49716 21882 49728
rect 23768 49688 23796 49728
rect 23937 49725 23949 49759
rect 23983 49725 23995 49759
rect 31726 49756 31754 49864
rect 37550 49756 37556 49768
rect 31726 49728 37556 49756
rect 23937 49719 23995 49725
rect 23952 49688 23980 49719
rect 37550 49716 37556 49728
rect 37608 49716 37614 49768
rect 21048 49660 21772 49688
rect 22066 49660 23520 49688
rect 23768 49660 23980 49688
rect 21048 49648 21054 49660
rect 21468 49632 21496 49660
rect 14356 49623 14414 49629
rect 14356 49589 14368 49623
rect 14402 49620 14414 49623
rect 16390 49620 16396 49632
rect 14402 49592 16396 49620
rect 14402 49589 14414 49592
rect 14356 49583 14414 49589
rect 16390 49580 16396 49592
rect 16448 49580 16454 49632
rect 19968 49623 20026 49629
rect 19968 49589 19980 49623
rect 20014 49620 20026 49623
rect 21082 49620 21088 49632
rect 20014 49592 21088 49620
rect 20014 49589 20026 49592
rect 19968 49583 20026 49589
rect 21082 49580 21088 49592
rect 21140 49580 21146 49632
rect 21450 49580 21456 49632
rect 21508 49580 21514 49632
rect 21542 49580 21548 49632
rect 21600 49620 21606 49632
rect 22066 49620 22094 49660
rect 21600 49592 22094 49620
rect 23492 49620 23520 49660
rect 27154 49620 27160 49632
rect 23492 49592 27160 49620
rect 21600 49580 21606 49592
rect 27154 49580 27160 49592
rect 27212 49580 27218 49632
rect 1104 49530 49864 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 32950 49530
rect 33002 49478 33014 49530
rect 33066 49478 33078 49530
rect 33130 49478 33142 49530
rect 33194 49478 33206 49530
rect 33258 49478 42950 49530
rect 43002 49478 43014 49530
rect 43066 49478 43078 49530
rect 43130 49478 43142 49530
rect 43194 49478 43206 49530
rect 43258 49478 49864 49530
rect 1104 49456 49864 49478
rect 9950 49376 9956 49428
rect 10008 49416 10014 49428
rect 12989 49419 13047 49425
rect 12989 49416 13001 49419
rect 10008 49388 13001 49416
rect 10008 49376 10014 49388
rect 12989 49385 13001 49388
rect 13035 49385 13047 49419
rect 15838 49416 15844 49428
rect 12989 49379 13047 49385
rect 13648 49388 15844 49416
rect 11790 49308 11796 49360
rect 11848 49308 11854 49360
rect 12529 49351 12587 49357
rect 12529 49317 12541 49351
rect 12575 49348 12587 49351
rect 12618 49348 12624 49360
rect 12575 49320 12624 49348
rect 12575 49317 12587 49320
rect 12529 49311 12587 49317
rect 12618 49308 12624 49320
rect 12676 49308 12682 49360
rect 1302 49240 1308 49292
rect 1360 49280 1366 49292
rect 2041 49283 2099 49289
rect 2041 49280 2053 49283
rect 1360 49252 2053 49280
rect 1360 49240 1366 49252
rect 2041 49249 2053 49252
rect 2087 49249 2099 49283
rect 2041 49243 2099 49249
rect 3602 49240 3608 49292
rect 3660 49280 3666 49292
rect 13648 49289 13676 49388
rect 15838 49376 15844 49388
rect 15896 49376 15902 49428
rect 16482 49376 16488 49428
rect 16540 49376 16546 49428
rect 18506 49416 18512 49428
rect 16776 49388 18512 49416
rect 13814 49308 13820 49360
rect 13872 49348 13878 49360
rect 15933 49351 15991 49357
rect 15933 49348 15945 49351
rect 13872 49320 15945 49348
rect 13872 49308 13878 49320
rect 15933 49317 15945 49320
rect 15979 49317 15991 49351
rect 16500 49348 16528 49376
rect 15933 49311 15991 49317
rect 16408 49320 16528 49348
rect 13633 49283 13691 49289
rect 3660 49252 13584 49280
rect 3660 49240 3666 49252
rect 1765 49215 1823 49221
rect 1765 49181 1777 49215
rect 1811 49212 1823 49215
rect 3418 49212 3424 49224
rect 1811 49184 3424 49212
rect 1811 49181 1823 49184
rect 1765 49175 1823 49181
rect 3418 49172 3424 49184
rect 3476 49172 3482 49224
rect 13354 49172 13360 49224
rect 13412 49172 13418 49224
rect 13556 49212 13584 49252
rect 13633 49249 13645 49283
rect 13679 49249 13691 49283
rect 14918 49280 14924 49292
rect 13633 49243 13691 49249
rect 14568 49252 14924 49280
rect 14568 49212 14596 49252
rect 14918 49240 14924 49252
rect 14976 49240 14982 49292
rect 15010 49240 15016 49292
rect 15068 49280 15074 49292
rect 16408 49289 16436 49320
rect 15289 49283 15347 49289
rect 15289 49280 15301 49283
rect 15068 49252 15301 49280
rect 15068 49240 15074 49252
rect 15289 49249 15301 49252
rect 15335 49249 15347 49283
rect 15289 49243 15347 49249
rect 16393 49283 16451 49289
rect 16393 49249 16405 49283
rect 16439 49249 16451 49283
rect 16393 49243 16451 49249
rect 16482 49240 16488 49292
rect 16540 49240 16546 49292
rect 13556 49184 14596 49212
rect 14642 49172 14648 49224
rect 14700 49212 14706 49224
rect 15105 49215 15163 49221
rect 15105 49212 15117 49215
rect 14700 49184 15117 49212
rect 14700 49172 14706 49184
rect 15105 49181 15117 49184
rect 15151 49181 15163 49215
rect 15105 49175 15163 49181
rect 15197 49215 15255 49221
rect 15197 49181 15209 49215
rect 15243 49212 15255 49215
rect 16776 49212 16804 49388
rect 18506 49376 18512 49388
rect 18564 49376 18570 49428
rect 21542 49376 21548 49428
rect 21600 49376 21606 49428
rect 21634 49376 21640 49428
rect 21692 49416 21698 49428
rect 21692 49388 23520 49416
rect 21692 49376 21698 49388
rect 18598 49308 18604 49360
rect 18656 49348 18662 49360
rect 19334 49348 19340 49360
rect 18656 49320 19340 49348
rect 18656 49308 18662 49320
rect 19334 49308 19340 49320
rect 19392 49308 19398 49360
rect 19702 49308 19708 49360
rect 19760 49308 19766 49360
rect 21560 49348 21588 49376
rect 20824 49320 21588 49348
rect 17034 49240 17040 49292
rect 17092 49280 17098 49292
rect 17129 49283 17187 49289
rect 17129 49280 17141 49283
rect 17092 49252 17141 49280
rect 17092 49240 17098 49252
rect 17129 49249 17141 49252
rect 17175 49249 17187 49283
rect 17129 49243 17187 49249
rect 17405 49283 17463 49289
rect 17405 49249 17417 49283
rect 17451 49280 17463 49283
rect 17770 49280 17776 49292
rect 17451 49252 17776 49280
rect 17451 49249 17463 49252
rect 17405 49243 17463 49249
rect 17770 49240 17776 49252
rect 17828 49240 17834 49292
rect 18874 49240 18880 49292
rect 18932 49240 18938 49292
rect 20824 49289 20852 49320
rect 20809 49283 20867 49289
rect 20809 49249 20821 49283
rect 20855 49249 20867 49283
rect 20809 49243 20867 49249
rect 20901 49283 20959 49289
rect 20901 49249 20913 49283
rect 20947 49249 20959 49283
rect 20901 49243 20959 49249
rect 15243 49184 16804 49212
rect 15243 49181 15255 49184
rect 15197 49175 15255 49181
rect 19058 49172 19064 49224
rect 19116 49212 19122 49224
rect 20916 49212 20944 49243
rect 21450 49240 21456 49292
rect 21508 49280 21514 49292
rect 21545 49283 21603 49289
rect 21545 49280 21557 49283
rect 21508 49252 21557 49280
rect 21508 49240 21514 49252
rect 21545 49249 21557 49252
rect 21591 49249 21603 49283
rect 21545 49243 21603 49249
rect 21821 49283 21879 49289
rect 21821 49249 21833 49283
rect 21867 49280 21879 49283
rect 22554 49280 22560 49292
rect 21867 49252 22560 49280
rect 21867 49249 21879 49252
rect 21821 49243 21879 49249
rect 22554 49240 22560 49252
rect 22612 49240 22618 49292
rect 23492 49280 23520 49388
rect 24949 49283 25007 49289
rect 24949 49280 24961 49283
rect 23492 49252 24961 49280
rect 24949 49249 24961 49252
rect 24995 49249 25007 49283
rect 24949 49243 25007 49249
rect 26050 49240 26056 49292
rect 26108 49240 26114 49292
rect 23382 49212 23388 49224
rect 19116 49184 20944 49212
rect 22954 49184 23388 49212
rect 19116 49172 19122 49184
rect 23382 49172 23388 49184
rect 23440 49172 23446 49224
rect 24857 49215 24915 49221
rect 24857 49181 24869 49215
rect 24903 49212 24915 49215
rect 30466 49212 30472 49224
rect 24903 49184 30472 49212
rect 24903 49181 24915 49184
rect 24857 49175 24915 49181
rect 30466 49172 30472 49184
rect 30524 49172 30530 49224
rect 9766 49104 9772 49156
rect 9824 49144 9830 49156
rect 11609 49147 11667 49153
rect 11609 49144 11621 49147
rect 9824 49116 11621 49144
rect 9824 49104 9830 49116
rect 11609 49113 11621 49116
rect 11655 49113 11667 49147
rect 11609 49107 11667 49113
rect 12345 49147 12403 49153
rect 12345 49113 12357 49147
rect 12391 49144 12403 49147
rect 12710 49144 12716 49156
rect 12391 49116 12716 49144
rect 12391 49113 12403 49116
rect 12345 49107 12403 49113
rect 12710 49104 12716 49116
rect 12768 49104 12774 49156
rect 13449 49147 13507 49153
rect 13449 49113 13461 49147
rect 13495 49144 13507 49147
rect 13495 49116 16436 49144
rect 13495 49113 13507 49116
rect 13449 49107 13507 49113
rect 13538 49036 13544 49088
rect 13596 49076 13602 49088
rect 14737 49079 14795 49085
rect 14737 49076 14749 49079
rect 13596 49048 14749 49076
rect 13596 49036 13602 49048
rect 14737 49045 14749 49048
rect 14783 49045 14795 49079
rect 14737 49039 14795 49045
rect 14918 49036 14924 49088
rect 14976 49076 14982 49088
rect 16114 49076 16120 49088
rect 14976 49048 16120 49076
rect 14976 49036 14982 49048
rect 16114 49036 16120 49048
rect 16172 49076 16178 49088
rect 16301 49079 16359 49085
rect 16301 49076 16313 49079
rect 16172 49048 16313 49076
rect 16172 49036 16178 49048
rect 16301 49045 16313 49048
rect 16347 49045 16359 49079
rect 16408 49076 16436 49116
rect 18414 49104 18420 49156
rect 18472 49104 18478 49156
rect 18690 49104 18696 49156
rect 18748 49144 18754 49156
rect 19521 49147 19579 49153
rect 19521 49144 19533 49147
rect 18748 49116 19533 49144
rect 18748 49104 18754 49116
rect 19521 49113 19533 49116
rect 19567 49113 19579 49147
rect 19521 49107 19579 49113
rect 20717 49147 20775 49153
rect 20717 49113 20729 49147
rect 20763 49144 20775 49147
rect 20763 49116 22094 49144
rect 20763 49113 20775 49116
rect 20717 49107 20775 49113
rect 17494 49076 17500 49088
rect 16408 49048 17500 49076
rect 16301 49039 16359 49045
rect 17494 49036 17500 49048
rect 17552 49036 17558 49088
rect 17770 49036 17776 49088
rect 17828 49076 17834 49088
rect 20349 49079 20407 49085
rect 20349 49076 20361 49079
rect 17828 49048 20361 49076
rect 17828 49036 17834 49048
rect 20349 49045 20361 49048
rect 20395 49045 20407 49079
rect 22066 49076 22094 49116
rect 23198 49104 23204 49156
rect 23256 49144 23262 49156
rect 23256 49116 24440 49144
rect 23256 49104 23262 49116
rect 22186 49076 22192 49088
rect 22066 49048 22192 49076
rect 20349 49039 20407 49045
rect 22186 49036 22192 49048
rect 22244 49036 22250 49088
rect 22554 49036 22560 49088
rect 22612 49076 22618 49088
rect 24412 49085 24440 49116
rect 24762 49104 24768 49156
rect 24820 49144 24826 49156
rect 24820 49116 25912 49144
rect 24820 49104 24826 49116
rect 25884 49088 25912 49116
rect 23293 49079 23351 49085
rect 23293 49076 23305 49079
rect 22612 49048 23305 49076
rect 22612 49036 22618 49048
rect 23293 49045 23305 49048
rect 23339 49045 23351 49079
rect 23293 49039 23351 49045
rect 24397 49079 24455 49085
rect 24397 49045 24409 49079
rect 24443 49045 24455 49079
rect 24397 49039 24455 49045
rect 25498 49036 25504 49088
rect 25556 49036 25562 49088
rect 25866 49036 25872 49088
rect 25924 49036 25930 49088
rect 25961 49079 26019 49085
rect 25961 49045 25973 49079
rect 26007 49076 26019 49079
rect 33778 49076 33784 49088
rect 26007 49048 33784 49076
rect 26007 49045 26019 49048
rect 25961 49039 26019 49045
rect 33778 49036 33784 49048
rect 33836 49036 33842 49088
rect 1104 48986 49864 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 27950 48986
rect 28002 48934 28014 48986
rect 28066 48934 28078 48986
rect 28130 48934 28142 48986
rect 28194 48934 28206 48986
rect 28258 48934 37950 48986
rect 38002 48934 38014 48986
rect 38066 48934 38078 48986
rect 38130 48934 38142 48986
rect 38194 48934 38206 48986
rect 38258 48934 47950 48986
rect 48002 48934 48014 48986
rect 48066 48934 48078 48986
rect 48130 48934 48142 48986
rect 48194 48934 48206 48986
rect 48258 48934 49864 48986
rect 1104 48912 49864 48934
rect 9214 48832 9220 48884
rect 9272 48872 9278 48884
rect 9585 48875 9643 48881
rect 9585 48872 9597 48875
rect 9272 48844 9597 48872
rect 9272 48832 9278 48844
rect 9585 48841 9597 48844
rect 9631 48841 9643 48875
rect 14090 48872 14096 48884
rect 9585 48835 9643 48841
rect 13004 48844 14096 48872
rect 9769 48739 9827 48745
rect 9769 48705 9781 48739
rect 9815 48736 9827 48739
rect 11238 48736 11244 48748
rect 9815 48708 11244 48736
rect 9815 48705 9827 48708
rect 9769 48699 9827 48705
rect 11238 48696 11244 48708
rect 11296 48696 11302 48748
rect 13004 48745 13032 48844
rect 14090 48832 14096 48844
rect 14148 48832 14154 48884
rect 15933 48875 15991 48881
rect 15933 48841 15945 48875
rect 15979 48872 15991 48875
rect 16298 48872 16304 48884
rect 15979 48844 16304 48872
rect 15979 48841 15991 48844
rect 15933 48835 15991 48841
rect 16298 48832 16304 48844
rect 16356 48832 16362 48884
rect 17773 48875 17831 48881
rect 17773 48841 17785 48875
rect 17819 48872 17831 48875
rect 17819 48844 19564 48872
rect 17819 48841 17831 48844
rect 17773 48835 17831 48841
rect 14734 48804 14740 48816
rect 14490 48776 14740 48804
rect 14734 48764 14740 48776
rect 14792 48764 14798 48816
rect 16025 48807 16083 48813
rect 16025 48773 16037 48807
rect 16071 48804 16083 48807
rect 18598 48804 18604 48816
rect 16071 48776 18604 48804
rect 16071 48773 16083 48776
rect 16025 48767 16083 48773
rect 18598 48764 18604 48776
rect 18656 48764 18662 48816
rect 19536 48804 19564 48844
rect 19886 48832 19892 48884
rect 19944 48872 19950 48884
rect 20165 48875 20223 48881
rect 20165 48872 20177 48875
rect 19944 48844 20177 48872
rect 19944 48832 19950 48844
rect 20165 48841 20177 48844
rect 20211 48841 20223 48875
rect 20165 48835 20223 48841
rect 21082 48832 21088 48884
rect 21140 48872 21146 48884
rect 23290 48872 23296 48884
rect 21140 48844 23296 48872
rect 21140 48832 21146 48844
rect 23290 48832 23296 48844
rect 23348 48872 23354 48884
rect 23753 48875 23811 48881
rect 23753 48872 23765 48875
rect 23348 48844 23765 48872
rect 23348 48832 23354 48844
rect 23753 48841 23765 48844
rect 23799 48841 23811 48875
rect 23753 48835 23811 48841
rect 25041 48875 25099 48881
rect 25041 48841 25053 48875
rect 25087 48872 25099 48875
rect 25961 48875 26019 48881
rect 25961 48872 25973 48875
rect 25087 48844 25973 48872
rect 25087 48841 25099 48844
rect 25041 48835 25099 48841
rect 25961 48841 25973 48844
rect 26007 48872 26019 48875
rect 28902 48872 28908 48884
rect 26007 48844 28908 48872
rect 26007 48841 26019 48844
rect 25961 48835 26019 48841
rect 28902 48832 28908 48844
rect 28960 48832 28966 48884
rect 21266 48804 21272 48816
rect 19168 48776 19380 48804
rect 19536 48776 21272 48804
rect 12989 48739 13047 48745
rect 12989 48705 13001 48739
rect 13035 48705 13047 48739
rect 12989 48699 13047 48705
rect 16114 48696 16120 48748
rect 16172 48736 16178 48748
rect 17681 48739 17739 48745
rect 17681 48736 17693 48739
rect 16172 48708 17693 48736
rect 16172 48696 16178 48708
rect 17681 48705 17693 48708
rect 17727 48736 17739 48739
rect 17727 48708 18460 48736
rect 17727 48705 17739 48708
rect 17681 48699 17739 48705
rect 13265 48671 13323 48677
rect 13265 48637 13277 48671
rect 13311 48668 13323 48671
rect 15010 48668 15016 48680
rect 13311 48640 15016 48668
rect 13311 48637 13323 48640
rect 13265 48631 13323 48637
rect 15010 48628 15016 48640
rect 15068 48628 15074 48680
rect 16206 48628 16212 48680
rect 16264 48628 16270 48680
rect 17865 48671 17923 48677
rect 17865 48637 17877 48671
rect 17911 48637 17923 48671
rect 18432 48668 18460 48708
rect 18506 48696 18512 48748
rect 18564 48736 18570 48748
rect 19168 48736 19196 48776
rect 18564 48708 19196 48736
rect 19245 48739 19303 48745
rect 18564 48696 18570 48708
rect 19245 48705 19257 48739
rect 19291 48705 19303 48739
rect 19352 48736 19380 48776
rect 21266 48764 21272 48776
rect 21324 48764 21330 48816
rect 21450 48764 21456 48816
rect 21508 48764 21514 48816
rect 20349 48739 20407 48745
rect 20349 48736 20361 48739
rect 19352 48708 20361 48736
rect 19245 48699 19303 48705
rect 20349 48705 20361 48708
rect 20395 48705 20407 48739
rect 21468 48736 21496 48764
rect 21910 48736 21916 48748
rect 21468 48708 21916 48736
rect 20349 48699 20407 48705
rect 19150 48668 19156 48680
rect 18432 48640 19156 48668
rect 17865 48631 17923 48637
rect 16666 48560 16672 48612
rect 16724 48600 16730 48612
rect 16724 48572 17448 48600
rect 16724 48560 16730 48572
rect 12529 48535 12587 48541
rect 12529 48501 12541 48535
rect 12575 48532 12587 48535
rect 13354 48532 13360 48544
rect 12575 48504 13360 48532
rect 12575 48501 12587 48504
rect 12529 48495 12587 48501
rect 13354 48492 13360 48504
rect 13412 48492 13418 48544
rect 14642 48492 14648 48544
rect 14700 48532 14706 48544
rect 14737 48535 14795 48541
rect 14737 48532 14749 48535
rect 14700 48504 14749 48532
rect 14700 48492 14706 48504
rect 14737 48501 14749 48504
rect 14783 48501 14795 48535
rect 14737 48495 14795 48501
rect 15194 48492 15200 48544
rect 15252 48532 15258 48544
rect 15565 48535 15623 48541
rect 15565 48532 15577 48535
rect 15252 48504 15577 48532
rect 15252 48492 15258 48504
rect 15565 48501 15577 48504
rect 15611 48501 15623 48535
rect 15565 48495 15623 48501
rect 17310 48492 17316 48544
rect 17368 48492 17374 48544
rect 17420 48532 17448 48572
rect 17494 48560 17500 48612
rect 17552 48600 17558 48612
rect 17880 48600 17908 48631
rect 19150 48628 19156 48640
rect 19208 48628 19214 48680
rect 17552 48572 17908 48600
rect 17552 48560 17558 48572
rect 18877 48535 18935 48541
rect 18877 48532 18889 48535
rect 17420 48504 18889 48532
rect 18877 48501 18889 48504
rect 18923 48501 18935 48535
rect 19260 48532 19288 48699
rect 21910 48696 21916 48708
rect 21968 48736 21974 48748
rect 22005 48739 22063 48745
rect 22005 48736 22017 48739
rect 21968 48708 22017 48736
rect 21968 48696 21974 48708
rect 22005 48705 22017 48708
rect 22051 48705 22063 48739
rect 22005 48699 22063 48705
rect 23382 48696 23388 48748
rect 23440 48696 23446 48748
rect 24854 48696 24860 48748
rect 24912 48736 24918 48748
rect 25869 48739 25927 48745
rect 25869 48736 25881 48739
rect 24912 48708 25881 48736
rect 24912 48696 24918 48708
rect 25869 48705 25881 48708
rect 25915 48736 25927 48739
rect 30742 48736 30748 48748
rect 25915 48708 30748 48736
rect 25915 48705 25927 48708
rect 25869 48699 25927 48705
rect 30742 48696 30748 48708
rect 30800 48696 30806 48748
rect 19337 48671 19395 48677
rect 19337 48637 19349 48671
rect 19383 48637 19395 48671
rect 19337 48631 19395 48637
rect 19521 48671 19579 48677
rect 19521 48637 19533 48671
rect 19567 48668 19579 48671
rect 20254 48668 20260 48680
rect 19567 48640 20260 48668
rect 19567 48637 19579 48640
rect 19521 48631 19579 48637
rect 19352 48600 19380 48631
rect 20254 48628 20260 48640
rect 20312 48628 20318 48680
rect 21450 48628 21456 48680
rect 21508 48668 21514 48680
rect 22281 48671 22339 48677
rect 22281 48668 22293 48671
rect 21508 48640 22293 48668
rect 21508 48628 21514 48640
rect 22281 48637 22293 48640
rect 22327 48637 22339 48671
rect 22281 48631 22339 48637
rect 22370 48628 22376 48680
rect 22428 48668 22434 48680
rect 23658 48668 23664 48680
rect 22428 48640 23664 48668
rect 22428 48628 22434 48640
rect 23658 48628 23664 48640
rect 23716 48628 23722 48680
rect 24762 48628 24768 48680
rect 24820 48668 24826 48680
rect 26053 48671 26111 48677
rect 26053 48668 26065 48671
rect 24820 48640 26065 48668
rect 24820 48628 24826 48640
rect 26053 48637 26065 48640
rect 26099 48637 26111 48671
rect 26053 48631 26111 48637
rect 19352 48572 22094 48600
rect 20714 48532 20720 48544
rect 19260 48504 20720 48532
rect 18877 48495 18935 48501
rect 20714 48492 20720 48504
rect 20772 48492 20778 48544
rect 20990 48492 20996 48544
rect 21048 48492 21054 48544
rect 22066 48532 22094 48572
rect 22462 48532 22468 48544
rect 22066 48504 22468 48532
rect 22462 48492 22468 48504
rect 22520 48492 22526 48544
rect 24946 48492 24952 48544
rect 25004 48532 25010 48544
rect 25501 48535 25559 48541
rect 25501 48532 25513 48535
rect 25004 48504 25513 48532
rect 25004 48492 25010 48504
rect 25501 48501 25513 48504
rect 25547 48501 25559 48535
rect 25501 48495 25559 48501
rect 1104 48442 49864 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 32950 48442
rect 33002 48390 33014 48442
rect 33066 48390 33078 48442
rect 33130 48390 33142 48442
rect 33194 48390 33206 48442
rect 33258 48390 42950 48442
rect 43002 48390 43014 48442
rect 43066 48390 43078 48442
rect 43130 48390 43142 48442
rect 43194 48390 43206 48442
rect 43258 48390 49864 48442
rect 1104 48368 49864 48390
rect 12710 48288 12716 48340
rect 12768 48328 12774 48340
rect 13262 48328 13268 48340
rect 12768 48300 13268 48328
rect 12768 48288 12774 48300
rect 13262 48288 13268 48300
rect 13320 48288 13326 48340
rect 16390 48288 16396 48340
rect 16448 48288 16454 48340
rect 19426 48288 19432 48340
rect 19484 48328 19490 48340
rect 25498 48328 25504 48340
rect 19484 48300 25504 48328
rect 19484 48288 19490 48300
rect 25498 48288 25504 48300
rect 25556 48288 25562 48340
rect 24029 48263 24087 48269
rect 20272 48232 22416 48260
rect 1302 48152 1308 48204
rect 1360 48192 1366 48204
rect 2041 48195 2099 48201
rect 2041 48192 2053 48195
rect 1360 48164 2053 48192
rect 1360 48152 1366 48164
rect 2041 48161 2053 48164
rect 2087 48161 2099 48195
rect 2041 48155 2099 48161
rect 13630 48152 13636 48204
rect 13688 48152 13694 48204
rect 14090 48152 14096 48204
rect 14148 48192 14154 48204
rect 14645 48195 14703 48201
rect 14645 48192 14657 48195
rect 14148 48164 14657 48192
rect 14148 48152 14154 48164
rect 14645 48161 14657 48164
rect 14691 48161 14703 48195
rect 14645 48155 14703 48161
rect 17034 48152 17040 48204
rect 17092 48192 17098 48204
rect 17129 48195 17187 48201
rect 17129 48192 17141 48195
rect 17092 48164 17141 48192
rect 17092 48152 17098 48164
rect 17129 48161 17141 48164
rect 17175 48161 17187 48195
rect 17129 48155 17187 48161
rect 17402 48152 17408 48204
rect 17460 48192 17466 48204
rect 18874 48192 18880 48204
rect 17460 48164 18880 48192
rect 17460 48152 17466 48164
rect 18874 48152 18880 48164
rect 18932 48152 18938 48204
rect 20272 48201 20300 48232
rect 20257 48195 20315 48201
rect 20257 48161 20269 48195
rect 20303 48161 20315 48195
rect 20257 48155 20315 48161
rect 20530 48152 20536 48204
rect 20588 48192 20594 48204
rect 20588 48164 21404 48192
rect 20588 48152 20594 48164
rect 1765 48127 1823 48133
rect 1765 48093 1777 48127
rect 1811 48124 1823 48127
rect 3878 48124 3884 48136
rect 1811 48096 3884 48124
rect 1811 48093 1823 48096
rect 1765 48087 1823 48093
rect 3878 48084 3884 48096
rect 3936 48084 3942 48136
rect 12526 48084 12532 48136
rect 12584 48084 12590 48136
rect 13354 48084 13360 48136
rect 13412 48084 13418 48136
rect 13449 48127 13507 48133
rect 13449 48093 13461 48127
rect 13495 48124 13507 48127
rect 13814 48124 13820 48136
rect 13495 48096 13820 48124
rect 13495 48093 13507 48096
rect 13449 48087 13507 48093
rect 13814 48084 13820 48096
rect 13872 48084 13878 48136
rect 19981 48127 20039 48133
rect 19981 48093 19993 48127
rect 20027 48124 20039 48127
rect 20990 48124 20996 48136
rect 20027 48096 20996 48124
rect 20027 48093 20039 48096
rect 19981 48087 20039 48093
rect 20990 48084 20996 48096
rect 21048 48084 21054 48136
rect 21266 48084 21272 48136
rect 21324 48084 21330 48136
rect 21376 48124 21404 48164
rect 21910 48152 21916 48204
rect 21968 48192 21974 48204
rect 22388 48192 22416 48232
rect 24029 48229 24041 48263
rect 24075 48260 24087 48263
rect 24854 48260 24860 48272
rect 24075 48232 24860 48260
rect 24075 48229 24087 48232
rect 24029 48223 24087 48229
rect 24854 48220 24860 48232
rect 24912 48260 24918 48272
rect 26050 48260 26056 48272
rect 24912 48232 26056 48260
rect 24912 48220 24918 48232
rect 26050 48220 26056 48232
rect 26108 48220 26114 48272
rect 22554 48192 22560 48204
rect 21968 48164 22324 48192
rect 22388 48164 22560 48192
rect 21968 48152 21974 48164
rect 22296 48136 22324 48164
rect 22554 48152 22560 48164
rect 22612 48152 22618 48204
rect 26329 48195 26387 48201
rect 26329 48192 26341 48195
rect 24136 48164 26341 48192
rect 21376 48096 22094 48124
rect 14918 48016 14924 48068
rect 14976 48016 14982 48068
rect 16206 48056 16212 48068
rect 16146 48028 16212 48056
rect 16206 48016 16212 48028
rect 16264 48056 16270 48068
rect 17862 48056 17868 48068
rect 16264 48028 17868 48056
rect 16264 48016 16270 48028
rect 17862 48016 17868 48028
rect 17920 48016 17926 48068
rect 20073 48059 20131 48065
rect 18708 48028 19656 48056
rect 12618 47948 12624 48000
rect 12676 47988 12682 48000
rect 12989 47991 13047 47997
rect 12989 47988 13001 47991
rect 12676 47960 13001 47988
rect 12676 47948 12682 47960
rect 12989 47957 13001 47960
rect 13035 47957 13047 47991
rect 12989 47951 13047 47957
rect 16758 47948 16764 48000
rect 16816 47988 16822 48000
rect 18708 47988 18736 48028
rect 16816 47960 18736 47988
rect 18877 47991 18935 47997
rect 16816 47948 16822 47960
rect 18877 47957 18889 47991
rect 18923 47988 18935 47991
rect 18966 47988 18972 48000
rect 18923 47960 18972 47988
rect 18923 47957 18935 47960
rect 18877 47951 18935 47957
rect 18966 47948 18972 47960
rect 19024 47948 19030 48000
rect 19628 47997 19656 48028
rect 20073 48025 20085 48059
rect 20119 48056 20131 48059
rect 21726 48056 21732 48068
rect 20119 48028 21732 48056
rect 20119 48025 20131 48028
rect 20073 48019 20131 48025
rect 21726 48016 21732 48028
rect 21784 48016 21790 48068
rect 19613 47991 19671 47997
rect 19613 47957 19625 47991
rect 19659 47957 19671 47991
rect 19613 47951 19671 47957
rect 21085 47991 21143 47997
rect 21085 47957 21097 47991
rect 21131 47988 21143 47991
rect 21174 47988 21180 48000
rect 21131 47960 21180 47988
rect 21131 47957 21143 47960
rect 21085 47951 21143 47957
rect 21174 47948 21180 47960
rect 21232 47948 21238 48000
rect 22066 47988 22094 48096
rect 22278 48084 22284 48136
rect 22336 48084 22342 48136
rect 24136 48124 24164 48164
rect 26329 48161 26341 48164
rect 26375 48161 26387 48195
rect 26329 48155 26387 48161
rect 23860 48096 24164 48124
rect 23566 48016 23572 48068
rect 23624 48016 23630 48068
rect 23860 47988 23888 48096
rect 25866 48084 25872 48136
rect 25924 48124 25930 48136
rect 26145 48127 26203 48133
rect 26145 48124 26157 48127
rect 25924 48096 26157 48124
rect 25924 48084 25930 48096
rect 26145 48093 26157 48096
rect 26191 48124 26203 48127
rect 32858 48124 32864 48136
rect 26191 48096 32864 48124
rect 26191 48093 26203 48096
rect 26145 48087 26203 48093
rect 32858 48084 32864 48096
rect 32916 48084 32922 48136
rect 25317 48059 25375 48065
rect 25317 48025 25329 48059
rect 25363 48056 25375 48059
rect 26237 48059 26295 48065
rect 26237 48056 26249 48059
rect 25363 48028 26249 48056
rect 25363 48025 25375 48028
rect 25317 48019 25375 48025
rect 26237 48025 26249 48028
rect 26283 48056 26295 48059
rect 26283 48028 35894 48056
rect 26283 48025 26295 48028
rect 26237 48019 26295 48025
rect 22066 47960 23888 47988
rect 25774 47948 25780 48000
rect 25832 47948 25838 48000
rect 35866 47988 35894 48028
rect 48958 48016 48964 48068
rect 49016 48016 49022 48068
rect 40034 47988 40040 48000
rect 35866 47960 40040 47988
rect 40034 47948 40040 47960
rect 40092 47948 40098 48000
rect 49050 47948 49056 48000
rect 49108 47948 49114 48000
rect 1104 47898 49864 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 27950 47898
rect 28002 47846 28014 47898
rect 28066 47846 28078 47898
rect 28130 47846 28142 47898
rect 28194 47846 28206 47898
rect 28258 47846 37950 47898
rect 38002 47846 38014 47898
rect 38066 47846 38078 47898
rect 38130 47846 38142 47898
rect 38194 47846 38206 47898
rect 38258 47846 47950 47898
rect 48002 47846 48014 47898
rect 48066 47846 48078 47898
rect 48130 47846 48142 47898
rect 48194 47846 48206 47898
rect 48258 47846 49864 47898
rect 1104 47824 49864 47846
rect 9677 47787 9735 47793
rect 9677 47753 9689 47787
rect 9723 47784 9735 47787
rect 9858 47784 9864 47796
rect 9723 47756 9864 47784
rect 9723 47753 9735 47756
rect 9677 47747 9735 47753
rect 9858 47744 9864 47756
rect 9916 47744 9922 47796
rect 10321 47787 10379 47793
rect 10321 47753 10333 47787
rect 10367 47784 10379 47787
rect 10502 47784 10508 47796
rect 10367 47756 10508 47784
rect 10367 47753 10379 47756
rect 10321 47747 10379 47753
rect 10502 47744 10508 47756
rect 10560 47744 10566 47796
rect 10686 47744 10692 47796
rect 10744 47784 10750 47796
rect 11701 47787 11759 47793
rect 11701 47784 11713 47787
rect 10744 47756 11713 47784
rect 10744 47744 10750 47756
rect 11701 47753 11713 47756
rect 11747 47753 11759 47787
rect 11701 47747 11759 47753
rect 12526 47744 12532 47796
rect 12584 47784 12590 47796
rect 15933 47787 15991 47793
rect 15933 47784 15945 47787
rect 12584 47756 15945 47784
rect 12584 47744 12590 47756
rect 15933 47753 15945 47756
rect 15979 47753 15991 47787
rect 15933 47747 15991 47753
rect 16025 47787 16083 47793
rect 16025 47753 16037 47787
rect 16071 47784 16083 47787
rect 19518 47784 19524 47796
rect 16071 47756 19524 47784
rect 16071 47753 16083 47756
rect 16025 47747 16083 47753
rect 19518 47744 19524 47756
rect 19576 47744 19582 47796
rect 22278 47784 22284 47796
rect 19720 47756 22284 47784
rect 11606 47716 11612 47728
rect 10520 47688 11612 47716
rect 1765 47651 1823 47657
rect 1765 47617 1777 47651
rect 1811 47648 1823 47651
rect 4154 47648 4160 47660
rect 1811 47620 4160 47648
rect 1811 47617 1823 47620
rect 1765 47611 1823 47617
rect 4154 47608 4160 47620
rect 4212 47608 4218 47660
rect 9858 47608 9864 47660
rect 9916 47608 9922 47660
rect 10520 47657 10548 47688
rect 11606 47676 11612 47688
rect 11664 47676 11670 47728
rect 13722 47716 13728 47728
rect 12406 47688 13728 47716
rect 10505 47651 10563 47657
rect 10505 47617 10517 47651
rect 10551 47617 10563 47651
rect 10505 47611 10563 47617
rect 11149 47651 11207 47657
rect 11149 47617 11161 47651
rect 11195 47617 11207 47651
rect 11149 47611 11207 47617
rect 11885 47651 11943 47657
rect 11885 47617 11897 47651
rect 11931 47648 11943 47651
rect 12406 47648 12434 47688
rect 13722 47676 13728 47688
rect 13780 47676 13786 47728
rect 16206 47716 16212 47728
rect 14858 47688 16212 47716
rect 11931 47620 12434 47648
rect 11931 47617 11943 47620
rect 11885 47611 11943 47617
rect 1302 47540 1308 47592
rect 1360 47580 1366 47592
rect 2041 47583 2099 47589
rect 2041 47580 2053 47583
rect 1360 47552 2053 47580
rect 1360 47540 1366 47552
rect 2041 47549 2053 47552
rect 2087 47549 2099 47583
rect 11164 47580 11192 47611
rect 14734 47608 14740 47660
rect 14792 47608 14798 47660
rect 12526 47580 12532 47592
rect 11164 47552 12532 47580
rect 2041 47543 2099 47549
rect 12526 47540 12532 47552
rect 12584 47540 12590 47592
rect 13357 47583 13415 47589
rect 13357 47549 13369 47583
rect 13403 47549 13415 47583
rect 13357 47543 13415 47549
rect 8386 47472 8392 47524
rect 8444 47512 8450 47524
rect 10965 47515 11023 47521
rect 10965 47512 10977 47515
rect 8444 47484 10977 47512
rect 8444 47472 8450 47484
rect 10965 47481 10977 47484
rect 11011 47481 11023 47515
rect 10965 47475 11023 47481
rect 13372 47444 13400 47543
rect 13630 47540 13636 47592
rect 13688 47540 13694 47592
rect 13998 47540 14004 47592
rect 14056 47580 14062 47592
rect 14752 47580 14780 47608
rect 14936 47580 14964 47688
rect 16206 47676 16212 47688
rect 16264 47676 16270 47728
rect 17402 47676 17408 47728
rect 17460 47676 17466 47728
rect 17954 47676 17960 47728
rect 18012 47716 18018 47728
rect 18012 47688 18170 47716
rect 18012 47676 18018 47688
rect 17420 47648 17448 47676
rect 19720 47657 19748 47756
rect 22278 47744 22284 47756
rect 22336 47784 22342 47796
rect 25317 47787 25375 47793
rect 22336 47756 23060 47784
rect 22336 47744 22342 47756
rect 16224 47620 17448 47648
rect 19705 47651 19763 47657
rect 14056 47552 14688 47580
rect 14752 47552 14964 47580
rect 14056 47540 14062 47552
rect 14660 47512 14688 47552
rect 15010 47540 15016 47592
rect 15068 47580 15074 47592
rect 16224 47589 16252 47620
rect 19705 47617 19717 47651
rect 19751 47617 19763 47651
rect 19705 47611 19763 47617
rect 20990 47608 20996 47660
rect 21048 47648 21054 47660
rect 23032 47657 23060 47756
rect 25317 47753 25329 47787
rect 25363 47784 25375 47787
rect 26237 47787 26295 47793
rect 26237 47784 26249 47787
rect 25363 47756 26249 47784
rect 25363 47753 25375 47756
rect 25317 47747 25375 47753
rect 26237 47753 26249 47756
rect 26283 47784 26295 47787
rect 30374 47784 30380 47796
rect 26283 47756 30380 47784
rect 26283 47753 26295 47756
rect 26237 47747 26295 47753
rect 30374 47744 30380 47756
rect 30432 47744 30438 47796
rect 48958 47744 48964 47796
rect 49016 47784 49022 47796
rect 49142 47784 49148 47796
rect 49016 47756 49148 47784
rect 49016 47744 49022 47756
rect 49142 47744 49148 47756
rect 49200 47744 49206 47796
rect 23566 47676 23572 47728
rect 23624 47716 23630 47728
rect 23624 47688 23782 47716
rect 23624 47676 23630 47688
rect 23017 47651 23075 47657
rect 21048 47620 21114 47648
rect 21048 47608 21054 47620
rect 23017 47617 23029 47651
rect 23063 47617 23075 47651
rect 23017 47611 23075 47617
rect 26142 47608 26148 47660
rect 26200 47608 26206 47660
rect 15105 47583 15163 47589
rect 15105 47580 15117 47583
rect 15068 47552 15117 47580
rect 15068 47540 15074 47552
rect 15105 47549 15117 47552
rect 15151 47549 15163 47583
rect 15105 47543 15163 47549
rect 16209 47583 16267 47589
rect 16209 47549 16221 47583
rect 16255 47549 16267 47583
rect 16209 47543 16267 47549
rect 17126 47540 17132 47592
rect 17184 47580 17190 47592
rect 17405 47583 17463 47589
rect 17405 47580 17417 47583
rect 17184 47552 17417 47580
rect 17184 47540 17190 47552
rect 17405 47549 17417 47552
rect 17451 47549 17463 47583
rect 17405 47543 17463 47549
rect 17681 47583 17739 47589
rect 17681 47549 17693 47583
rect 17727 47580 17739 47583
rect 18966 47580 18972 47592
rect 17727 47552 18972 47580
rect 17727 47549 17739 47552
rect 17681 47543 17739 47549
rect 18966 47540 18972 47552
rect 19024 47540 19030 47592
rect 19981 47583 20039 47589
rect 19981 47549 19993 47583
rect 20027 47580 20039 47583
rect 20622 47580 20628 47592
rect 20027 47552 20628 47580
rect 20027 47549 20039 47552
rect 19981 47543 20039 47549
rect 20622 47540 20628 47552
rect 20680 47540 20686 47592
rect 20714 47540 20720 47592
rect 20772 47580 20778 47592
rect 22189 47583 22247 47589
rect 22189 47580 22201 47583
rect 20772 47552 22201 47580
rect 20772 47540 20778 47552
rect 22189 47549 22201 47552
rect 22235 47549 22247 47583
rect 23293 47583 23351 47589
rect 23293 47580 23305 47583
rect 22189 47543 22247 47549
rect 23124 47552 23305 47580
rect 17310 47512 17316 47524
rect 14660 47484 17316 47512
rect 17310 47472 17316 47484
rect 17368 47472 17374 47524
rect 23124 47512 23152 47552
rect 23293 47549 23305 47552
rect 23339 47580 23351 47583
rect 24026 47580 24032 47592
rect 23339 47552 24032 47580
rect 23339 47549 23351 47552
rect 23293 47543 23351 47549
rect 24026 47540 24032 47552
rect 24084 47540 24090 47592
rect 24762 47540 24768 47592
rect 24820 47540 24826 47592
rect 26329 47583 26387 47589
rect 26329 47549 26341 47583
rect 26375 47549 26387 47583
rect 26329 47543 26387 47549
rect 21008 47484 23152 47512
rect 14274 47444 14280 47456
rect 13372 47416 14280 47444
rect 14274 47404 14280 47416
rect 14332 47404 14338 47456
rect 14734 47404 14740 47456
rect 14792 47444 14798 47456
rect 15565 47447 15623 47453
rect 15565 47444 15577 47447
rect 14792 47416 15577 47444
rect 14792 47404 14798 47416
rect 15565 47413 15577 47416
rect 15611 47413 15623 47447
rect 15565 47407 15623 47413
rect 17402 47404 17408 47456
rect 17460 47444 17466 47456
rect 19153 47447 19211 47453
rect 19153 47444 19165 47447
rect 17460 47416 19165 47444
rect 17460 47404 17466 47416
rect 19153 47413 19165 47416
rect 19199 47413 19211 47447
rect 19153 47407 19211 47413
rect 19242 47404 19248 47456
rect 19300 47444 19306 47456
rect 21008 47444 21036 47484
rect 24302 47472 24308 47524
rect 24360 47512 24366 47524
rect 26344 47512 26372 47543
rect 24360 47484 26372 47512
rect 24360 47472 24366 47484
rect 19300 47416 21036 47444
rect 19300 47404 19306 47416
rect 21450 47404 21456 47456
rect 21508 47404 21514 47456
rect 22462 47404 22468 47456
rect 22520 47444 22526 47456
rect 25777 47447 25835 47453
rect 25777 47444 25789 47447
rect 22520 47416 25789 47444
rect 22520 47404 22526 47416
rect 25777 47413 25789 47416
rect 25823 47413 25835 47447
rect 25777 47407 25835 47413
rect 1104 47354 49864 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 32950 47354
rect 33002 47302 33014 47354
rect 33066 47302 33078 47354
rect 33130 47302 33142 47354
rect 33194 47302 33206 47354
rect 33258 47302 42950 47354
rect 43002 47302 43014 47354
rect 43066 47302 43078 47354
rect 43130 47302 43142 47354
rect 43194 47302 43206 47354
rect 43258 47302 49864 47354
rect 1104 47280 49864 47302
rect 10778 47200 10784 47252
rect 10836 47240 10842 47252
rect 11149 47243 11207 47249
rect 11149 47240 11161 47243
rect 10836 47212 11161 47240
rect 10836 47200 10842 47212
rect 11149 47209 11161 47212
rect 11195 47209 11207 47243
rect 13538 47240 13544 47252
rect 11149 47203 11207 47209
rect 12406 47212 13544 47240
rect 8754 47132 8760 47184
rect 8812 47172 8818 47184
rect 11793 47175 11851 47181
rect 11793 47172 11805 47175
rect 8812 47144 11805 47172
rect 8812 47132 8818 47144
rect 11793 47141 11805 47144
rect 11839 47141 11851 47175
rect 12406 47172 12434 47212
rect 13538 47200 13544 47212
rect 13596 47200 13602 47252
rect 16298 47240 16304 47252
rect 14200 47212 16304 47240
rect 11793 47135 11851 47141
rect 12268 47144 12434 47172
rect 12268 47113 12296 47144
rect 12710 47132 12716 47184
rect 12768 47172 12774 47184
rect 12989 47175 13047 47181
rect 12989 47172 13001 47175
rect 12768 47144 13001 47172
rect 12768 47132 12774 47144
rect 12989 47141 13001 47144
rect 13035 47141 13047 47175
rect 13906 47172 13912 47184
rect 12989 47135 13047 47141
rect 13372 47144 13912 47172
rect 12253 47107 12311 47113
rect 12253 47073 12265 47107
rect 12299 47073 12311 47107
rect 12253 47067 12311 47073
rect 12345 47107 12403 47113
rect 12345 47073 12357 47107
rect 12391 47104 12403 47107
rect 13372 47104 13400 47144
rect 13906 47132 13912 47144
rect 13964 47132 13970 47184
rect 12391 47076 13400 47104
rect 12391 47073 12403 47076
rect 12345 47067 12403 47073
rect 13630 47064 13636 47116
rect 13688 47104 13694 47116
rect 14200 47104 14228 47212
rect 16298 47200 16304 47212
rect 16356 47200 16362 47252
rect 18877 47243 18935 47249
rect 18877 47209 18889 47243
rect 18923 47240 18935 47243
rect 19058 47240 19064 47252
rect 18923 47212 19064 47240
rect 18923 47209 18935 47212
rect 18877 47203 18935 47209
rect 19058 47200 19064 47212
rect 19116 47200 19122 47252
rect 21361 47243 21419 47249
rect 21361 47209 21373 47243
rect 21407 47240 21419 47243
rect 21634 47240 21640 47252
rect 21407 47212 21640 47240
rect 21407 47209 21419 47212
rect 21361 47203 21419 47209
rect 21634 47200 21640 47212
rect 21692 47200 21698 47252
rect 24026 47200 24032 47252
rect 24084 47200 24090 47252
rect 16022 47132 16028 47184
rect 16080 47132 16086 47184
rect 16390 47132 16396 47184
rect 16448 47172 16454 47184
rect 16448 47144 17264 47172
rect 16448 47132 16454 47144
rect 13688 47076 14228 47104
rect 13688 47064 13694 47076
rect 14274 47064 14280 47116
rect 14332 47104 14338 47116
rect 14550 47104 14556 47116
rect 14332 47076 14556 47104
rect 14332 47064 14338 47076
rect 14550 47064 14556 47076
rect 14608 47104 14614 47116
rect 17129 47107 17187 47113
rect 17129 47104 17141 47107
rect 14608 47076 17141 47104
rect 14608 47064 14614 47076
rect 17129 47073 17141 47076
rect 17175 47073 17187 47107
rect 17236 47104 17264 47144
rect 17402 47104 17408 47116
rect 17236 47076 17408 47104
rect 17129 47067 17187 47073
rect 17402 47064 17408 47076
rect 17460 47064 17466 47116
rect 22557 47107 22615 47113
rect 22557 47073 22569 47107
rect 22603 47104 22615 47107
rect 24854 47104 24860 47116
rect 22603 47076 24860 47104
rect 22603 47073 22615 47076
rect 22557 47067 22615 47073
rect 24854 47064 24860 47076
rect 24912 47064 24918 47116
rect 11333 47039 11391 47045
rect 11333 47005 11345 47039
rect 11379 47036 11391 47039
rect 12434 47036 12440 47048
rect 11379 47008 12440 47036
rect 11379 47005 11391 47008
rect 11333 46999 11391 47005
rect 12434 46996 12440 47008
rect 12492 46996 12498 47048
rect 12526 46996 12532 47048
rect 12584 47036 12590 47048
rect 13449 47039 13507 47045
rect 12584 47008 13400 47036
rect 12584 46996 12590 47008
rect 12161 46971 12219 46977
rect 12161 46937 12173 46971
rect 12207 46968 12219 46971
rect 12894 46968 12900 46980
rect 12207 46940 12900 46968
rect 12207 46937 12219 46940
rect 12161 46931 12219 46937
rect 12894 46928 12900 46940
rect 12952 46928 12958 46980
rect 13372 46968 13400 47008
rect 13449 47005 13461 47039
rect 13495 47036 13507 47039
rect 13998 47036 14004 47048
rect 13495 47008 14004 47036
rect 13495 47005 13507 47008
rect 13449 46999 13507 47005
rect 13998 46996 14004 47008
rect 14056 46996 14062 47048
rect 16022 46996 16028 47048
rect 16080 47036 16086 47048
rect 16669 47039 16727 47045
rect 16669 47036 16681 47039
rect 16080 47008 16681 47036
rect 16080 46996 16086 47008
rect 16669 47005 16681 47008
rect 16715 47005 16727 47039
rect 16669 46999 16727 47005
rect 19610 46996 19616 47048
rect 19668 46996 19674 47048
rect 22278 46996 22284 47048
rect 22336 46996 22342 47048
rect 13372 46940 13492 46968
rect 13354 46860 13360 46912
rect 13412 46860 13418 46912
rect 13464 46900 13492 46940
rect 13906 46928 13912 46980
rect 13964 46968 13970 46980
rect 14553 46971 14611 46977
rect 14553 46968 14565 46971
rect 13964 46940 14565 46968
rect 13964 46928 13970 46940
rect 14553 46937 14565 46940
rect 14599 46968 14611 46971
rect 14642 46968 14648 46980
rect 14599 46940 14648 46968
rect 14599 46937 14611 46940
rect 14553 46931 14611 46937
rect 14642 46928 14648 46940
rect 14700 46928 14706 46980
rect 16206 46968 16212 46980
rect 15778 46940 16212 46968
rect 16206 46928 16212 46940
rect 16264 46968 16270 46980
rect 17862 46968 17868 46980
rect 16264 46940 17868 46968
rect 16264 46928 16270 46940
rect 17862 46928 17868 46940
rect 17920 46928 17926 46980
rect 19242 46928 19248 46980
rect 19300 46968 19306 46980
rect 19889 46971 19947 46977
rect 19889 46968 19901 46971
rect 19300 46940 19901 46968
rect 19300 46928 19306 46940
rect 19889 46937 19901 46940
rect 19935 46937 19947 46971
rect 19889 46931 19947 46937
rect 20898 46928 20904 46980
rect 20956 46928 20962 46980
rect 23566 46928 23572 46980
rect 23624 46928 23630 46980
rect 13538 46900 13544 46912
rect 13464 46872 13544 46900
rect 13538 46860 13544 46872
rect 13596 46860 13602 46912
rect 18322 46860 18328 46912
rect 18380 46900 18386 46912
rect 18782 46900 18788 46912
rect 18380 46872 18788 46900
rect 18380 46860 18386 46872
rect 18782 46860 18788 46872
rect 18840 46860 18846 46912
rect 1104 46810 49864 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 27950 46810
rect 28002 46758 28014 46810
rect 28066 46758 28078 46810
rect 28130 46758 28142 46810
rect 28194 46758 28206 46810
rect 28258 46758 37950 46810
rect 38002 46758 38014 46810
rect 38066 46758 38078 46810
rect 38130 46758 38142 46810
rect 38194 46758 38206 46810
rect 38258 46758 47950 46810
rect 48002 46758 48014 46810
rect 48066 46758 48078 46810
rect 48130 46758 48142 46810
rect 48194 46758 48206 46810
rect 48258 46758 49864 46810
rect 1104 46736 49864 46758
rect 2314 46656 2320 46708
rect 2372 46696 2378 46708
rect 4249 46699 4307 46705
rect 4249 46696 4261 46699
rect 2372 46668 4261 46696
rect 2372 46656 2378 46668
rect 4249 46665 4261 46668
rect 4295 46665 4307 46699
rect 4249 46659 4307 46665
rect 5166 46656 5172 46708
rect 5224 46656 5230 46708
rect 10962 46656 10968 46708
rect 11020 46656 11026 46708
rect 13817 46699 13875 46705
rect 13817 46665 13829 46699
rect 13863 46696 13875 46699
rect 13863 46668 16160 46696
rect 13863 46665 13875 46668
rect 13817 46659 13875 46665
rect 16132 46628 16160 46668
rect 16298 46656 16304 46708
rect 16356 46656 16362 46708
rect 19702 46696 19708 46708
rect 17512 46668 19708 46696
rect 16574 46628 16580 46640
rect 16132 46600 16580 46628
rect 16574 46588 16580 46600
rect 16632 46588 16638 46640
rect 1765 46563 1823 46569
rect 1765 46529 1777 46563
rect 1811 46560 1823 46563
rect 4157 46563 4215 46569
rect 1811 46532 2774 46560
rect 1811 46529 1823 46532
rect 1765 46523 1823 46529
rect 1302 46452 1308 46504
rect 1360 46492 1366 46504
rect 2041 46495 2099 46501
rect 2041 46492 2053 46495
rect 1360 46464 2053 46492
rect 1360 46452 1366 46464
rect 2041 46461 2053 46464
rect 2087 46461 2099 46495
rect 2746 46492 2774 46532
rect 4157 46529 4169 46563
rect 4203 46560 4215 46563
rect 4522 46560 4528 46572
rect 4203 46532 4528 46560
rect 4203 46529 4215 46532
rect 4157 46523 4215 46529
rect 4522 46520 4528 46532
rect 4580 46520 4586 46572
rect 5077 46563 5135 46569
rect 5077 46529 5089 46563
rect 5123 46560 5135 46563
rect 9582 46560 9588 46572
rect 5123 46532 9588 46560
rect 5123 46529 5135 46532
rect 5077 46523 5135 46529
rect 9582 46520 9588 46532
rect 9640 46520 9646 46572
rect 11149 46563 11207 46569
rect 11149 46529 11161 46563
rect 11195 46560 11207 46563
rect 12526 46560 12532 46572
rect 11195 46532 12532 46560
rect 11195 46529 11207 46532
rect 11149 46523 11207 46529
rect 12526 46520 12532 46532
rect 12584 46520 12590 46572
rect 12894 46520 12900 46572
rect 12952 46520 12958 46572
rect 13725 46563 13783 46569
rect 13725 46529 13737 46563
rect 13771 46560 13783 46563
rect 14458 46560 14464 46572
rect 13771 46532 14464 46560
rect 13771 46529 13783 46532
rect 13725 46523 13783 46529
rect 14458 46520 14464 46532
rect 14516 46520 14522 46572
rect 16206 46560 16212 46572
rect 15962 46532 16212 46560
rect 16206 46520 16212 46532
rect 16264 46520 16270 46572
rect 17126 46520 17132 46572
rect 17184 46560 17190 46572
rect 17512 46569 17540 46668
rect 19702 46656 19708 46668
rect 19760 46656 19766 46708
rect 20806 46656 20812 46708
rect 20864 46696 20870 46708
rect 21453 46699 21511 46705
rect 21453 46696 21465 46699
rect 20864 46668 21465 46696
rect 20864 46656 20870 46668
rect 21453 46665 21465 46668
rect 21499 46696 21511 46699
rect 21818 46696 21824 46708
rect 21499 46668 21824 46696
rect 21499 46665 21511 46668
rect 21453 46659 21511 46665
rect 21818 46656 21824 46668
rect 21876 46656 21882 46708
rect 23566 46656 23572 46708
rect 23624 46696 23630 46708
rect 24121 46699 24179 46705
rect 23624 46668 23796 46696
rect 23624 46656 23630 46668
rect 17862 46588 17868 46640
rect 17920 46628 17926 46640
rect 17920 46600 18262 46628
rect 17920 46588 17926 46600
rect 20714 46588 20720 46640
rect 20772 46588 20778 46640
rect 17497 46563 17555 46569
rect 17497 46560 17509 46563
rect 17184 46532 17509 46560
rect 17184 46520 17190 46532
rect 17497 46529 17509 46532
rect 17543 46529 17555 46563
rect 23768 46546 23796 46668
rect 24121 46665 24133 46699
rect 24167 46696 24179 46699
rect 24302 46696 24308 46708
rect 24167 46668 24308 46696
rect 24167 46665 24179 46668
rect 24121 46659 24179 46665
rect 24302 46656 24308 46668
rect 24360 46656 24366 46708
rect 17497 46523 17555 46529
rect 25406 46520 25412 46572
rect 25464 46560 25470 46572
rect 25501 46563 25559 46569
rect 25501 46560 25513 46563
rect 25464 46532 25513 46560
rect 25464 46520 25470 46532
rect 25501 46529 25513 46532
rect 25547 46529 25559 46563
rect 25501 46523 25559 46529
rect 25593 46563 25651 46569
rect 25593 46529 25605 46563
rect 25639 46560 25651 46563
rect 33502 46560 33508 46572
rect 25639 46532 33508 46560
rect 25639 46529 25651 46532
rect 25593 46523 25651 46529
rect 4430 46492 4436 46504
rect 2746 46464 4436 46492
rect 2041 46455 2099 46461
rect 4430 46452 4436 46464
rect 4488 46452 4494 46504
rect 13998 46452 14004 46504
rect 14056 46452 14062 46504
rect 14550 46452 14556 46504
rect 14608 46452 14614 46504
rect 14829 46495 14887 46501
rect 14829 46461 14841 46495
rect 14875 46492 14887 46495
rect 17402 46492 17408 46504
rect 14875 46464 17408 46492
rect 14875 46461 14887 46464
rect 14829 46455 14887 46461
rect 17402 46452 17408 46464
rect 17460 46452 17466 46504
rect 17773 46495 17831 46501
rect 17773 46461 17785 46495
rect 17819 46492 17831 46495
rect 19058 46492 19064 46504
rect 17819 46464 19064 46492
rect 17819 46461 17831 46464
rect 17773 46455 17831 46461
rect 19058 46452 19064 46464
rect 19116 46452 19122 46504
rect 19702 46452 19708 46504
rect 19760 46452 19766 46504
rect 19978 46452 19984 46504
rect 20036 46452 20042 46504
rect 22278 46452 22284 46504
rect 22336 46492 22342 46504
rect 22373 46495 22431 46501
rect 22373 46492 22385 46495
rect 22336 46464 22385 46492
rect 22336 46452 22342 46464
rect 22373 46461 22385 46464
rect 22419 46461 22431 46495
rect 22373 46455 22431 46461
rect 22646 46452 22652 46504
rect 22704 46452 22710 46504
rect 24673 46495 24731 46501
rect 24673 46461 24685 46495
rect 24719 46492 24731 46495
rect 25608 46492 25636 46523
rect 33502 46520 33508 46532
rect 33560 46520 33566 46572
rect 24719 46464 25636 46492
rect 25685 46495 25743 46501
rect 24719 46461 24731 46464
rect 24673 46455 24731 46461
rect 25685 46461 25697 46495
rect 25731 46461 25743 46495
rect 25685 46455 25743 46461
rect 11330 46384 11336 46436
rect 11388 46424 11394 46436
rect 13357 46427 13415 46433
rect 13357 46424 13369 46427
rect 11388 46396 13369 46424
rect 11388 46384 11394 46396
rect 13357 46393 13369 46396
rect 13403 46393 13415 46427
rect 13357 46387 13415 46393
rect 24026 46384 24032 46436
rect 24084 46424 24090 46436
rect 25700 46424 25728 46455
rect 24084 46396 25728 46424
rect 24084 46384 24090 46396
rect 17034 46316 17040 46368
rect 17092 46316 17098 46368
rect 18414 46316 18420 46368
rect 18472 46356 18478 46368
rect 19242 46356 19248 46368
rect 18472 46328 19248 46356
rect 18472 46316 18478 46328
rect 19242 46316 19248 46328
rect 19300 46316 19306 46368
rect 25130 46316 25136 46368
rect 25188 46316 25194 46368
rect 1104 46266 49864 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 32950 46266
rect 33002 46214 33014 46266
rect 33066 46214 33078 46266
rect 33130 46214 33142 46266
rect 33194 46214 33206 46266
rect 33258 46214 42950 46266
rect 43002 46214 43014 46266
rect 43066 46214 43078 46266
rect 43130 46214 43142 46266
rect 43194 46214 43206 46266
rect 43258 46214 49864 46266
rect 1104 46192 49864 46214
rect 3326 46112 3332 46164
rect 3384 46152 3390 46164
rect 4157 46155 4215 46161
rect 4157 46152 4169 46155
rect 3384 46124 4169 46152
rect 3384 46112 3390 46124
rect 4157 46121 4169 46124
rect 4203 46121 4215 46155
rect 4157 46115 4215 46121
rect 7834 46112 7840 46164
rect 7892 46152 7898 46164
rect 8021 46155 8079 46161
rect 8021 46152 8033 46155
rect 7892 46124 8033 46152
rect 7892 46112 7898 46124
rect 8021 46121 8033 46124
rect 8067 46121 8079 46155
rect 8021 46115 8079 46121
rect 11054 46112 11060 46164
rect 11112 46152 11118 46164
rect 11241 46155 11299 46161
rect 11241 46152 11253 46155
rect 11112 46124 11253 46152
rect 11112 46112 11118 46124
rect 11241 46121 11253 46124
rect 11287 46121 11299 46155
rect 11241 46115 11299 46121
rect 13354 46112 13360 46164
rect 13412 46152 13418 46164
rect 13725 46155 13783 46161
rect 13725 46152 13737 46155
rect 13412 46124 13737 46152
rect 13412 46112 13418 46124
rect 13725 46121 13737 46124
rect 13771 46121 13783 46155
rect 13725 46115 13783 46121
rect 13998 46112 14004 46164
rect 14056 46152 14062 46164
rect 14918 46152 14924 46164
rect 14056 46124 14924 46152
rect 14056 46112 14062 46124
rect 14918 46112 14924 46124
rect 14976 46152 14982 46164
rect 16301 46155 16359 46161
rect 16301 46152 16313 46155
rect 14976 46124 16313 46152
rect 14976 46112 14982 46124
rect 16301 46121 16313 46124
rect 16347 46121 16359 46155
rect 16301 46115 16359 46121
rect 17402 46112 17408 46164
rect 17460 46152 17466 46164
rect 18877 46155 18935 46161
rect 18877 46152 18889 46155
rect 17460 46124 18889 46152
rect 17460 46112 17466 46124
rect 18877 46121 18889 46124
rect 18923 46121 18935 46155
rect 18877 46115 18935 46121
rect 20336 46155 20394 46161
rect 20336 46121 20348 46155
rect 20382 46152 20394 46155
rect 21634 46152 21640 46164
rect 20382 46124 21640 46152
rect 20382 46121 20394 46124
rect 20336 46115 20394 46121
rect 21634 46112 21640 46124
rect 21692 46112 21698 46164
rect 1302 45976 1308 46028
rect 1360 46016 1366 46028
rect 2041 46019 2099 46025
rect 2041 46016 2053 46019
rect 1360 45988 2053 46016
rect 1360 45976 1366 45988
rect 2041 45985 2053 45988
rect 2087 45985 2099 46019
rect 2041 45979 2099 45985
rect 14829 46019 14887 46025
rect 14829 45985 14841 46019
rect 14875 46016 14887 46019
rect 16114 46016 16120 46028
rect 14875 45988 16120 46016
rect 14875 45985 14887 45988
rect 14829 45979 14887 45985
rect 16114 45976 16120 45988
rect 16172 45976 16178 46028
rect 17126 45976 17132 46028
rect 17184 45976 17190 46028
rect 17405 46019 17463 46025
rect 17405 45985 17417 46019
rect 17451 46016 17463 46019
rect 19518 46016 19524 46028
rect 17451 45988 19524 46016
rect 17451 45985 17463 45988
rect 17405 45979 17463 45985
rect 19518 45976 19524 45988
rect 19576 45976 19582 46028
rect 19702 45976 19708 46028
rect 19760 46016 19766 46028
rect 20073 46019 20131 46025
rect 20073 46016 20085 46019
rect 19760 45988 20085 46016
rect 19760 45976 19766 45988
rect 20073 45985 20085 45988
rect 20119 46016 20131 46019
rect 20346 46016 20352 46028
rect 20119 45988 20352 46016
rect 20119 45985 20131 45988
rect 20073 45979 20131 45985
rect 20346 45976 20352 45988
rect 20404 45976 20410 46028
rect 22557 46019 22615 46025
rect 22557 45985 22569 46019
rect 22603 46016 22615 46019
rect 24762 46016 24768 46028
rect 22603 45988 24768 46016
rect 22603 45985 22615 45988
rect 22557 45979 22615 45985
rect 24762 45976 24768 45988
rect 24820 45976 24826 46028
rect 1765 45951 1823 45957
rect 1765 45917 1777 45951
rect 1811 45948 1823 45951
rect 3694 45948 3700 45960
rect 1811 45920 3700 45948
rect 1811 45917 1823 45920
rect 1765 45911 1823 45917
rect 3694 45908 3700 45920
rect 3752 45908 3758 45960
rect 7742 45908 7748 45960
rect 7800 45948 7806 45960
rect 8205 45951 8263 45957
rect 8205 45948 8217 45951
rect 7800 45920 8217 45948
rect 7800 45908 7806 45920
rect 8205 45917 8217 45920
rect 8251 45917 8263 45951
rect 8205 45911 8263 45917
rect 11422 45908 11428 45960
rect 11480 45908 11486 45960
rect 14550 45908 14556 45960
rect 14608 45908 14614 45960
rect 19334 45908 19340 45960
rect 19392 45948 19398 45960
rect 19613 45951 19671 45957
rect 19613 45948 19625 45951
rect 19392 45920 19625 45948
rect 19392 45908 19398 45920
rect 19613 45917 19625 45920
rect 19659 45917 19671 45951
rect 19613 45911 19671 45917
rect 22278 45908 22284 45960
rect 22336 45908 22342 45960
rect 47854 45908 47860 45960
rect 47912 45948 47918 45960
rect 47949 45951 48007 45957
rect 47949 45948 47961 45951
rect 47912 45920 47961 45948
rect 47912 45908 47918 45920
rect 47949 45917 47961 45920
rect 47995 45917 48007 45951
rect 47949 45911 48007 45917
rect 49142 45908 49148 45960
rect 49200 45908 49206 45960
rect 4065 45883 4123 45889
rect 4065 45849 4077 45883
rect 4111 45880 4123 45883
rect 5442 45880 5448 45892
rect 4111 45852 5448 45880
rect 4111 45849 4123 45852
rect 4065 45843 4123 45849
rect 5442 45840 5448 45852
rect 5500 45840 5506 45892
rect 14568 45880 14596 45908
rect 16206 45880 16212 45892
rect 14568 45852 14688 45880
rect 16054 45852 16212 45880
rect 14660 45812 14688 45852
rect 16206 45840 16212 45852
rect 16264 45880 16270 45892
rect 17862 45880 17868 45892
rect 16264 45852 17868 45880
rect 16264 45840 16270 45852
rect 17862 45840 17868 45852
rect 17920 45840 17926 45892
rect 20806 45840 20812 45892
rect 20864 45840 20870 45892
rect 23566 45840 23572 45892
rect 23624 45840 23630 45892
rect 15102 45812 15108 45824
rect 14660 45784 15108 45812
rect 15102 45772 15108 45784
rect 15160 45772 15166 45824
rect 19978 45772 19984 45824
rect 20036 45812 20042 45824
rect 21821 45815 21879 45821
rect 21821 45812 21833 45815
rect 20036 45784 21833 45812
rect 20036 45772 20042 45784
rect 21821 45781 21833 45784
rect 21867 45781 21879 45815
rect 21821 45775 21879 45781
rect 22646 45772 22652 45824
rect 22704 45812 22710 45824
rect 24029 45815 24087 45821
rect 24029 45812 24041 45815
rect 22704 45784 24041 45812
rect 22704 45772 22710 45784
rect 24029 45781 24041 45784
rect 24075 45781 24087 45815
rect 24029 45775 24087 45781
rect 1104 45722 49864 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 27950 45722
rect 28002 45670 28014 45722
rect 28066 45670 28078 45722
rect 28130 45670 28142 45722
rect 28194 45670 28206 45722
rect 28258 45670 37950 45722
rect 38002 45670 38014 45722
rect 38066 45670 38078 45722
rect 38130 45670 38142 45722
rect 38194 45670 38206 45722
rect 38258 45670 47950 45722
rect 48002 45670 48014 45722
rect 48066 45670 48078 45722
rect 48130 45670 48142 45722
rect 48194 45670 48206 45722
rect 48258 45670 49864 45722
rect 1104 45648 49864 45670
rect 19337 45611 19395 45617
rect 15856 45580 16160 45608
rect 2682 45500 2688 45552
rect 2740 45500 2746 45552
rect 3878 45500 3884 45552
rect 3936 45500 3942 45552
rect 4614 45500 4620 45552
rect 4672 45500 4678 45552
rect 12618 45540 12624 45552
rect 9232 45512 12624 45540
rect 2498 45432 2504 45484
rect 2556 45432 2562 45484
rect 3697 45475 3755 45481
rect 3697 45441 3709 45475
rect 3743 45441 3755 45475
rect 3697 45435 3755 45441
rect 4433 45475 4491 45481
rect 4433 45441 4445 45475
rect 4479 45472 4491 45475
rect 5718 45472 5724 45484
rect 4479 45444 5724 45472
rect 4479 45441 4491 45444
rect 4433 45435 4491 45441
rect 3712 45404 3740 45435
rect 5718 45432 5724 45444
rect 5776 45472 5782 45484
rect 6822 45472 6828 45484
rect 5776 45444 6828 45472
rect 5776 45432 5782 45444
rect 6822 45432 6828 45444
rect 6880 45432 6886 45484
rect 8113 45475 8171 45481
rect 8113 45441 8125 45475
rect 8159 45472 8171 45475
rect 9122 45472 9128 45484
rect 8159 45444 9128 45472
rect 8159 45441 8171 45444
rect 8113 45435 8171 45441
rect 9122 45432 9128 45444
rect 9180 45432 9186 45484
rect 9232 45481 9260 45512
rect 12618 45500 12624 45512
rect 12676 45500 12682 45552
rect 15856 45540 15884 45580
rect 12728 45512 15884 45540
rect 15933 45543 15991 45549
rect 12728 45481 12756 45512
rect 15933 45509 15945 45543
rect 15979 45540 15991 45543
rect 16022 45540 16028 45552
rect 15979 45512 16028 45540
rect 15979 45509 15991 45512
rect 15933 45503 15991 45509
rect 16022 45500 16028 45512
rect 16080 45500 16086 45552
rect 16132 45540 16160 45580
rect 19337 45577 19349 45611
rect 19383 45608 19395 45611
rect 19426 45608 19432 45620
rect 19383 45580 19432 45608
rect 19383 45577 19395 45580
rect 19337 45571 19395 45577
rect 19426 45568 19432 45580
rect 19484 45568 19490 45620
rect 23750 45568 23756 45620
rect 23808 45608 23814 45620
rect 25406 45608 25412 45620
rect 23808 45580 25412 45608
rect 23808 45568 23814 45580
rect 25406 45568 25412 45580
rect 25464 45568 25470 45620
rect 16666 45540 16672 45552
rect 16132 45512 16672 45540
rect 16666 45500 16672 45512
rect 16724 45500 16730 45552
rect 18782 45540 18788 45552
rect 17420 45512 18788 45540
rect 17420 45484 17448 45512
rect 18782 45500 18788 45512
rect 18840 45540 18846 45552
rect 20073 45543 20131 45549
rect 20073 45540 20085 45543
rect 18840 45512 20085 45540
rect 18840 45500 18846 45512
rect 20073 45509 20085 45512
rect 20119 45509 20131 45543
rect 20073 45503 20131 45509
rect 23566 45500 23572 45552
rect 23624 45500 23630 45552
rect 9217 45475 9275 45481
rect 9217 45441 9229 45475
rect 9263 45441 9275 45475
rect 9217 45435 9275 45441
rect 11885 45475 11943 45481
rect 11885 45441 11897 45475
rect 11931 45472 11943 45475
rect 12713 45475 12771 45481
rect 11931 45444 12434 45472
rect 11931 45441 11943 45444
rect 11885 45435 11943 45441
rect 6178 45404 6184 45416
rect 3712 45376 6184 45404
rect 6178 45364 6184 45376
rect 6236 45404 6242 45416
rect 12406 45404 12434 45444
rect 12713 45441 12725 45475
rect 12759 45441 12771 45475
rect 12713 45435 12771 45441
rect 14461 45475 14519 45481
rect 14461 45441 14473 45475
rect 14507 45472 14519 45475
rect 14642 45472 14648 45484
rect 14507 45444 14648 45472
rect 14507 45441 14519 45444
rect 14461 45435 14519 45441
rect 14642 45432 14648 45444
rect 14700 45432 14706 45484
rect 15105 45475 15163 45481
rect 15105 45441 15117 45475
rect 15151 45472 15163 45475
rect 16482 45472 16488 45484
rect 15151 45444 16488 45472
rect 15151 45441 15163 45444
rect 15105 45435 15163 45441
rect 16482 45432 16488 45444
rect 16540 45432 16546 45484
rect 17402 45432 17408 45484
rect 17460 45432 17466 45484
rect 19245 45475 19303 45481
rect 19245 45441 19257 45475
rect 19291 45472 19303 45475
rect 22189 45475 22247 45481
rect 22189 45472 22201 45475
rect 19291 45444 22201 45472
rect 19291 45441 19303 45444
rect 19245 45435 19303 45441
rect 22189 45441 22201 45444
rect 22235 45441 22247 45475
rect 22189 45435 22247 45441
rect 15194 45404 15200 45416
rect 6236 45376 9076 45404
rect 12406 45376 15200 45404
rect 6236 45364 6242 45376
rect 7650 45296 7656 45348
rect 7708 45336 7714 45348
rect 9048 45345 9076 45376
rect 15194 45364 15200 45376
rect 15252 45364 15258 45416
rect 15930 45364 15936 45416
rect 15988 45404 15994 45416
rect 16025 45407 16083 45413
rect 16025 45404 16037 45407
rect 15988 45376 16037 45404
rect 15988 45364 15994 45376
rect 16025 45373 16037 45376
rect 16071 45373 16083 45407
rect 16025 45367 16083 45373
rect 16114 45364 16120 45416
rect 16172 45364 16178 45416
rect 18233 45407 18291 45413
rect 18233 45373 18245 45407
rect 18279 45404 18291 45407
rect 18322 45404 18328 45416
rect 18279 45376 18328 45404
rect 18279 45373 18291 45376
rect 18233 45367 18291 45373
rect 18322 45364 18328 45376
rect 18380 45364 18386 45416
rect 19429 45407 19487 45413
rect 19429 45373 19441 45407
rect 19475 45373 19487 45407
rect 19429 45367 19487 45373
rect 7929 45339 7987 45345
rect 7929 45336 7941 45339
rect 7708 45308 7941 45336
rect 7708 45296 7714 45308
rect 7929 45305 7941 45308
rect 7975 45305 7987 45339
rect 7929 45299 7987 45305
rect 9033 45339 9091 45345
rect 9033 45305 9045 45339
rect 9079 45305 9091 45339
rect 9033 45299 9091 45305
rect 10870 45296 10876 45348
rect 10928 45336 10934 45348
rect 12529 45339 12587 45345
rect 12529 45336 12541 45339
rect 10928 45308 12541 45336
rect 10928 45296 10934 45308
rect 12529 45305 12541 45308
rect 12575 45305 12587 45339
rect 12529 45299 12587 45305
rect 14182 45296 14188 45348
rect 14240 45336 14246 45348
rect 14240 45308 14412 45336
rect 14240 45296 14246 45308
rect 7006 45228 7012 45280
rect 7064 45268 7070 45280
rect 11701 45271 11759 45277
rect 11701 45268 11713 45271
rect 7064 45240 11713 45268
rect 7064 45228 7070 45240
rect 11701 45237 11713 45240
rect 11747 45237 11759 45271
rect 11701 45231 11759 45237
rect 12802 45228 12808 45280
rect 12860 45268 12866 45280
rect 14277 45271 14335 45277
rect 14277 45268 14289 45271
rect 12860 45240 14289 45268
rect 12860 45228 12866 45240
rect 14277 45237 14289 45240
rect 14323 45237 14335 45271
rect 14384 45268 14412 45308
rect 14458 45296 14464 45348
rect 14516 45336 14522 45348
rect 15565 45339 15623 45345
rect 15565 45336 15577 45339
rect 14516 45308 15577 45336
rect 14516 45296 14522 45308
rect 15565 45305 15577 45308
rect 15611 45305 15623 45339
rect 15565 45299 15623 45305
rect 19150 45296 19156 45348
rect 19208 45336 19214 45348
rect 19444 45336 19472 45367
rect 20346 45364 20352 45416
rect 20404 45404 20410 45416
rect 20901 45407 20959 45413
rect 20901 45404 20913 45407
rect 20404 45376 20913 45404
rect 20404 45364 20410 45376
rect 20901 45373 20913 45376
rect 20947 45404 20959 45407
rect 22278 45404 22284 45416
rect 20947 45376 22284 45404
rect 20947 45373 20959 45376
rect 20901 45367 20959 45373
rect 22278 45364 22284 45376
rect 22336 45404 22342 45416
rect 22830 45404 22836 45416
rect 22336 45376 22836 45404
rect 22336 45364 22342 45376
rect 22830 45364 22836 45376
rect 22888 45364 22894 45416
rect 23109 45407 23167 45413
rect 23109 45373 23121 45407
rect 23155 45404 23167 45407
rect 24302 45404 24308 45416
rect 23155 45376 24308 45404
rect 23155 45373 23167 45376
rect 23109 45367 23167 45373
rect 24302 45364 24308 45376
rect 24360 45364 24366 45416
rect 21450 45336 21456 45348
rect 19208 45308 19472 45336
rect 20732 45308 21456 45336
rect 19208 45296 19214 45308
rect 14921 45271 14979 45277
rect 14921 45268 14933 45271
rect 14384 45240 14933 45268
rect 14277 45231 14335 45237
rect 14921 45237 14933 45240
rect 14967 45237 14979 45271
rect 14921 45231 14979 45237
rect 15010 45228 15016 45280
rect 15068 45268 15074 45280
rect 18877 45271 18935 45277
rect 18877 45268 18889 45271
rect 15068 45240 18889 45268
rect 15068 45228 15074 45240
rect 18877 45237 18889 45240
rect 18923 45237 18935 45271
rect 18877 45231 18935 45237
rect 19242 45228 19248 45280
rect 19300 45268 19306 45280
rect 20732 45268 20760 45308
rect 21450 45296 21456 45308
rect 21508 45296 21514 45348
rect 19300 45240 20760 45268
rect 19300 45228 19306 45240
rect 20806 45228 20812 45280
rect 20864 45268 20870 45280
rect 23566 45268 23572 45280
rect 20864 45240 23572 45268
rect 20864 45228 20870 45240
rect 23566 45228 23572 45240
rect 23624 45228 23630 45280
rect 24578 45228 24584 45280
rect 24636 45228 24642 45280
rect 1104 45178 49864 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 32950 45178
rect 33002 45126 33014 45178
rect 33066 45126 33078 45178
rect 33130 45126 33142 45178
rect 33194 45126 33206 45178
rect 33258 45126 42950 45178
rect 43002 45126 43014 45178
rect 43066 45126 43078 45178
rect 43130 45126 43142 45178
rect 43194 45126 43206 45178
rect 43258 45126 49864 45178
rect 1104 45104 49864 45126
rect 3418 45024 3424 45076
rect 3476 45064 3482 45076
rect 4157 45067 4215 45073
rect 4157 45064 4169 45067
rect 3476 45036 4169 45064
rect 3476 45024 3482 45036
rect 4157 45033 4169 45036
rect 4203 45033 4215 45067
rect 4157 45027 4215 45033
rect 4706 45024 4712 45076
rect 4764 45064 4770 45076
rect 4893 45067 4951 45073
rect 4893 45064 4905 45067
rect 4764 45036 4905 45064
rect 4764 45024 4770 45036
rect 4893 45033 4905 45036
rect 4939 45033 4951 45067
rect 4893 45027 4951 45033
rect 5442 45024 5448 45076
rect 5500 45064 5506 45076
rect 9125 45067 9183 45073
rect 9125 45064 9137 45067
rect 5500 45036 9137 45064
rect 5500 45024 5506 45036
rect 9125 45033 9137 45036
rect 9171 45033 9183 45067
rect 9125 45027 9183 45033
rect 11057 45067 11115 45073
rect 11057 45033 11069 45067
rect 11103 45064 11115 45067
rect 11882 45064 11888 45076
rect 11103 45036 11888 45064
rect 11103 45033 11115 45036
rect 11057 45027 11115 45033
rect 11882 45024 11888 45036
rect 11940 45024 11946 45076
rect 12434 45024 12440 45076
rect 12492 45064 12498 45076
rect 13630 45064 13636 45076
rect 12492 45036 13636 45064
rect 12492 45024 12498 45036
rect 13630 45024 13636 45036
rect 13688 45024 13694 45076
rect 14366 45024 14372 45076
rect 14424 45064 14430 45076
rect 15105 45067 15163 45073
rect 15105 45064 15117 45067
rect 14424 45036 15117 45064
rect 14424 45024 14430 45036
rect 15105 45033 15117 45036
rect 15151 45033 15163 45067
rect 16758 45064 16764 45076
rect 15105 45027 15163 45033
rect 15212 45036 16764 45064
rect 12710 44996 12716 45008
rect 9324 44968 12716 44996
rect 1302 44888 1308 44940
rect 1360 44928 1366 44940
rect 2041 44931 2099 44937
rect 2041 44928 2053 44931
rect 1360 44900 2053 44928
rect 1360 44888 1366 44900
rect 2041 44897 2053 44900
rect 2087 44897 2099 44931
rect 2041 44891 2099 44897
rect 1765 44863 1823 44869
rect 1765 44829 1777 44863
rect 1811 44860 1823 44863
rect 4338 44860 4344 44872
rect 1811 44832 4344 44860
rect 1811 44829 1823 44832
rect 1765 44823 1823 44829
rect 4338 44820 4344 44832
rect 4396 44820 4402 44872
rect 5810 44860 5816 44872
rect 4724 44832 5816 44860
rect 4065 44795 4123 44801
rect 4065 44761 4077 44795
rect 4111 44792 4123 44795
rect 4724 44792 4752 44832
rect 5810 44820 5816 44832
rect 5868 44820 5874 44872
rect 9324 44869 9352 44968
rect 12710 44956 12716 44968
rect 12768 44956 12774 45008
rect 13078 44956 13084 45008
rect 13136 44956 13142 45008
rect 14734 44928 14740 44940
rect 10612 44900 14740 44928
rect 9309 44863 9367 44869
rect 9309 44829 9321 44863
rect 9355 44829 9367 44863
rect 9309 44823 9367 44829
rect 9950 44820 9956 44872
rect 10008 44820 10014 44872
rect 10612 44869 10640 44900
rect 14734 44888 14740 44900
rect 14792 44888 14798 44940
rect 10597 44863 10655 44869
rect 10597 44829 10609 44863
rect 10643 44829 10655 44863
rect 10597 44823 10655 44829
rect 11241 44863 11299 44869
rect 11241 44829 11253 44863
rect 11287 44829 11299 44863
rect 11241 44823 11299 44829
rect 11885 44863 11943 44869
rect 11885 44829 11897 44863
rect 11931 44860 11943 44863
rect 12434 44860 12440 44872
rect 11931 44832 12440 44860
rect 11931 44829 11943 44832
rect 11885 44823 11943 44829
rect 4111 44764 4752 44792
rect 4801 44795 4859 44801
rect 4111 44761 4123 44764
rect 4065 44755 4123 44761
rect 4801 44761 4813 44795
rect 4847 44792 4859 44795
rect 4982 44792 4988 44804
rect 4847 44764 4988 44792
rect 4847 44761 4859 44764
rect 4801 44755 4859 44761
rect 4982 44752 4988 44764
rect 5040 44752 5046 44804
rect 5626 44752 5632 44804
rect 5684 44792 5690 44804
rect 5684 44764 10456 44792
rect 5684 44752 5690 44764
rect 5534 44684 5540 44736
rect 5592 44724 5598 44736
rect 6362 44724 6368 44736
rect 5592 44696 6368 44724
rect 5592 44684 5598 44696
rect 6362 44684 6368 44696
rect 6420 44724 6426 44736
rect 10428 44733 10456 44764
rect 9769 44727 9827 44733
rect 9769 44724 9781 44727
rect 6420 44696 9781 44724
rect 6420 44684 6426 44696
rect 9769 44693 9781 44696
rect 9815 44693 9827 44727
rect 9769 44687 9827 44693
rect 10413 44727 10471 44733
rect 10413 44693 10425 44727
rect 10459 44693 10471 44727
rect 11256 44724 11284 44823
rect 12434 44820 12440 44832
rect 12492 44820 12498 44872
rect 12526 44820 12532 44872
rect 12584 44820 12590 44872
rect 13265 44863 13323 44869
rect 13265 44829 13277 44863
rect 13311 44860 13323 44863
rect 13311 44832 14412 44860
rect 13311 44829 13323 44832
rect 13265 44823 13323 44829
rect 12342 44752 12348 44804
rect 12400 44792 12406 44804
rect 14384 44792 14412 44832
rect 14458 44820 14464 44872
rect 14516 44820 14522 44872
rect 15212 44792 15240 45036
rect 16758 45024 16764 45036
rect 16816 45024 16822 45076
rect 22738 45064 22744 45076
rect 18616 45036 22744 45064
rect 16850 44996 16856 45008
rect 16316 44968 16856 44996
rect 15289 44863 15347 44869
rect 15289 44829 15301 44863
rect 15335 44860 15347 44863
rect 16316 44860 16344 44968
rect 16850 44956 16856 44968
rect 16908 44956 16914 45008
rect 16945 44999 17003 45005
rect 16945 44965 16957 44999
rect 16991 44965 17003 44999
rect 16945 44959 17003 44965
rect 16390 44888 16396 44940
rect 16448 44888 16454 44940
rect 16960 44928 16988 44959
rect 17126 44956 17132 45008
rect 17184 44996 17190 45008
rect 18141 44999 18199 45005
rect 18141 44996 18153 44999
rect 17184 44968 18153 44996
rect 17184 44956 17190 44968
rect 18141 44965 18153 44968
rect 18187 44965 18199 44999
rect 18141 44959 18199 44965
rect 16500 44900 16988 44928
rect 17589 44931 17647 44937
rect 15335 44832 16344 44860
rect 15335 44829 15347 44832
rect 15289 44823 15347 44829
rect 12400 44764 14320 44792
rect 14384 44764 15240 44792
rect 12400 44752 12406 44764
rect 13446 44724 13452 44736
rect 11256 44696 13452 44724
rect 10413 44687 10471 44693
rect 13446 44684 13452 44696
rect 13504 44684 13510 44736
rect 14292 44733 14320 44764
rect 15378 44752 15384 44804
rect 15436 44792 15442 44804
rect 16500 44792 16528 44900
rect 17589 44897 17601 44931
rect 17635 44928 17647 44931
rect 18414 44928 18420 44940
rect 17635 44900 18420 44928
rect 17635 44897 17647 44900
rect 17589 44891 17647 44897
rect 18414 44888 18420 44900
rect 18472 44888 18478 44940
rect 18616 44937 18644 45036
rect 22738 45024 22744 45036
rect 22796 45024 22802 45076
rect 18601 44931 18659 44937
rect 18601 44897 18613 44931
rect 18647 44897 18659 44931
rect 18601 44891 18659 44897
rect 18785 44931 18843 44937
rect 18785 44897 18797 44931
rect 18831 44928 18843 44931
rect 19242 44928 19248 44940
rect 18831 44900 19248 44928
rect 18831 44897 18843 44900
rect 18785 44891 18843 44897
rect 19242 44888 19248 44900
rect 19300 44888 19306 44940
rect 19429 44931 19487 44937
rect 19429 44897 19441 44931
rect 19475 44928 19487 44931
rect 19702 44928 19708 44940
rect 19475 44900 19708 44928
rect 19475 44897 19487 44900
rect 19429 44891 19487 44897
rect 19702 44888 19708 44900
rect 19760 44888 19766 44940
rect 22281 44931 22339 44937
rect 22281 44897 22293 44931
rect 22327 44928 22339 44931
rect 22646 44928 22652 44940
rect 22327 44900 22652 44928
rect 22327 44897 22339 44900
rect 22281 44891 22339 44897
rect 22646 44888 22652 44900
rect 22704 44888 22710 44940
rect 27433 44931 27491 44937
rect 27433 44897 27445 44931
rect 27479 44928 27491 44931
rect 27614 44928 27620 44940
rect 27479 44900 27620 44928
rect 27479 44897 27491 44900
rect 27433 44891 27491 44897
rect 27614 44888 27620 44900
rect 27672 44888 27678 44940
rect 17034 44820 17040 44872
rect 17092 44860 17098 44872
rect 17313 44863 17371 44869
rect 17313 44860 17325 44863
rect 17092 44832 17325 44860
rect 17092 44820 17098 44832
rect 17313 44829 17325 44832
rect 17359 44829 17371 44863
rect 17313 44823 17371 44829
rect 17405 44863 17463 44869
rect 17405 44829 17417 44863
rect 17451 44860 17463 44863
rect 17770 44860 17776 44872
rect 17451 44832 17776 44860
rect 17451 44829 17463 44832
rect 17405 44823 17463 44829
rect 17770 44820 17776 44832
rect 17828 44820 17834 44872
rect 18509 44863 18567 44869
rect 18509 44829 18521 44863
rect 18555 44860 18567 44863
rect 19334 44860 19340 44872
rect 18555 44832 19340 44860
rect 18555 44829 18567 44832
rect 18509 44823 18567 44829
rect 19334 44820 19340 44832
rect 19392 44820 19398 44872
rect 20806 44820 20812 44872
rect 20864 44820 20870 44872
rect 22097 44863 22155 44869
rect 22097 44829 22109 44863
rect 22143 44860 22155 44863
rect 24946 44860 24952 44872
rect 22143 44832 24952 44860
rect 22143 44829 22155 44832
rect 22097 44823 22155 44829
rect 24946 44820 24952 44832
rect 25004 44820 25010 44872
rect 26329 44863 26387 44869
rect 26329 44829 26341 44863
rect 26375 44860 26387 44863
rect 27157 44863 27215 44869
rect 27157 44860 27169 44863
rect 26375 44832 27169 44860
rect 26375 44829 26387 44832
rect 26329 44823 26387 44829
rect 27157 44829 27169 44832
rect 27203 44860 27215 44863
rect 46842 44860 46848 44872
rect 27203 44832 46848 44860
rect 27203 44829 27215 44832
rect 27157 44823 27215 44829
rect 19610 44792 19616 44804
rect 15436 44764 16528 44792
rect 16868 44764 19616 44792
rect 15436 44752 15442 44764
rect 14277 44727 14335 44733
rect 14277 44693 14289 44727
rect 14323 44693 14335 44727
rect 14277 44687 14335 44693
rect 15286 44684 15292 44736
rect 15344 44724 15350 44736
rect 15749 44727 15807 44733
rect 15749 44724 15761 44727
rect 15344 44696 15761 44724
rect 15344 44684 15350 44696
rect 15749 44693 15761 44696
rect 15795 44693 15807 44727
rect 15749 44687 15807 44693
rect 16114 44684 16120 44736
rect 16172 44684 16178 44736
rect 16209 44727 16267 44733
rect 16209 44693 16221 44727
rect 16255 44724 16267 44727
rect 16868 44724 16896 44764
rect 19610 44752 19616 44764
rect 19668 44752 19674 44804
rect 19702 44752 19708 44804
rect 19760 44752 19766 44804
rect 23658 44752 23664 44804
rect 23716 44792 23722 44804
rect 26344 44792 26372 44823
rect 46842 44820 46848 44832
rect 46900 44820 46906 44872
rect 44358 44792 44364 44804
rect 23716 44764 26372 44792
rect 28966 44764 44364 44792
rect 23716 44752 23722 44764
rect 16255 44696 16896 44724
rect 16255 44693 16267 44696
rect 16209 44687 16267 44693
rect 19518 44684 19524 44736
rect 19576 44724 19582 44736
rect 20070 44724 20076 44736
rect 19576 44696 20076 44724
rect 19576 44684 19582 44696
rect 20070 44684 20076 44696
rect 20128 44724 20134 44736
rect 21177 44727 21235 44733
rect 21177 44724 21189 44727
rect 20128 44696 21189 44724
rect 20128 44684 20134 44696
rect 21177 44693 21189 44696
rect 21223 44693 21235 44727
rect 21177 44687 21235 44693
rect 21634 44684 21640 44736
rect 21692 44684 21698 44736
rect 22002 44684 22008 44736
rect 22060 44684 22066 44736
rect 26786 44684 26792 44736
rect 26844 44684 26850 44736
rect 27246 44684 27252 44736
rect 27304 44724 27310 44736
rect 27985 44727 28043 44733
rect 27985 44724 27997 44727
rect 27304 44696 27997 44724
rect 27304 44684 27310 44696
rect 27985 44693 27997 44696
rect 28031 44724 28043 44727
rect 28966 44724 28994 44764
rect 44358 44752 44364 44764
rect 44416 44752 44422 44804
rect 28031 44696 28994 44724
rect 28031 44693 28043 44696
rect 27985 44687 28043 44693
rect 1104 44634 49864 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 27950 44634
rect 28002 44582 28014 44634
rect 28066 44582 28078 44634
rect 28130 44582 28142 44634
rect 28194 44582 28206 44634
rect 28258 44582 37950 44634
rect 38002 44582 38014 44634
rect 38066 44582 38078 44634
rect 38130 44582 38142 44634
rect 38194 44582 38206 44634
rect 38258 44582 47950 44634
rect 48002 44582 48014 44634
rect 48066 44582 48078 44634
rect 48130 44582 48142 44634
rect 48194 44582 48206 44634
rect 48258 44582 49864 44634
rect 1104 44560 49864 44582
rect 4154 44480 4160 44532
rect 4212 44520 4218 44532
rect 4525 44523 4583 44529
rect 4525 44520 4537 44523
rect 4212 44492 4537 44520
rect 4212 44480 4218 44492
rect 4525 44489 4537 44492
rect 4571 44489 4583 44523
rect 4525 44483 4583 44489
rect 6822 44480 6828 44532
rect 6880 44520 6886 44532
rect 8573 44523 8631 44529
rect 8573 44520 8585 44523
rect 6880 44492 8585 44520
rect 6880 44480 6886 44492
rect 8573 44489 8585 44492
rect 8619 44489 8631 44523
rect 8573 44483 8631 44489
rect 11974 44480 11980 44532
rect 12032 44520 12038 44532
rect 12805 44523 12863 44529
rect 12805 44520 12817 44523
rect 12032 44492 12817 44520
rect 12032 44480 12038 44492
rect 12805 44489 12817 44492
rect 12851 44489 12863 44523
rect 12805 44483 12863 44489
rect 13906 44480 13912 44532
rect 13964 44520 13970 44532
rect 17126 44520 17132 44532
rect 13964 44492 17132 44520
rect 13964 44480 13970 44492
rect 17126 44480 17132 44492
rect 17184 44480 17190 44532
rect 17497 44523 17555 44529
rect 17497 44489 17509 44523
rect 17543 44520 17555 44523
rect 18690 44520 18696 44532
rect 17543 44492 18696 44520
rect 17543 44489 17555 44492
rect 17497 44483 17555 44489
rect 18690 44480 18696 44492
rect 18748 44480 18754 44532
rect 20257 44523 20315 44529
rect 20257 44489 20269 44523
rect 20303 44489 20315 44523
rect 23290 44520 23296 44532
rect 20257 44483 20315 44489
rect 20364 44492 23296 44520
rect 3789 44455 3847 44461
rect 3789 44421 3801 44455
rect 3835 44452 3847 44455
rect 4246 44452 4252 44464
rect 3835 44424 4252 44452
rect 3835 44421 3847 44424
rect 3789 44415 3847 44421
rect 4246 44412 4252 44424
rect 4304 44412 4310 44464
rect 4433 44455 4491 44461
rect 4433 44421 4445 44455
rect 4479 44452 4491 44455
rect 5534 44452 5540 44464
rect 4479 44424 5540 44452
rect 4479 44421 4491 44424
rect 4433 44415 4491 44421
rect 5534 44412 5540 44424
rect 5592 44412 5598 44464
rect 9309 44455 9367 44461
rect 9309 44421 9321 44455
rect 9355 44452 9367 44455
rect 9950 44452 9956 44464
rect 9355 44424 9956 44452
rect 9355 44421 9367 44424
rect 9309 44415 9367 44421
rect 9950 44412 9956 44424
rect 10008 44452 10014 44464
rect 10410 44452 10416 44464
rect 10008 44424 10416 44452
rect 10008 44412 10014 44424
rect 10410 44412 10416 44424
rect 10468 44412 10474 44464
rect 13078 44452 13084 44464
rect 12406 44424 13084 44452
rect 1765 44387 1823 44393
rect 1765 44353 1777 44387
rect 1811 44384 1823 44387
rect 1811 44356 2774 44384
rect 1811 44353 1823 44356
rect 1765 44347 1823 44353
rect 2038 44276 2044 44328
rect 2096 44276 2102 44328
rect 2746 44316 2774 44356
rect 3510 44344 3516 44396
rect 3568 44384 3574 44396
rect 3605 44387 3663 44393
rect 3605 44384 3617 44387
rect 3568 44356 3617 44384
rect 3568 44344 3574 44356
rect 3605 44353 3617 44356
rect 3651 44353 3663 44387
rect 3605 44347 3663 44353
rect 8754 44344 8760 44396
rect 8812 44344 8818 44396
rect 10226 44344 10232 44396
rect 10284 44384 10290 44396
rect 12406 44384 12434 44424
rect 13078 44412 13084 44424
rect 13136 44412 13142 44464
rect 19886 44412 19892 44464
rect 19944 44452 19950 44464
rect 20272 44452 20300 44483
rect 19944 44424 20300 44452
rect 19944 44412 19950 44424
rect 10284 44356 12434 44384
rect 10284 44344 10290 44356
rect 12802 44344 12808 44396
rect 12860 44384 12866 44396
rect 12989 44387 13047 44393
rect 12989 44384 13001 44387
rect 12860 44356 13001 44384
rect 12860 44344 12866 44356
rect 12989 44353 13001 44356
rect 13035 44353 13047 44387
rect 12989 44347 13047 44353
rect 16114 44344 16120 44396
rect 16172 44384 16178 44396
rect 17037 44387 17095 44393
rect 17037 44384 17049 44387
rect 16172 44356 17049 44384
rect 16172 44344 16178 44356
rect 17037 44353 17049 44356
rect 17083 44353 17095 44387
rect 17037 44347 17095 44353
rect 17681 44387 17739 44393
rect 17681 44353 17693 44387
rect 17727 44353 17739 44387
rect 17681 44347 17739 44353
rect 4154 44316 4160 44328
rect 2746 44288 4160 44316
rect 4154 44276 4160 44288
rect 4212 44276 4218 44328
rect 17696 44316 17724 44347
rect 17770 44344 17776 44396
rect 17828 44384 17834 44396
rect 18325 44387 18383 44393
rect 18325 44384 18337 44387
rect 17828 44356 18337 44384
rect 17828 44344 17834 44356
rect 18325 44353 18337 44356
rect 18371 44353 18383 44387
rect 18325 44347 18383 44353
rect 19150 44344 19156 44396
rect 19208 44344 19214 44396
rect 19245 44387 19303 44393
rect 19245 44353 19257 44387
rect 19291 44384 19303 44387
rect 20364 44384 20392 44492
rect 23290 44480 23296 44492
rect 23348 44480 23354 44532
rect 20438 44412 20444 44464
rect 20496 44452 20502 44464
rect 20717 44455 20775 44461
rect 20717 44452 20729 44455
rect 20496 44424 20729 44452
rect 20496 44412 20502 44424
rect 20717 44421 20729 44424
rect 20763 44421 20775 44455
rect 20717 44415 20775 44421
rect 23566 44412 23572 44464
rect 23624 44452 23630 44464
rect 23842 44452 23848 44464
rect 23624 44424 23848 44452
rect 23624 44412 23630 44424
rect 23842 44412 23848 44424
rect 23900 44452 23906 44464
rect 23900 44424 25622 44452
rect 23900 44412 23906 44424
rect 19291 44356 20392 44384
rect 20625 44387 20683 44393
rect 19291 44353 19303 44356
rect 19245 44347 19303 44353
rect 20625 44353 20637 44387
rect 20671 44384 20683 44387
rect 20898 44384 20904 44396
rect 20671 44356 20904 44384
rect 20671 44353 20683 44356
rect 20625 44347 20683 44353
rect 20898 44344 20904 44356
rect 20956 44344 20962 44396
rect 22002 44344 22008 44396
rect 22060 44384 22066 44396
rect 22189 44387 22247 44393
rect 22189 44384 22201 44387
rect 22060 44356 22201 44384
rect 22060 44344 22066 44356
rect 22189 44353 22201 44356
rect 22235 44353 22247 44387
rect 22189 44347 22247 44353
rect 22830 44344 22836 44396
rect 22888 44384 22894 44396
rect 24857 44387 24915 44393
rect 24857 44384 24869 44387
rect 22888 44356 24869 44384
rect 22888 44344 22894 44356
rect 24857 44353 24869 44356
rect 24903 44353 24915 44387
rect 24857 44347 24915 44353
rect 18414 44316 18420 44328
rect 17696 44288 18420 44316
rect 18414 44276 18420 44288
rect 18472 44276 18478 44328
rect 19429 44319 19487 44325
rect 19429 44285 19441 44319
rect 19475 44316 19487 44319
rect 19978 44316 19984 44328
rect 19475 44288 19984 44316
rect 19475 44285 19487 44288
rect 19429 44279 19487 44285
rect 19978 44276 19984 44288
rect 20036 44276 20042 44328
rect 20809 44319 20867 44325
rect 20809 44285 20821 44319
rect 20855 44285 20867 44319
rect 20809 44279 20867 44285
rect 25133 44319 25191 44325
rect 25133 44285 25145 44319
rect 25179 44316 25191 44319
rect 27614 44316 27620 44328
rect 25179 44288 27620 44316
rect 25179 44285 25191 44288
rect 25133 44279 25191 44285
rect 13814 44208 13820 44260
rect 13872 44248 13878 44260
rect 18785 44251 18843 44257
rect 18785 44248 18797 44251
rect 13872 44220 18797 44248
rect 13872 44208 13878 44220
rect 18785 44217 18797 44220
rect 18831 44217 18843 44251
rect 18785 44211 18843 44217
rect 19702 44208 19708 44260
rect 19760 44248 19766 44260
rect 20530 44248 20536 44260
rect 19760 44220 20536 44248
rect 19760 44208 19766 44220
rect 20530 44208 20536 44220
rect 20588 44248 20594 44260
rect 20824 44248 20852 44279
rect 27614 44276 27620 44288
rect 27672 44276 27678 44328
rect 20588 44220 20852 44248
rect 20588 44208 20594 44220
rect 9398 44140 9404 44192
rect 9456 44140 9462 44192
rect 10778 44140 10784 44192
rect 10836 44180 10842 44192
rect 11057 44183 11115 44189
rect 11057 44180 11069 44183
rect 10836 44152 11069 44180
rect 10836 44140 10842 44152
rect 11057 44149 11069 44152
rect 11103 44149 11115 44183
rect 11057 44143 11115 44149
rect 12342 44140 12348 44192
rect 12400 44140 12406 44192
rect 18141 44183 18199 44189
rect 18141 44149 18153 44183
rect 18187 44180 18199 44183
rect 21358 44180 21364 44192
rect 18187 44152 21364 44180
rect 18187 44149 18199 44152
rect 18141 44143 18199 44149
rect 21358 44140 21364 44152
rect 21416 44140 21422 44192
rect 25222 44140 25228 44192
rect 25280 44180 25286 44192
rect 26605 44183 26663 44189
rect 26605 44180 26617 44183
rect 25280 44152 26617 44180
rect 25280 44140 25286 44152
rect 26605 44149 26617 44152
rect 26651 44149 26663 44183
rect 26605 44143 26663 44149
rect 1104 44090 49864 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 32950 44090
rect 33002 44038 33014 44090
rect 33066 44038 33078 44090
rect 33130 44038 33142 44090
rect 33194 44038 33206 44090
rect 33258 44038 42950 44090
rect 43002 44038 43014 44090
rect 43066 44038 43078 44090
rect 43130 44038 43142 44090
rect 43194 44038 43206 44090
rect 43258 44038 49864 44090
rect 1104 44016 49864 44038
rect 4430 43936 4436 43988
rect 4488 43976 4494 43988
rect 5077 43979 5135 43985
rect 5077 43976 5089 43979
rect 4488 43948 5089 43976
rect 4488 43936 4494 43948
rect 5077 43945 5089 43948
rect 5123 43945 5135 43979
rect 5077 43939 5135 43945
rect 5810 43936 5816 43988
rect 5868 43976 5874 43988
rect 10689 43979 10747 43985
rect 10689 43976 10701 43979
rect 5868 43948 10701 43976
rect 5868 43936 5874 43948
rect 10689 43945 10701 43948
rect 10735 43945 10747 43979
rect 10689 43939 10747 43945
rect 11238 43936 11244 43988
rect 11296 43936 11302 43988
rect 13449 43979 13507 43985
rect 13449 43976 13461 43979
rect 11348 43948 13461 43976
rect 9674 43868 9680 43920
rect 9732 43908 9738 43920
rect 11348 43908 11376 43948
rect 13449 43945 13461 43948
rect 13495 43945 13507 43979
rect 13449 43939 13507 43945
rect 17678 43936 17684 43988
rect 17736 43936 17742 43988
rect 18877 43979 18935 43985
rect 18877 43945 18889 43979
rect 18923 43976 18935 43979
rect 19150 43976 19156 43988
rect 18923 43948 19156 43976
rect 18923 43945 18935 43948
rect 18877 43939 18935 43945
rect 19150 43936 19156 43948
rect 19208 43936 19214 43988
rect 20898 43936 20904 43988
rect 20956 43936 20962 43988
rect 24026 43936 24032 43988
rect 24084 43936 24090 43988
rect 24946 43936 24952 43988
rect 25004 43976 25010 43988
rect 26789 43979 26847 43985
rect 26789 43976 26801 43979
rect 25004 43948 26801 43976
rect 25004 43936 25010 43948
rect 26789 43945 26801 43948
rect 26835 43976 26847 43979
rect 26835 43948 27936 43976
rect 26835 43945 26847 43948
rect 26789 43939 26847 43945
rect 14277 43911 14335 43917
rect 14277 43908 14289 43911
rect 9732 43880 11376 43908
rect 11440 43880 14289 43908
rect 9732 43868 9738 43880
rect 7282 43800 7288 43852
rect 7340 43840 7346 43852
rect 11440 43840 11468 43880
rect 14277 43877 14289 43880
rect 14323 43877 14335 43911
rect 21634 43908 21640 43920
rect 14277 43871 14335 43877
rect 17052 43880 21640 43908
rect 7340 43812 11468 43840
rect 7340 43800 7346 43812
rect 11790 43800 11796 43852
rect 11848 43800 11854 43852
rect 13814 43840 13820 43852
rect 13004 43812 13820 43840
rect 4985 43775 5043 43781
rect 4985 43741 4997 43775
rect 5031 43772 5043 43775
rect 7006 43772 7012 43784
rect 5031 43744 7012 43772
rect 5031 43741 5043 43744
rect 4985 43735 5043 43741
rect 7006 43732 7012 43744
rect 7064 43772 7070 43784
rect 7650 43772 7656 43784
rect 7064 43744 7656 43772
rect 7064 43732 7070 43744
rect 7650 43732 7656 43744
rect 7708 43732 7714 43784
rect 10597 43775 10655 43781
rect 10597 43741 10609 43775
rect 10643 43772 10655 43775
rect 11330 43772 11336 43784
rect 10643 43744 11336 43772
rect 10643 43741 10655 43744
rect 10597 43735 10655 43741
rect 11330 43732 11336 43744
rect 11388 43732 11394 43784
rect 11609 43775 11667 43781
rect 11609 43741 11621 43775
rect 11655 43772 11667 43775
rect 12526 43772 12532 43784
rect 11655 43744 12532 43772
rect 11655 43741 11667 43744
rect 11609 43735 11667 43741
rect 12526 43732 12532 43744
rect 12584 43732 12590 43784
rect 13004 43781 13032 43812
rect 13814 43800 13820 43812
rect 13872 43800 13878 43852
rect 13998 43800 14004 43852
rect 14056 43840 14062 43852
rect 17052 43840 17080 43880
rect 21634 43868 21640 43880
rect 21692 43868 21698 43920
rect 24854 43868 24860 43920
rect 24912 43908 24918 43920
rect 24912 43880 27016 43908
rect 24912 43868 24918 43880
rect 14056 43812 17080 43840
rect 14056 43800 14062 43812
rect 20070 43800 20076 43852
rect 20128 43800 20134 43852
rect 22557 43843 22615 43849
rect 22557 43809 22569 43843
rect 22603 43840 22615 43843
rect 23566 43840 23572 43852
rect 22603 43812 23572 43840
rect 22603 43809 22615 43812
rect 22557 43803 22615 43809
rect 23566 43800 23572 43812
rect 23624 43840 23630 43852
rect 24578 43840 24584 43852
rect 23624 43812 24584 43840
rect 23624 43800 23630 43812
rect 24578 43800 24584 43812
rect 24636 43800 24642 43852
rect 25222 43800 25228 43852
rect 25280 43800 25286 43852
rect 12989 43775 13047 43781
rect 12989 43741 13001 43775
rect 13035 43741 13047 43775
rect 12989 43735 13047 43741
rect 13633 43775 13691 43781
rect 13633 43741 13645 43775
rect 13679 43772 13691 43775
rect 13906 43772 13912 43784
rect 13679 43744 13912 43772
rect 13679 43741 13691 43744
rect 13633 43735 13691 43741
rect 13906 43732 13912 43744
rect 13964 43732 13970 43784
rect 14461 43775 14519 43781
rect 14461 43741 14473 43775
rect 14507 43772 14519 43775
rect 15010 43772 15016 43784
rect 14507 43744 15016 43772
rect 14507 43741 14519 43744
rect 14461 43735 14519 43741
rect 15010 43732 15016 43744
rect 15068 43732 15074 43784
rect 15194 43732 15200 43784
rect 15252 43772 15258 43784
rect 15470 43772 15476 43784
rect 15252 43744 15476 43772
rect 15252 43732 15258 43744
rect 15470 43732 15476 43744
rect 15528 43732 15534 43784
rect 17218 43732 17224 43784
rect 17276 43772 17282 43784
rect 17865 43775 17923 43781
rect 17865 43772 17877 43775
rect 17276 43744 17877 43772
rect 17276 43732 17282 43744
rect 17865 43741 17877 43744
rect 17911 43741 17923 43775
rect 17865 43735 17923 43741
rect 19886 43732 19892 43784
rect 19944 43732 19950 43784
rect 21818 43732 21824 43784
rect 21876 43732 21882 43784
rect 22278 43732 22284 43784
rect 22336 43732 22342 43784
rect 25041 43775 25099 43781
rect 25041 43741 25053 43775
rect 25087 43772 25099 43775
rect 26786 43772 26792 43784
rect 25087 43744 26792 43772
rect 25087 43741 25099 43744
rect 25041 43735 25099 43741
rect 26786 43732 26792 43744
rect 26844 43732 26850 43784
rect 26988 43772 27016 43880
rect 27614 43800 27620 43852
rect 27672 43840 27678 43852
rect 27801 43843 27859 43849
rect 27801 43840 27813 43843
rect 27672 43812 27813 43840
rect 27672 43800 27678 43812
rect 27801 43809 27813 43812
rect 27847 43809 27859 43843
rect 27801 43803 27859 43809
rect 27709 43775 27767 43781
rect 26988 43744 27660 43772
rect 11701 43707 11759 43713
rect 11701 43673 11713 43707
rect 11747 43704 11759 43707
rect 13354 43704 13360 43716
rect 11747 43676 13360 43704
rect 11747 43673 11759 43676
rect 11701 43667 11759 43673
rect 13354 43664 13360 43676
rect 13412 43664 13418 43716
rect 15746 43664 15752 43716
rect 15804 43664 15810 43716
rect 16022 43664 16028 43716
rect 16080 43704 16086 43716
rect 16206 43704 16212 43716
rect 16080 43676 16212 43704
rect 16080 43664 16086 43676
rect 16206 43664 16212 43676
rect 16264 43664 16270 43716
rect 23842 43704 23848 43716
rect 23782 43676 23848 43704
rect 23842 43664 23848 43676
rect 23900 43664 23906 43716
rect 27632 43713 27660 43744
rect 27709 43741 27721 43775
rect 27755 43772 27767 43775
rect 27908 43772 27936 43948
rect 27755 43744 31754 43772
rect 27755 43741 27767 43744
rect 27709 43735 27767 43741
rect 24949 43707 25007 43713
rect 23952 43676 24716 43704
rect 7466 43596 7472 43648
rect 7524 43636 7530 43648
rect 12805 43639 12863 43645
rect 12805 43636 12817 43639
rect 7524 43608 12817 43636
rect 7524 43596 7530 43608
rect 12805 43605 12817 43608
rect 12851 43605 12863 43639
rect 12805 43599 12863 43605
rect 13262 43596 13268 43648
rect 13320 43636 13326 43648
rect 16666 43636 16672 43648
rect 13320 43608 16672 43636
rect 13320 43596 13326 43608
rect 16666 43596 16672 43608
rect 16724 43596 16730 43648
rect 16758 43596 16764 43648
rect 16816 43636 16822 43648
rect 17221 43639 17279 43645
rect 17221 43636 17233 43639
rect 16816 43608 17233 43636
rect 16816 43596 16822 43608
rect 17221 43605 17233 43608
rect 17267 43605 17279 43639
rect 17221 43599 17279 43605
rect 17310 43596 17316 43648
rect 17368 43636 17374 43648
rect 19521 43639 19579 43645
rect 19521 43636 19533 43639
rect 17368 43608 19533 43636
rect 17368 43596 17374 43608
rect 19521 43605 19533 43608
rect 19567 43605 19579 43639
rect 19521 43599 19579 43605
rect 19981 43639 20039 43645
rect 19981 43605 19993 43639
rect 20027 43636 20039 43639
rect 23952 43636 23980 43676
rect 20027 43608 23980 43636
rect 20027 43605 20039 43608
rect 19981 43599 20039 43605
rect 24578 43596 24584 43648
rect 24636 43596 24642 43648
rect 24688 43636 24716 43676
rect 24949 43673 24961 43707
rect 24995 43704 25007 43707
rect 27617 43707 27675 43713
rect 24995 43676 27292 43704
rect 24995 43673 25007 43676
rect 24949 43667 25007 43673
rect 25774 43636 25780 43648
rect 24688 43608 25780 43636
rect 25774 43596 25780 43608
rect 25832 43596 25838 43648
rect 27264 43645 27292 43676
rect 27617 43673 27629 43707
rect 27663 43704 27675 43707
rect 28445 43707 28503 43713
rect 28445 43704 28457 43707
rect 27663 43676 28457 43704
rect 27663 43673 27675 43676
rect 27617 43667 27675 43673
rect 28445 43673 28457 43676
rect 28491 43673 28503 43707
rect 31726 43704 31754 43744
rect 48590 43704 48596 43716
rect 31726 43676 48596 43704
rect 28445 43667 28503 43673
rect 27249 43639 27307 43645
rect 27249 43605 27261 43639
rect 27295 43605 27307 43639
rect 28460 43636 28488 43667
rect 48590 43664 48596 43676
rect 48648 43664 48654 43716
rect 49234 43636 49240 43648
rect 28460 43608 49240 43636
rect 27249 43599 27307 43605
rect 49234 43596 49240 43608
rect 49292 43596 49298 43648
rect 1104 43546 49864 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 27950 43546
rect 28002 43494 28014 43546
rect 28066 43494 28078 43546
rect 28130 43494 28142 43546
rect 28194 43494 28206 43546
rect 28258 43494 37950 43546
rect 38002 43494 38014 43546
rect 38066 43494 38078 43546
rect 38130 43494 38142 43546
rect 38194 43494 38206 43546
rect 38258 43494 47950 43546
rect 48002 43494 48014 43546
rect 48066 43494 48078 43546
rect 48130 43494 48142 43546
rect 48194 43494 48206 43546
rect 48258 43494 49864 43546
rect 1104 43472 49864 43494
rect 9766 43392 9772 43444
rect 9824 43392 9830 43444
rect 9858 43392 9864 43444
rect 9916 43432 9922 43444
rect 10413 43435 10471 43441
rect 10413 43432 10425 43435
rect 9916 43404 10425 43432
rect 9916 43392 9922 43404
rect 10413 43401 10425 43404
rect 10459 43401 10471 43435
rect 10413 43395 10471 43401
rect 10778 43392 10784 43444
rect 10836 43392 10842 43444
rect 11422 43392 11428 43444
rect 11480 43432 11486 43444
rect 11701 43435 11759 43441
rect 11701 43432 11713 43435
rect 11480 43404 11713 43432
rect 11480 43392 11486 43404
rect 11701 43401 11713 43404
rect 11747 43401 11759 43435
rect 11701 43395 11759 43401
rect 12069 43435 12127 43441
rect 12069 43401 12081 43435
rect 12115 43432 12127 43435
rect 12342 43432 12348 43444
rect 12115 43404 12348 43432
rect 12115 43401 12127 43404
rect 12069 43395 12127 43401
rect 12342 43392 12348 43404
rect 12400 43392 12406 43444
rect 13449 43435 13507 43441
rect 13449 43401 13461 43435
rect 13495 43401 13507 43435
rect 13449 43395 13507 43401
rect 10873 43367 10931 43373
rect 10873 43333 10885 43367
rect 10919 43364 10931 43367
rect 12526 43364 12532 43376
rect 10919 43336 12532 43364
rect 10919 43333 10931 43336
rect 10873 43327 10931 43333
rect 12526 43324 12532 43336
rect 12584 43324 12590 43376
rect 1765 43299 1823 43305
rect 1765 43265 1777 43299
rect 1811 43296 1823 43299
rect 5350 43296 5356 43308
rect 1811 43268 5356 43296
rect 1811 43265 1823 43268
rect 1765 43259 1823 43265
rect 5350 43256 5356 43268
rect 5408 43256 5414 43308
rect 9125 43299 9183 43305
rect 9125 43265 9137 43299
rect 9171 43296 9183 43299
rect 9214 43296 9220 43308
rect 9171 43268 9220 43296
rect 9171 43265 9183 43268
rect 9125 43259 9183 43265
rect 9214 43256 9220 43268
rect 9272 43256 9278 43308
rect 9953 43299 10011 43305
rect 9953 43265 9965 43299
rect 9999 43296 10011 43299
rect 10042 43296 10048 43308
rect 9999 43268 10048 43296
rect 9999 43265 10011 43268
rect 9953 43259 10011 43265
rect 10042 43256 10048 43268
rect 10100 43256 10106 43308
rect 10152 43268 12388 43296
rect 1302 43188 1308 43240
rect 1360 43228 1366 43240
rect 2041 43231 2099 43237
rect 2041 43228 2053 43231
rect 1360 43200 2053 43228
rect 1360 43188 1366 43200
rect 2041 43197 2053 43200
rect 2087 43197 2099 43231
rect 2041 43191 2099 43197
rect 5074 43188 5080 43240
rect 5132 43228 5138 43240
rect 10152 43228 10180 43268
rect 5132 43200 10180 43228
rect 5132 43188 5138 43200
rect 10962 43188 10968 43240
rect 11020 43188 11026 43240
rect 12158 43188 12164 43240
rect 12216 43188 12222 43240
rect 12250 43188 12256 43240
rect 12308 43188 12314 43240
rect 12360 43228 12388 43268
rect 13464 43228 13492 43395
rect 13538 43392 13544 43444
rect 13596 43432 13602 43444
rect 14829 43435 14887 43441
rect 14829 43432 14841 43435
rect 13596 43404 14841 43432
rect 13596 43392 13602 43404
rect 14829 43401 14841 43404
rect 14875 43401 14887 43435
rect 14829 43395 14887 43401
rect 15289 43435 15347 43441
rect 15289 43401 15301 43435
rect 15335 43432 15347 43435
rect 17678 43432 17684 43444
rect 15335 43404 17684 43432
rect 15335 43401 15347 43404
rect 15289 43395 15347 43401
rect 17678 43392 17684 43404
rect 17736 43392 17742 43444
rect 17862 43392 17868 43444
rect 17920 43432 17926 43444
rect 17920 43404 18460 43432
rect 17920 43392 17926 43404
rect 14185 43367 14243 43373
rect 14185 43333 14197 43367
rect 14231 43364 14243 43367
rect 17310 43364 17316 43376
rect 14231 43336 17316 43364
rect 14231 43333 14243 43336
rect 14185 43327 14243 43333
rect 17310 43324 17316 43336
rect 17368 43324 17374 43376
rect 18322 43364 18328 43376
rect 18156 43336 18328 43364
rect 13633 43299 13691 43305
rect 13633 43265 13645 43299
rect 13679 43296 13691 43299
rect 13998 43296 14004 43308
rect 13679 43268 14004 43296
rect 13679 43265 13691 43268
rect 13633 43259 13691 43265
rect 13998 43256 14004 43268
rect 14056 43256 14062 43308
rect 14918 43256 14924 43308
rect 14976 43296 14982 43308
rect 15197 43299 15255 43305
rect 15197 43296 15209 43299
rect 14976 43268 15209 43296
rect 14976 43256 14982 43268
rect 15197 43265 15209 43268
rect 15243 43265 15255 43299
rect 15197 43259 15255 43265
rect 15838 43256 15844 43308
rect 15896 43296 15902 43308
rect 16301 43299 16359 43305
rect 16301 43296 16313 43299
rect 15896 43268 16313 43296
rect 15896 43256 15902 43268
rect 16301 43265 16313 43268
rect 16347 43265 16359 43299
rect 16301 43259 16359 43265
rect 17034 43256 17040 43308
rect 17092 43256 17098 43308
rect 17586 43256 17592 43308
rect 17644 43296 17650 43308
rect 17681 43299 17739 43305
rect 17681 43296 17693 43299
rect 17644 43268 17693 43296
rect 17644 43256 17650 43268
rect 17681 43265 17693 43268
rect 17727 43265 17739 43299
rect 17681 43259 17739 43265
rect 12360 43200 13492 43228
rect 15381 43231 15439 43237
rect 15381 43197 15393 43231
rect 15427 43197 15439 43231
rect 15381 43191 15439 43197
rect 9766 43120 9772 43172
rect 9824 43160 9830 43172
rect 11514 43160 11520 43172
rect 9824 43132 11520 43160
rect 9824 43120 9830 43132
rect 11514 43120 11520 43132
rect 11572 43120 11578 43172
rect 14369 43163 14427 43169
rect 14369 43160 14381 43163
rect 13372 43132 14381 43160
rect 9214 43052 9220 43104
rect 9272 43052 9278 43104
rect 9582 43052 9588 43104
rect 9640 43092 9646 43104
rect 13372 43092 13400 43132
rect 14369 43129 14381 43132
rect 14415 43129 14427 43163
rect 15396 43160 15424 43191
rect 15470 43188 15476 43240
rect 15528 43228 15534 43240
rect 18156 43237 18184 43336
rect 18322 43324 18328 43336
rect 18380 43324 18386 43376
rect 18432 43364 18460 43404
rect 19702 43392 19708 43444
rect 19760 43432 19766 43444
rect 19889 43435 19947 43441
rect 19889 43432 19901 43435
rect 19760 43404 19901 43432
rect 19760 43392 19766 43404
rect 19889 43401 19901 43404
rect 19935 43401 19947 43435
rect 19889 43395 19947 43401
rect 20717 43435 20775 43441
rect 20717 43401 20729 43435
rect 20763 43432 20775 43435
rect 21266 43432 21272 43444
rect 20763 43404 21272 43432
rect 20763 43401 20775 43404
rect 20717 43395 20775 43401
rect 21266 43392 21272 43404
rect 21324 43392 21330 43444
rect 21818 43392 21824 43444
rect 21876 43432 21882 43444
rect 22373 43435 22431 43441
rect 22373 43432 22385 43435
rect 21876 43404 22385 43432
rect 21876 43392 21882 43404
rect 22373 43401 22385 43404
rect 22419 43401 22431 43435
rect 22373 43395 22431 43401
rect 22462 43392 22468 43444
rect 22520 43392 22526 43444
rect 21177 43367 21235 43373
rect 18432 43336 18906 43364
rect 21177 43333 21189 43367
rect 21223 43364 21235 43367
rect 24578 43364 24584 43376
rect 21223 43336 24584 43364
rect 21223 43333 21235 43336
rect 21177 43327 21235 43333
rect 24578 43324 24584 43336
rect 24636 43324 24642 43376
rect 20806 43256 20812 43308
rect 20864 43296 20870 43308
rect 21085 43299 21143 43305
rect 21085 43296 21097 43299
rect 20864 43268 21097 43296
rect 20864 43256 20870 43268
rect 21085 43265 21097 43268
rect 21131 43265 21143 43299
rect 21085 43259 21143 43265
rect 18141 43231 18199 43237
rect 18141 43228 18153 43231
rect 15528 43200 18153 43228
rect 15528 43188 15534 43200
rect 18141 43197 18153 43200
rect 18187 43197 18199 43231
rect 18417 43231 18475 43237
rect 18417 43228 18429 43231
rect 18141 43191 18199 43197
rect 18248 43200 18429 43228
rect 17310 43160 17316 43172
rect 15396 43132 17316 43160
rect 14369 43123 14427 43129
rect 17310 43120 17316 43132
rect 17368 43160 17374 43172
rect 18248 43160 18276 43200
rect 18417 43197 18429 43200
rect 18463 43197 18475 43231
rect 18417 43191 18475 43197
rect 21358 43188 21364 43240
rect 21416 43188 21422 43240
rect 22649 43231 22707 43237
rect 22649 43197 22661 43231
rect 22695 43228 22707 43231
rect 23566 43228 23572 43240
rect 22695 43200 23572 43228
rect 22695 43197 22707 43200
rect 22649 43191 22707 43197
rect 23566 43188 23572 43200
rect 23624 43188 23630 43240
rect 17368 43132 18276 43160
rect 17368 43120 17374 43132
rect 9640 43064 13400 43092
rect 9640 43052 9646 43064
rect 15562 43052 15568 43104
rect 15620 43092 15626 43104
rect 16117 43095 16175 43101
rect 16117 43092 16129 43095
rect 15620 43064 16129 43092
rect 15620 43052 15626 43064
rect 16117 43061 16129 43064
rect 16163 43061 16175 43095
rect 16117 43055 16175 43061
rect 16666 43052 16672 43104
rect 16724 43092 16730 43104
rect 17497 43095 17555 43101
rect 17497 43092 17509 43095
rect 16724 43064 17509 43092
rect 16724 43052 16730 43064
rect 17497 43061 17509 43064
rect 17543 43061 17555 43095
rect 17497 43055 17555 43061
rect 17862 43052 17868 43104
rect 17920 43092 17926 43104
rect 22005 43095 22063 43101
rect 22005 43092 22017 43095
rect 17920 43064 22017 43092
rect 17920 43052 17926 43064
rect 22005 43061 22017 43064
rect 22051 43061 22063 43095
rect 22005 43055 22063 43061
rect 1104 43002 49864 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 32950 43002
rect 33002 42950 33014 43002
rect 33066 42950 33078 43002
rect 33130 42950 33142 43002
rect 33194 42950 33206 43002
rect 33258 42950 42950 43002
rect 43002 42950 43014 43002
rect 43066 42950 43078 43002
rect 43130 42950 43142 43002
rect 43194 42950 43206 43002
rect 43258 42950 49864 43002
rect 1104 42928 49864 42950
rect 6996 42891 7054 42897
rect 6996 42857 7008 42891
rect 7042 42888 7054 42891
rect 8938 42888 8944 42900
rect 7042 42860 8944 42888
rect 7042 42857 7054 42860
rect 6996 42851 7054 42857
rect 8938 42848 8944 42860
rect 8996 42848 9002 42900
rect 11517 42891 11575 42897
rect 11517 42857 11529 42891
rect 11563 42888 11575 42891
rect 11790 42888 11796 42900
rect 11563 42860 11796 42888
rect 11563 42857 11575 42860
rect 11517 42851 11575 42857
rect 11790 42848 11796 42860
rect 11848 42888 11854 42900
rect 12234 42891 12292 42897
rect 12234 42888 12246 42891
rect 11848 42860 12246 42888
rect 11848 42848 11854 42860
rect 12234 42857 12246 42860
rect 12280 42857 12292 42891
rect 12234 42851 12292 42857
rect 14182 42848 14188 42900
rect 14240 42888 14246 42900
rect 16098 42891 16156 42897
rect 16098 42888 16110 42891
rect 14240 42860 16110 42888
rect 14240 42848 14246 42860
rect 16098 42857 16110 42860
rect 16144 42888 16156 42891
rect 16758 42888 16764 42900
rect 16144 42860 16764 42888
rect 16144 42857 16156 42860
rect 16098 42851 16156 42857
rect 16758 42848 16764 42860
rect 16816 42888 16822 42900
rect 20254 42888 20260 42900
rect 16816 42860 20260 42888
rect 16816 42848 16822 42860
rect 20254 42848 20260 42860
rect 20312 42848 20318 42900
rect 21072 42891 21130 42897
rect 21072 42857 21084 42891
rect 21118 42888 21130 42891
rect 24026 42888 24032 42900
rect 21118 42860 24032 42888
rect 21118 42857 21130 42860
rect 21072 42851 21130 42857
rect 24026 42848 24032 42860
rect 24084 42848 24090 42900
rect 1302 42712 1308 42764
rect 1360 42752 1366 42764
rect 2041 42755 2099 42761
rect 2041 42752 2053 42755
rect 1360 42724 2053 42752
rect 1360 42712 1366 42724
rect 2041 42721 2053 42724
rect 2087 42721 2099 42755
rect 2041 42715 2099 42721
rect 3694 42712 3700 42764
rect 3752 42752 3758 42764
rect 4801 42755 4859 42761
rect 4801 42752 4813 42755
rect 3752 42724 4813 42752
rect 3752 42712 3758 42724
rect 4801 42721 4813 42724
rect 4847 42721 4859 42755
rect 4801 42715 4859 42721
rect 6733 42755 6791 42761
rect 6733 42721 6745 42755
rect 6779 42752 6791 42755
rect 11977 42755 12035 42761
rect 11977 42752 11989 42755
rect 6779 42724 11989 42752
rect 6779 42721 6791 42724
rect 6733 42715 6791 42721
rect 11977 42721 11989 42724
rect 12023 42752 12035 42755
rect 15013 42755 15071 42761
rect 12023 42724 14872 42752
rect 12023 42721 12035 42724
rect 11977 42715 12035 42721
rect 1578 42644 1584 42696
rect 1636 42644 1642 42696
rect 4617 42687 4675 42693
rect 4617 42653 4629 42687
rect 4663 42684 4675 42687
rect 5626 42684 5632 42696
rect 4663 42656 5632 42684
rect 4663 42653 4675 42656
rect 4617 42647 4675 42653
rect 5626 42644 5632 42656
rect 5684 42684 5690 42696
rect 5994 42684 6000 42696
rect 5684 42656 6000 42684
rect 5684 42644 5690 42656
rect 5994 42644 6000 42656
rect 6052 42644 6058 42696
rect 9306 42644 9312 42696
rect 9364 42644 9370 42696
rect 9769 42687 9827 42693
rect 9769 42653 9781 42687
rect 9815 42653 9827 42687
rect 14844 42684 14872 42724
rect 15013 42721 15025 42755
rect 15059 42752 15071 42755
rect 15194 42752 15200 42764
rect 15059 42724 15200 42752
rect 15059 42721 15071 42724
rect 15013 42715 15071 42721
rect 15194 42712 15200 42724
rect 15252 42712 15258 42764
rect 17310 42712 17316 42764
rect 17368 42752 17374 42764
rect 17589 42755 17647 42761
rect 17589 42752 17601 42755
rect 17368 42724 17601 42752
rect 17368 42712 17374 42724
rect 17589 42721 17601 42724
rect 17635 42721 17647 42755
rect 17589 42715 17647 42721
rect 19978 42712 19984 42764
rect 20036 42712 20042 42764
rect 20809 42755 20867 42761
rect 20809 42721 20821 42755
rect 20855 42752 20867 42755
rect 21450 42752 21456 42764
rect 20855 42724 21456 42752
rect 20855 42721 20867 42724
rect 20809 42715 20867 42721
rect 21450 42712 21456 42724
rect 21508 42712 21514 42764
rect 21726 42712 21732 42764
rect 21784 42752 21790 42764
rect 21784 42724 22876 42752
rect 21784 42712 21790 42724
rect 15470 42684 15476 42696
rect 14844 42656 15476 42684
rect 9769 42647 9827 42653
rect 7558 42576 7564 42628
rect 7616 42576 7622 42628
rect 8312 42588 8616 42616
rect 7006 42508 7012 42560
rect 7064 42548 7070 42560
rect 8312 42548 8340 42588
rect 7064 42520 8340 42548
rect 7064 42508 7070 42520
rect 8478 42508 8484 42560
rect 8536 42508 8542 42560
rect 8588 42548 8616 42588
rect 8754 42576 8760 42628
rect 8812 42616 8818 42628
rect 9784 42616 9812 42647
rect 15470 42644 15476 42656
rect 15528 42684 15534 42696
rect 15841 42687 15899 42693
rect 15841 42684 15853 42687
rect 15528 42656 15853 42684
rect 15528 42644 15534 42656
rect 15841 42653 15853 42656
rect 15887 42653 15899 42687
rect 15841 42647 15899 42653
rect 18322 42644 18328 42696
rect 18380 42684 18386 42696
rect 18506 42684 18512 42696
rect 18380 42656 18512 42684
rect 18380 42644 18386 42656
rect 18506 42644 18512 42656
rect 18564 42644 18570 42696
rect 22848 42684 22876 42724
rect 22922 42712 22928 42764
rect 22980 42752 22986 42764
rect 48774 42752 48780 42764
rect 22980 42724 48780 42752
rect 22980 42712 22986 42724
rect 48774 42712 48780 42724
rect 48832 42712 48838 42764
rect 25130 42684 25136 42696
rect 22848 42656 25136 42684
rect 25130 42644 25136 42656
rect 25188 42644 25194 42696
rect 8812 42588 9812 42616
rect 10045 42619 10103 42625
rect 8812 42576 8818 42588
rect 10045 42585 10057 42619
rect 10091 42616 10103 42619
rect 10318 42616 10324 42628
rect 10091 42588 10324 42616
rect 10091 42585 10103 42588
rect 10045 42579 10103 42585
rect 10318 42576 10324 42588
rect 10376 42576 10382 42628
rect 11330 42616 11336 42628
rect 11270 42588 11336 42616
rect 11330 42576 11336 42588
rect 11388 42616 11394 42628
rect 12710 42616 12716 42628
rect 11388 42588 12716 42616
rect 11388 42576 11394 42588
rect 12710 42576 12716 42588
rect 12768 42576 12774 42628
rect 13814 42576 13820 42628
rect 13872 42616 13878 42628
rect 14737 42619 14795 42625
rect 14737 42616 14749 42619
rect 13872 42588 14749 42616
rect 13872 42576 13878 42588
rect 14737 42585 14749 42588
rect 14783 42585 14795 42619
rect 14737 42579 14795 42585
rect 16022 42576 16028 42628
rect 16080 42616 16086 42628
rect 18141 42619 18199 42625
rect 16080 42588 16606 42616
rect 16080 42576 16086 42588
rect 18141 42585 18153 42619
rect 18187 42616 18199 42619
rect 18690 42616 18696 42628
rect 18187 42588 18696 42616
rect 18187 42585 18199 42588
rect 18141 42579 18199 42585
rect 18690 42576 18696 42588
rect 18748 42576 18754 42628
rect 22462 42616 22468 42628
rect 22310 42588 22468 42616
rect 22462 42576 22468 42588
rect 22520 42616 22526 42628
rect 23842 42616 23848 42628
rect 22520 42588 23848 42616
rect 22520 42576 22526 42588
rect 23842 42576 23848 42588
rect 23900 42576 23906 42628
rect 9125 42551 9183 42557
rect 9125 42548 9137 42551
rect 8588 42520 9137 42548
rect 9125 42517 9137 42520
rect 9171 42517 9183 42551
rect 9125 42511 9183 42517
rect 13630 42508 13636 42560
rect 13688 42548 13694 42560
rect 13725 42551 13783 42557
rect 13725 42548 13737 42551
rect 13688 42520 13737 42548
rect 13688 42508 13694 42520
rect 13725 42517 13737 42520
rect 13771 42517 13783 42551
rect 13725 42511 13783 42517
rect 13906 42508 13912 42560
rect 13964 42548 13970 42560
rect 14369 42551 14427 42557
rect 14369 42548 14381 42551
rect 13964 42520 14381 42548
rect 13964 42508 13970 42520
rect 14369 42517 14381 42520
rect 14415 42517 14427 42551
rect 14369 42511 14427 42517
rect 14829 42551 14887 42557
rect 14829 42517 14841 42551
rect 14875 42548 14887 42551
rect 18506 42548 18512 42560
rect 14875 42520 18512 42548
rect 14875 42517 14887 42520
rect 14829 42511 14887 42517
rect 18506 42508 18512 42520
rect 18564 42508 18570 42560
rect 18782 42508 18788 42560
rect 18840 42508 18846 42560
rect 18966 42508 18972 42560
rect 19024 42548 19030 42560
rect 19429 42551 19487 42557
rect 19429 42548 19441 42551
rect 19024 42520 19441 42548
rect 19024 42508 19030 42520
rect 19429 42517 19441 42520
rect 19475 42517 19487 42551
rect 19429 42511 19487 42517
rect 19794 42508 19800 42560
rect 19852 42508 19858 42560
rect 19889 42551 19947 42557
rect 19889 42517 19901 42551
rect 19935 42548 19947 42551
rect 21726 42548 21732 42560
rect 19935 42520 21732 42548
rect 19935 42517 19947 42520
rect 19889 42511 19947 42517
rect 21726 42508 21732 42520
rect 21784 42508 21790 42560
rect 21910 42508 21916 42560
rect 21968 42548 21974 42560
rect 22557 42551 22615 42557
rect 22557 42548 22569 42551
rect 21968 42520 22569 42548
rect 21968 42508 21974 42520
rect 22557 42517 22569 42520
rect 22603 42517 22615 42551
rect 22557 42511 22615 42517
rect 1104 42458 49864 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 27950 42458
rect 28002 42406 28014 42458
rect 28066 42406 28078 42458
rect 28130 42406 28142 42458
rect 28194 42406 28206 42458
rect 28258 42406 37950 42458
rect 38002 42406 38014 42458
rect 38066 42406 38078 42458
rect 38130 42406 38142 42458
rect 38194 42406 38206 42458
rect 38258 42406 47950 42458
rect 48002 42406 48014 42458
rect 48066 42406 48078 42458
rect 48130 42406 48142 42458
rect 48194 42406 48206 42458
rect 48258 42406 49864 42458
rect 1104 42384 49864 42406
rect 4154 42304 4160 42356
rect 4212 42344 4218 42356
rect 4985 42347 5043 42353
rect 4985 42344 4997 42347
rect 4212 42316 4997 42344
rect 4212 42304 4218 42316
rect 4985 42313 4997 42316
rect 5031 42313 5043 42347
rect 4985 42307 5043 42313
rect 9306 42304 9312 42356
rect 9364 42344 9370 42356
rect 9364 42316 10916 42344
rect 9364 42304 9370 42316
rect 10888 42276 10916 42316
rect 12434 42304 12440 42356
rect 12492 42344 12498 42356
rect 13449 42347 13507 42353
rect 13449 42344 13461 42347
rect 12492 42316 13461 42344
rect 12492 42304 12498 42316
rect 13449 42313 13461 42316
rect 13495 42313 13507 42347
rect 13449 42307 13507 42313
rect 15194 42304 15200 42356
rect 15252 42344 15258 42356
rect 15746 42344 15752 42356
rect 15252 42316 15752 42344
rect 15252 42304 15258 42316
rect 15746 42304 15752 42316
rect 15804 42344 15810 42356
rect 16301 42347 16359 42353
rect 16301 42344 16313 42347
rect 15804 42316 16313 42344
rect 15804 42304 15810 42316
rect 16301 42313 16313 42316
rect 16347 42313 16359 42347
rect 16301 42307 16359 42313
rect 17221 42347 17279 42353
rect 17221 42313 17233 42347
rect 17267 42344 17279 42347
rect 18322 42344 18328 42356
rect 17267 42316 18328 42344
rect 17267 42313 17279 42316
rect 17221 42307 17279 42313
rect 18322 42304 18328 42316
rect 18380 42304 18386 42356
rect 18506 42304 18512 42356
rect 18564 42344 18570 42356
rect 20717 42347 20775 42353
rect 20717 42344 20729 42347
rect 18564 42316 20729 42344
rect 18564 42304 18570 42316
rect 20717 42313 20729 42316
rect 20763 42313 20775 42347
rect 20717 42307 20775 42313
rect 21082 42304 21088 42356
rect 21140 42304 21146 42356
rect 21358 42304 21364 42356
rect 21416 42344 21422 42356
rect 21818 42344 21824 42356
rect 21416 42316 21824 42344
rect 21416 42304 21422 42316
rect 21818 42304 21824 42316
rect 21876 42344 21882 42356
rect 24121 42347 24179 42353
rect 24121 42344 24133 42347
rect 21876 42316 24133 42344
rect 21876 42304 21882 42316
rect 24121 42313 24133 42316
rect 24167 42313 24179 42347
rect 24121 42307 24179 42313
rect 15102 42276 15108 42288
rect 10888 42248 15108 42276
rect 15102 42236 15108 42248
rect 15160 42236 15166 42288
rect 16390 42236 16396 42288
rect 16448 42276 16454 42288
rect 19702 42276 19708 42288
rect 16448 42248 19708 42276
rect 16448 42236 16454 42248
rect 19702 42236 19708 42248
rect 19760 42236 19766 42288
rect 20070 42236 20076 42288
rect 20128 42276 20134 42288
rect 21910 42276 21916 42288
rect 20128 42248 21916 42276
rect 20128 42236 20134 42248
rect 21910 42236 21916 42248
rect 21968 42236 21974 42288
rect 22922 42276 22928 42288
rect 22066 42248 22928 42276
rect 4893 42211 4951 42217
rect 4893 42177 4905 42211
rect 4939 42208 4951 42211
rect 4939 42180 7144 42208
rect 4939 42177 4951 42180
rect 4893 42171 4951 42177
rect 7116 42084 7144 42180
rect 8754 42168 8760 42220
rect 8812 42168 8818 42220
rect 11054 42208 11060 42220
rect 10166 42180 11060 42208
rect 11054 42168 11060 42180
rect 11112 42168 11118 42220
rect 11146 42168 11152 42220
rect 11204 42168 11210 42220
rect 11701 42211 11759 42217
rect 11701 42177 11713 42211
rect 11747 42208 11759 42211
rect 12158 42208 12164 42220
rect 11747 42180 12164 42208
rect 11747 42177 11759 42180
rect 11701 42171 11759 42177
rect 12158 42168 12164 42180
rect 12216 42168 12222 42220
rect 15930 42168 15936 42220
rect 15988 42168 15994 42220
rect 16758 42168 16764 42220
rect 16816 42208 16822 42220
rect 17405 42211 17463 42217
rect 17405 42208 17417 42211
rect 16816 42180 17417 42208
rect 16816 42168 16822 42180
rect 17405 42177 17417 42180
rect 17451 42177 17463 42211
rect 17405 42171 17463 42177
rect 17494 42168 17500 42220
rect 17552 42208 17558 42220
rect 18049 42211 18107 42217
rect 18049 42208 18061 42211
rect 17552 42180 18061 42208
rect 17552 42168 17558 42180
rect 18049 42177 18061 42180
rect 18095 42177 18107 42211
rect 18049 42171 18107 42177
rect 19337 42211 19395 42217
rect 19337 42177 19349 42211
rect 19383 42208 19395 42211
rect 19794 42208 19800 42220
rect 19383 42180 19800 42208
rect 19383 42177 19395 42180
rect 19337 42171 19395 42177
rect 19794 42168 19800 42180
rect 19852 42168 19858 42220
rect 19889 42211 19947 42217
rect 19889 42177 19901 42211
rect 19935 42177 19947 42211
rect 19889 42171 19947 42177
rect 19981 42211 20039 42217
rect 19981 42177 19993 42211
rect 20027 42208 20039 42211
rect 20162 42208 20168 42220
rect 20027 42180 20168 42208
rect 20027 42177 20039 42180
rect 19981 42171 20039 42177
rect 9030 42100 9036 42152
rect 9088 42100 9094 42152
rect 10410 42100 10416 42152
rect 10468 42140 10474 42152
rect 12437 42143 12495 42149
rect 12437 42140 12449 42143
rect 10468 42112 12449 42140
rect 10468 42100 10474 42112
rect 12437 42109 12449 42112
rect 12483 42109 12495 42143
rect 12437 42103 12495 42109
rect 13538 42100 13544 42152
rect 13596 42100 13602 42152
rect 13633 42143 13691 42149
rect 13633 42109 13645 42143
rect 13679 42109 13691 42143
rect 13633 42103 13691 42109
rect 7098 42032 7104 42084
rect 7156 42072 7162 42084
rect 7156 42044 8800 42072
rect 7156 42032 7162 42044
rect 8478 41964 8484 42016
rect 8536 42004 8542 42016
rect 8662 42004 8668 42016
rect 8536 41976 8668 42004
rect 8536 41964 8542 41976
rect 8662 41964 8668 41976
rect 8720 41964 8726 42016
rect 8772 42004 8800 42044
rect 10502 42032 10508 42084
rect 10560 42032 10566 42084
rect 11606 42032 11612 42084
rect 11664 42072 11670 42084
rect 13081 42075 13139 42081
rect 13081 42072 13093 42075
rect 11664 42044 13093 42072
rect 11664 42032 11670 42044
rect 13081 42041 13093 42044
rect 13127 42041 13139 42075
rect 13081 42035 13139 42041
rect 10965 42007 11023 42013
rect 10965 42004 10977 42007
rect 8772 41976 10977 42004
rect 10965 41973 10977 41976
rect 11011 41973 11023 42007
rect 10965 41967 11023 41973
rect 11974 41964 11980 42016
rect 12032 42004 12038 42016
rect 13648 42004 13676 42103
rect 14550 42100 14556 42152
rect 14608 42100 14614 42152
rect 14826 42100 14832 42152
rect 14884 42140 14890 42152
rect 17218 42140 17224 42152
rect 14884 42112 17224 42140
rect 14884 42100 14890 42112
rect 17218 42100 17224 42112
rect 17276 42100 17282 42152
rect 17862 42140 17868 42152
rect 17604 42112 17868 42140
rect 16022 42032 16028 42084
rect 16080 42072 16086 42084
rect 17604 42072 17632 42112
rect 17862 42100 17868 42112
rect 17920 42100 17926 42152
rect 18138 42100 18144 42152
rect 18196 42140 18202 42152
rect 18506 42140 18512 42152
rect 18196 42112 18512 42140
rect 18196 42100 18202 42112
rect 18506 42100 18512 42112
rect 18564 42100 18570 42152
rect 18690 42100 18696 42152
rect 18748 42140 18754 42152
rect 18969 42143 19027 42149
rect 18969 42140 18981 42143
rect 18748 42112 18981 42140
rect 18748 42100 18754 42112
rect 18969 42109 18981 42112
rect 19015 42140 19027 42143
rect 19904 42140 19932 42171
rect 20162 42168 20168 42180
rect 20220 42168 20226 42220
rect 20346 42168 20352 42220
rect 20404 42208 20410 42220
rect 20404 42180 21312 42208
rect 20404 42168 20410 42180
rect 19015 42112 19932 42140
rect 19015 42109 19027 42112
rect 18969 42103 19027 42109
rect 16080 42044 17632 42072
rect 16080 42032 16086 42044
rect 17678 42032 17684 42084
rect 17736 42072 17742 42084
rect 19521 42075 19579 42081
rect 19521 42072 19533 42075
rect 17736 42044 19533 42072
rect 17736 42032 17742 42044
rect 19521 42041 19533 42044
rect 19567 42041 19579 42075
rect 19904 42072 19932 42112
rect 20073 42143 20131 42149
rect 20073 42109 20085 42143
rect 20119 42140 20131 42143
rect 20254 42140 20260 42152
rect 20119 42112 20260 42140
rect 20119 42109 20131 42112
rect 20073 42103 20131 42109
rect 20254 42100 20260 42112
rect 20312 42100 20318 42152
rect 21284 42149 21312 42180
rect 21358 42168 21364 42220
rect 21416 42208 21422 42220
rect 22066 42208 22094 42248
rect 22922 42236 22928 42248
rect 22980 42236 22986 42288
rect 21416 42180 22094 42208
rect 21416 42168 21422 42180
rect 22278 42168 22284 42220
rect 22336 42208 22342 42220
rect 22373 42211 22431 42217
rect 22373 42208 22385 42211
rect 22336 42180 22385 42208
rect 22336 42168 22342 42180
rect 22373 42177 22385 42180
rect 22419 42177 22431 42211
rect 22373 42171 22431 42177
rect 23750 42168 23756 42220
rect 23808 42168 23814 42220
rect 21177 42143 21235 42149
rect 21177 42140 21189 42143
rect 21008 42112 21189 42140
rect 20898 42072 20904 42084
rect 19904 42044 20904 42072
rect 19521 42035 19579 42041
rect 20898 42032 20904 42044
rect 20956 42032 20962 42084
rect 21008 42072 21036 42112
rect 21177 42109 21189 42112
rect 21223 42109 21235 42143
rect 21177 42103 21235 42109
rect 21269 42143 21327 42149
rect 21269 42109 21281 42143
rect 21315 42109 21327 42143
rect 21269 42103 21327 42109
rect 21450 42100 21456 42152
rect 21508 42140 21514 42152
rect 22296 42140 22324 42168
rect 21508 42112 22324 42140
rect 21508 42100 21514 42112
rect 22646 42100 22652 42152
rect 22704 42140 22710 42152
rect 25222 42140 25228 42152
rect 22704 42112 25228 42140
rect 22704 42100 22710 42112
rect 25222 42100 25228 42112
rect 25280 42100 25286 42152
rect 22370 42072 22376 42084
rect 21008 42044 22376 42072
rect 12032 41976 13676 42004
rect 12032 41964 12038 41976
rect 13722 41964 13728 42016
rect 13780 42004 13786 42016
rect 14274 42004 14280 42016
rect 13780 41976 14280 42004
rect 13780 41964 13786 41976
rect 14274 41964 14280 41976
rect 14332 41964 14338 42016
rect 15562 41964 15568 42016
rect 15620 42004 15626 42016
rect 17865 42007 17923 42013
rect 17865 42004 17877 42007
rect 15620 41976 17877 42004
rect 15620 41964 15626 41976
rect 17865 41973 17877 41976
rect 17911 41973 17923 42007
rect 17865 41967 17923 41973
rect 17954 41964 17960 42016
rect 18012 42004 18018 42016
rect 19242 42004 19248 42016
rect 18012 41976 19248 42004
rect 18012 41964 18018 41976
rect 19242 41964 19248 41976
rect 19300 41964 19306 42016
rect 19702 41964 19708 42016
rect 19760 42004 19766 42016
rect 21008 42004 21036 42044
rect 22370 42032 22376 42044
rect 22428 42032 22434 42084
rect 24670 42032 24676 42084
rect 24728 42072 24734 42084
rect 48958 42072 48964 42084
rect 24728 42044 48964 42072
rect 24728 42032 24734 42044
rect 48958 42032 48964 42044
rect 49016 42032 49022 42084
rect 19760 41976 21036 42004
rect 19760 41964 19766 41976
rect 21082 41964 21088 42016
rect 21140 42004 21146 42016
rect 22281 42007 22339 42013
rect 22281 42004 22293 42007
rect 21140 41976 22293 42004
rect 21140 41964 21146 41976
rect 22281 41973 22293 41976
rect 22327 42004 22339 42007
rect 24688 42004 24716 42032
rect 22327 41976 24716 42004
rect 22327 41973 22339 41976
rect 22281 41967 22339 41973
rect 1104 41914 49864 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 32950 41914
rect 33002 41862 33014 41914
rect 33066 41862 33078 41914
rect 33130 41862 33142 41914
rect 33194 41862 33206 41914
rect 33258 41862 42950 41914
rect 43002 41862 43014 41914
rect 43066 41862 43078 41914
rect 43130 41862 43142 41914
rect 43194 41862 43206 41914
rect 43258 41862 49864 41914
rect 1104 41840 49864 41862
rect 4338 41760 4344 41812
rect 4396 41800 4402 41812
rect 4801 41803 4859 41809
rect 4801 41800 4813 41803
rect 4396 41772 4813 41800
rect 4396 41760 4402 41772
rect 4801 41769 4813 41772
rect 4847 41769 4859 41803
rect 10870 41800 10876 41812
rect 4801 41763 4859 41769
rect 10060 41772 10876 41800
rect 1762 41692 1768 41744
rect 1820 41732 1826 41744
rect 9953 41735 10011 41741
rect 9953 41732 9965 41735
rect 1820 41704 9965 41732
rect 1820 41692 1826 41704
rect 9953 41701 9965 41704
rect 9999 41701 10011 41735
rect 9953 41695 10011 41701
rect 1302 41624 1308 41676
rect 1360 41664 1366 41676
rect 2041 41667 2099 41673
rect 2041 41664 2053 41667
rect 1360 41636 2053 41664
rect 1360 41624 1366 41636
rect 2041 41633 2053 41636
rect 2087 41633 2099 41667
rect 9398 41664 9404 41676
rect 2041 41627 2099 41633
rect 2746 41636 9404 41664
rect 1765 41599 1823 41605
rect 1765 41565 1777 41599
rect 1811 41596 1823 41599
rect 2746 41596 2774 41636
rect 9398 41624 9404 41636
rect 9456 41624 9462 41676
rect 10060 41664 10088 41772
rect 10870 41760 10876 41772
rect 10928 41760 10934 41812
rect 11146 41760 11152 41812
rect 11204 41800 11210 41812
rect 11204 41772 12572 41800
rect 11204 41760 11210 41772
rect 11974 41732 11980 41744
rect 11716 41704 11980 41732
rect 9692 41636 10088 41664
rect 1811 41568 2774 41596
rect 4709 41599 4767 41605
rect 1811 41565 1823 41568
rect 1765 41559 1823 41565
rect 4709 41565 4721 41599
rect 4755 41596 4767 41599
rect 7006 41596 7012 41608
rect 4755 41568 7012 41596
rect 4755 41565 4767 41568
rect 4709 41559 4767 41565
rect 7006 41556 7012 41568
rect 7064 41556 7070 41608
rect 8294 41556 8300 41608
rect 8352 41596 8358 41608
rect 8573 41599 8631 41605
rect 8573 41596 8585 41599
rect 8352 41568 8585 41596
rect 8352 41556 8358 41568
rect 8573 41565 8585 41568
rect 8619 41565 8631 41599
rect 8573 41559 8631 41565
rect 6457 41531 6515 41537
rect 6457 41497 6469 41531
rect 6503 41528 6515 41531
rect 9692 41528 9720 41636
rect 10410 41624 10416 41676
rect 10468 41624 10474 41676
rect 10689 41667 10747 41673
rect 10689 41633 10701 41667
rect 10735 41664 10747 41667
rect 11716 41664 11744 41704
rect 11974 41692 11980 41704
rect 12032 41692 12038 41744
rect 12544 41732 12572 41772
rect 12618 41760 12624 41812
rect 12676 41800 12682 41812
rect 12989 41803 13047 41809
rect 12989 41800 13001 41803
rect 12676 41772 13001 41800
rect 12676 41760 12682 41772
rect 12989 41769 13001 41772
rect 13035 41769 13047 41803
rect 17954 41800 17960 41812
rect 12989 41763 13047 41769
rect 13556 41772 17960 41800
rect 12544 41704 13400 41732
rect 10735 41636 11744 41664
rect 10735 41633 10747 41636
rect 10689 41627 10747 41633
rect 11882 41624 11888 41676
rect 11940 41664 11946 41676
rect 11940 41636 13308 41664
rect 11940 41624 11946 41636
rect 9766 41556 9772 41608
rect 9824 41556 9830 41608
rect 12710 41596 12716 41608
rect 11822 41568 12716 41596
rect 12710 41556 12716 41568
rect 12768 41556 12774 41608
rect 6503 41500 9720 41528
rect 6503 41497 6515 41500
rect 6457 41491 6515 41497
rect 10594 41488 10600 41540
rect 10652 41528 10658 41540
rect 13280 41528 13308 41636
rect 13372 41596 13400 41704
rect 13449 41667 13507 41673
rect 13449 41633 13461 41667
rect 13495 41664 13507 41667
rect 13556 41664 13584 41772
rect 17954 41760 17960 41772
rect 18012 41760 18018 41812
rect 18049 41803 18107 41809
rect 18049 41769 18061 41803
rect 18095 41800 18107 41803
rect 20806 41800 20812 41812
rect 18095 41772 20812 41800
rect 18095 41769 18107 41772
rect 18049 41763 18107 41769
rect 20806 41760 20812 41772
rect 20864 41760 20870 41812
rect 20990 41760 20996 41812
rect 21048 41760 21054 41812
rect 22370 41760 22376 41812
rect 22428 41800 22434 41812
rect 24946 41800 24952 41812
rect 22428 41772 24952 41800
rect 22428 41760 22434 41772
rect 24946 41760 24952 41772
rect 25004 41760 25010 41812
rect 14274 41692 14280 41744
rect 14332 41692 14338 41744
rect 15378 41732 15384 41744
rect 14384 41704 15384 41732
rect 13495 41636 13584 41664
rect 13633 41667 13691 41673
rect 13495 41633 13507 41636
rect 13449 41627 13507 41633
rect 13633 41633 13645 41667
rect 13679 41664 13691 41667
rect 14090 41664 14096 41676
rect 13679 41636 14096 41664
rect 13679 41633 13691 41636
rect 13633 41627 13691 41633
rect 14090 41624 14096 41636
rect 14148 41624 14154 41676
rect 14384 41596 14412 41704
rect 15378 41692 15384 41704
rect 15436 41692 15442 41744
rect 17218 41692 17224 41744
rect 17276 41732 17282 41744
rect 17494 41732 17500 41744
rect 17276 41704 17500 41732
rect 17276 41692 17282 41704
rect 17494 41692 17500 41704
rect 17552 41692 17558 41744
rect 17773 41735 17831 41741
rect 17773 41701 17785 41735
rect 17819 41732 17831 41735
rect 18138 41732 18144 41744
rect 17819 41704 18144 41732
rect 17819 41701 17831 41704
rect 17773 41695 17831 41701
rect 18138 41692 18144 41704
rect 18196 41692 18202 41744
rect 22646 41732 22652 41744
rect 18708 41704 22652 41732
rect 14734 41624 14740 41676
rect 14792 41624 14798 41676
rect 14921 41667 14979 41673
rect 14921 41633 14933 41667
rect 14967 41664 14979 41667
rect 15746 41664 15752 41676
rect 14967 41636 15752 41664
rect 14967 41633 14979 41636
rect 14921 41627 14979 41633
rect 15746 41624 15752 41636
rect 15804 41624 15810 41676
rect 18230 41624 18236 41676
rect 18288 41664 18294 41676
rect 18708 41673 18736 41704
rect 22646 41692 22652 41704
rect 22704 41692 22710 41744
rect 24854 41732 24860 41744
rect 23492 41704 24860 41732
rect 18509 41667 18567 41673
rect 18509 41664 18521 41667
rect 18288 41636 18521 41664
rect 18288 41624 18294 41636
rect 18509 41633 18521 41636
rect 18555 41633 18567 41667
rect 18509 41627 18567 41633
rect 18693 41667 18751 41673
rect 18693 41633 18705 41667
rect 18739 41633 18751 41667
rect 21545 41667 21603 41673
rect 21545 41664 21557 41667
rect 18693 41627 18751 41633
rect 19168 41636 21557 41664
rect 13372 41568 14412 41596
rect 14550 41556 14556 41608
rect 14608 41596 14614 41608
rect 15473 41599 15531 41605
rect 15473 41596 15485 41599
rect 14608 41568 15485 41596
rect 14608 41556 14614 41568
rect 15473 41565 15485 41568
rect 15519 41565 15531 41599
rect 15473 41559 15531 41565
rect 17957 41599 18015 41605
rect 17957 41565 17969 41599
rect 18003 41596 18015 41599
rect 18322 41596 18328 41608
rect 18003 41568 18328 41596
rect 18003 41565 18015 41568
rect 17957 41559 18015 41565
rect 18322 41556 18328 41568
rect 18380 41556 18386 41608
rect 18417 41599 18475 41605
rect 18417 41565 18429 41599
rect 18463 41596 18475 41599
rect 19061 41599 19119 41605
rect 19061 41596 19073 41599
rect 18463 41592 18644 41596
rect 18708 41592 19073 41596
rect 18463 41568 19073 41592
rect 18463 41565 18475 41568
rect 18417 41559 18475 41565
rect 18616 41564 18736 41568
rect 19061 41565 19073 41568
rect 19107 41565 19119 41599
rect 19061 41559 19119 41565
rect 14645 41531 14703 41537
rect 14645 41528 14657 41531
rect 10652 41500 10916 41528
rect 10652 41488 10658 41500
rect 5534 41420 5540 41472
rect 5592 41460 5598 41472
rect 6549 41463 6607 41469
rect 6549 41460 6561 41463
rect 5592 41432 6561 41460
rect 5592 41420 5598 41432
rect 6549 41429 6561 41432
rect 6595 41429 6607 41463
rect 10888 41460 10916 41500
rect 11992 41500 12434 41528
rect 13280 41500 14657 41528
rect 11992 41460 12020 41500
rect 10888 41432 12020 41460
rect 12161 41463 12219 41469
rect 6549 41423 6607 41429
rect 12161 41429 12173 41463
rect 12207 41460 12219 41463
rect 12250 41460 12256 41472
rect 12207 41432 12256 41460
rect 12207 41429 12219 41432
rect 12161 41423 12219 41429
rect 12250 41420 12256 41432
rect 12308 41420 12314 41472
rect 12406 41460 12434 41500
rect 14645 41497 14657 41500
rect 14691 41497 14703 41531
rect 19168 41528 19196 41636
rect 21545 41633 21557 41636
rect 21591 41633 21603 41667
rect 21545 41627 21603 41633
rect 22094 41624 22100 41676
rect 22152 41664 22158 41676
rect 22557 41667 22615 41673
rect 22557 41664 22569 41667
rect 22152 41636 22569 41664
rect 22152 41624 22158 41636
rect 22557 41633 22569 41636
rect 22603 41633 22615 41667
rect 22557 41627 22615 41633
rect 20165 41599 20223 41605
rect 20165 41565 20177 41599
rect 20211 41596 20223 41599
rect 20714 41596 20720 41608
rect 20211 41568 20720 41596
rect 20211 41565 20223 41568
rect 20165 41559 20223 41565
rect 20714 41556 20720 41568
rect 20772 41556 20778 41608
rect 20901 41599 20959 41605
rect 20901 41565 20913 41599
rect 20947 41596 20959 41599
rect 20990 41596 20996 41608
rect 20947 41568 20996 41596
rect 20947 41565 20959 41568
rect 20901 41559 20959 41565
rect 20990 41556 20996 41568
rect 21048 41556 21054 41608
rect 23492 41596 23520 41704
rect 24854 41692 24860 41704
rect 24912 41692 24918 41744
rect 23566 41624 23572 41676
rect 23624 41664 23630 41676
rect 23842 41664 23848 41676
rect 23624 41636 23848 41664
rect 23624 41624 23630 41636
rect 23842 41624 23848 41636
rect 23900 41624 23906 41676
rect 21376 41568 23520 41596
rect 14645 41491 14703 41497
rect 15948 41500 16238 41528
rect 17052 41500 19196 41528
rect 15948 41472 15976 41500
rect 13357 41463 13415 41469
rect 13357 41460 13369 41463
rect 12406 41432 13369 41460
rect 13357 41429 13369 41432
rect 13403 41429 13415 41463
rect 13357 41423 13415 41429
rect 15930 41420 15936 41472
rect 15988 41420 15994 41472
rect 16114 41420 16120 41472
rect 16172 41460 16178 41472
rect 17052 41460 17080 41500
rect 21376 41472 21404 41568
rect 23658 41556 23664 41608
rect 23716 41556 23722 41608
rect 21453 41531 21511 41537
rect 21453 41497 21465 41531
rect 21499 41528 21511 41531
rect 22186 41528 22192 41540
rect 21499 41500 22192 41528
rect 21499 41497 21511 41500
rect 21453 41491 21511 41497
rect 22186 41488 22192 41500
rect 22244 41488 22250 41540
rect 22373 41531 22431 41537
rect 22373 41497 22385 41531
rect 22419 41528 22431 41531
rect 24486 41528 24492 41540
rect 22419 41500 24492 41528
rect 22419 41497 22431 41500
rect 22373 41491 22431 41497
rect 24486 41488 24492 41500
rect 24544 41488 24550 41540
rect 16172 41432 17080 41460
rect 16172 41420 16178 41432
rect 17494 41420 17500 41472
rect 17552 41460 17558 41472
rect 20346 41460 20352 41472
rect 17552 41432 20352 41460
rect 17552 41420 17558 41432
rect 20346 41420 20352 41432
rect 20404 41420 20410 41472
rect 20898 41420 20904 41472
rect 20956 41460 20962 41472
rect 21266 41460 21272 41472
rect 20956 41432 21272 41460
rect 20956 41420 20962 41432
rect 21266 41420 21272 41432
rect 21324 41420 21330 41472
rect 21358 41420 21364 41472
rect 21416 41420 21422 41472
rect 21634 41420 21640 41472
rect 21692 41460 21698 41472
rect 22005 41463 22063 41469
rect 22005 41460 22017 41463
rect 21692 41432 22017 41460
rect 21692 41420 21698 41432
rect 22005 41429 22017 41432
rect 22051 41429 22063 41463
rect 22005 41423 22063 41429
rect 22465 41463 22523 41469
rect 22465 41429 22477 41463
rect 22511 41460 22523 41463
rect 23293 41463 23351 41469
rect 23293 41460 23305 41463
rect 22511 41432 23305 41460
rect 22511 41429 22523 41432
rect 22465 41423 22523 41429
rect 23293 41429 23305 41432
rect 23339 41429 23351 41463
rect 23293 41423 23351 41429
rect 23750 41420 23756 41472
rect 23808 41460 23814 41472
rect 27246 41460 27252 41472
rect 23808 41432 27252 41460
rect 23808 41420 23814 41432
rect 27246 41420 27252 41432
rect 27304 41420 27310 41472
rect 1104 41370 49864 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 27950 41370
rect 28002 41318 28014 41370
rect 28066 41318 28078 41370
rect 28130 41318 28142 41370
rect 28194 41318 28206 41370
rect 28258 41318 37950 41370
rect 38002 41318 38014 41370
rect 38066 41318 38078 41370
rect 38130 41318 38142 41370
rect 38194 41318 38206 41370
rect 38258 41318 47950 41370
rect 48002 41318 48014 41370
rect 48066 41318 48078 41370
rect 48130 41318 48142 41370
rect 48194 41318 48206 41370
rect 48258 41318 49864 41370
rect 1104 41296 49864 41318
rect 10318 41256 10324 41268
rect 6748 41228 10324 41256
rect 6748 41197 6776 41228
rect 10318 41216 10324 41228
rect 10376 41216 10382 41268
rect 11514 41216 11520 41268
rect 11572 41256 11578 41268
rect 12066 41256 12072 41268
rect 11572 41228 12072 41256
rect 11572 41216 11578 41228
rect 12066 41216 12072 41228
rect 12124 41216 12130 41268
rect 14550 41256 14556 41268
rect 12360 41228 14556 41256
rect 6733 41191 6791 41197
rect 6733 41157 6745 41191
rect 6779 41157 6791 41191
rect 9214 41188 9220 41200
rect 6733 41151 6791 41157
rect 6840 41160 9220 41188
rect 1765 41123 1823 41129
rect 1765 41089 1777 41123
rect 1811 41120 1823 41123
rect 6840 41120 6868 41160
rect 9214 41148 9220 41160
rect 9272 41148 9278 41200
rect 11330 41188 11336 41200
rect 10902 41160 11336 41188
rect 11330 41148 11336 41160
rect 11388 41148 11394 41200
rect 1811 41092 6868 41120
rect 1811 41089 1823 41092
rect 1765 41083 1823 41089
rect 7834 41080 7840 41132
rect 7892 41120 7898 41132
rect 8021 41123 8079 41129
rect 8021 41120 8033 41123
rect 7892 41092 8033 41120
rect 7892 41080 7898 41092
rect 8021 41089 8033 41092
rect 8067 41089 8079 41123
rect 8021 41083 8079 41089
rect 8478 41080 8484 41132
rect 8536 41120 8542 41132
rect 9401 41123 9459 41129
rect 9401 41120 9413 41123
rect 8536 41092 9413 41120
rect 8536 41080 8542 41092
rect 9401 41089 9413 41092
rect 9447 41089 9459 41123
rect 9401 41083 9459 41089
rect 11698 41080 11704 41132
rect 11756 41120 11762 41132
rect 12360 41129 12388 41228
rect 14550 41216 14556 41228
rect 14608 41216 14614 41268
rect 15746 41216 15752 41268
rect 15804 41256 15810 41268
rect 16301 41259 16359 41265
rect 16301 41256 16313 41259
rect 15804 41228 16313 41256
rect 15804 41216 15810 41228
rect 16301 41225 16313 41228
rect 16347 41225 16359 41259
rect 16301 41219 16359 41225
rect 16482 41216 16488 41268
rect 16540 41256 16546 41268
rect 16853 41259 16911 41265
rect 16853 41256 16865 41259
rect 16540 41228 16865 41256
rect 16540 41216 16546 41228
rect 16853 41225 16865 41228
rect 16899 41225 16911 41259
rect 16853 41219 16911 41225
rect 19242 41216 19248 41268
rect 19300 41216 19306 41268
rect 19613 41259 19671 41265
rect 19613 41225 19625 41259
rect 19659 41256 19671 41259
rect 20533 41259 20591 41265
rect 20533 41256 20545 41259
rect 19659 41228 20545 41256
rect 19659 41225 19671 41228
rect 19613 41219 19671 41225
rect 20533 41225 20545 41228
rect 20579 41256 20591 41259
rect 24394 41256 24400 41268
rect 20579 41228 24400 41256
rect 20579 41225 20591 41228
rect 20533 41219 20591 41225
rect 24394 41216 24400 41228
rect 24452 41216 24458 41268
rect 24486 41216 24492 41268
rect 24544 41216 24550 41268
rect 24854 41216 24860 41268
rect 24912 41216 24918 41268
rect 24946 41216 24952 41268
rect 25004 41216 25010 41268
rect 46106 41256 46112 41268
rect 31726 41228 46112 41256
rect 12710 41148 12716 41200
rect 12768 41188 12774 41200
rect 12768 41160 13110 41188
rect 12768 41148 12774 41160
rect 14568 41129 14596 41216
rect 19518 41188 19524 41200
rect 17420 41160 19524 41188
rect 12345 41123 12403 41129
rect 12345 41120 12357 41123
rect 11756 41092 12357 41120
rect 11756 41080 11762 41092
rect 12345 41089 12357 41092
rect 12391 41089 12403 41123
rect 12345 41083 12403 41089
rect 14553 41123 14611 41129
rect 14553 41089 14565 41123
rect 14599 41089 14611 41123
rect 14553 41083 14611 41089
rect 15930 41080 15936 41132
rect 15988 41080 15994 41132
rect 16482 41080 16488 41132
rect 16540 41120 16546 41132
rect 17221 41123 17279 41129
rect 17221 41120 17233 41123
rect 16540 41092 17233 41120
rect 16540 41080 16546 41092
rect 17221 41089 17233 41092
rect 17267 41089 17279 41123
rect 17221 41083 17279 41089
rect 1302 41012 1308 41064
rect 1360 41052 1366 41064
rect 2041 41055 2099 41061
rect 2041 41052 2053 41055
rect 1360 41024 2053 41052
rect 1360 41012 1366 41024
rect 2041 41021 2053 41024
rect 2087 41021 2099 41055
rect 2041 41015 2099 41021
rect 8570 41012 8576 41064
rect 8628 41052 8634 41064
rect 8757 41055 8815 41061
rect 8757 41052 8769 41055
rect 8628 41024 8769 41052
rect 8628 41012 8634 41024
rect 8757 41021 8769 41024
rect 8803 41021 8815 41055
rect 8757 41015 8815 41021
rect 9677 41055 9735 41061
rect 9677 41021 9689 41055
rect 9723 41052 9735 41055
rect 12250 41052 12256 41064
rect 9723 41024 12256 41052
rect 9723 41021 9735 41024
rect 9677 41015 9735 41021
rect 12250 41012 12256 41024
rect 12308 41012 12314 41064
rect 12621 41055 12679 41061
rect 12621 41052 12633 41055
rect 12406 41024 12633 41052
rect 6914 40944 6920 40996
rect 6972 40944 6978 40996
rect 11330 40944 11336 40996
rect 11388 40984 11394 40996
rect 12406 40984 12434 41024
rect 12621 41021 12633 41024
rect 12667 41052 12679 41055
rect 13630 41052 13636 41064
rect 12667 41024 13636 41052
rect 12667 41021 12679 41024
rect 12621 41015 12679 41021
rect 13630 41012 13636 41024
rect 13688 41012 13694 41064
rect 14090 41012 14096 41064
rect 14148 41012 14154 41064
rect 14182 41012 14188 41064
rect 14240 41052 14246 41064
rect 14829 41055 14887 41061
rect 14829 41052 14841 41055
rect 14240 41024 14841 41052
rect 14240 41012 14246 41024
rect 14829 41021 14841 41024
rect 14875 41021 14887 41055
rect 14829 41015 14887 41021
rect 16298 41012 16304 41064
rect 16356 41052 16362 41064
rect 17313 41055 17371 41061
rect 17313 41052 17325 41055
rect 16356 41024 17325 41052
rect 16356 41012 16362 41024
rect 17313 41021 17325 41024
rect 17359 41021 17371 41055
rect 17313 41015 17371 41021
rect 11388 40956 12434 40984
rect 11388 40944 11394 40956
rect 8202 40876 8208 40928
rect 8260 40916 8266 40928
rect 10686 40916 10692 40928
rect 8260 40888 10692 40916
rect 8260 40876 8266 40888
rect 10686 40876 10692 40888
rect 10744 40876 10750 40928
rect 10870 40876 10876 40928
rect 10928 40916 10934 40928
rect 11149 40919 11207 40925
rect 11149 40916 11161 40919
rect 10928 40888 11161 40916
rect 10928 40876 10934 40888
rect 11149 40885 11161 40888
rect 11195 40885 11207 40919
rect 11149 40879 11207 40885
rect 11882 40876 11888 40928
rect 11940 40876 11946 40928
rect 13630 40876 13636 40928
rect 13688 40916 13694 40928
rect 17420 40916 17448 41160
rect 19518 41148 19524 41160
rect 19576 41148 19582 41200
rect 22186 41148 22192 41200
rect 22244 41188 22250 41200
rect 23198 41188 23204 41200
rect 22244 41160 23204 41188
rect 22244 41148 22250 41160
rect 23198 41148 23204 41160
rect 23256 41188 23262 41200
rect 23477 41191 23535 41197
rect 23477 41188 23489 41191
rect 23256 41160 23489 41188
rect 23256 41148 23262 41160
rect 23477 41157 23489 41160
rect 23523 41157 23535 41191
rect 23477 41151 23535 41157
rect 23569 41191 23627 41197
rect 23569 41157 23581 41191
rect 23615 41188 23627 41191
rect 31726 41188 31754 41228
rect 46106 41216 46112 41228
rect 46164 41216 46170 41268
rect 23615 41160 31754 41188
rect 23615 41157 23627 41160
rect 23569 41151 23627 41157
rect 19705 41123 19763 41129
rect 19705 41120 19717 41123
rect 18708 41092 19717 41120
rect 17497 41055 17555 41061
rect 17497 41021 17509 41055
rect 17543 41052 17555 41055
rect 17862 41052 17868 41064
rect 17543 41024 17868 41052
rect 17543 41021 17555 41024
rect 17497 41015 17555 41021
rect 17862 41012 17868 41024
rect 17920 41012 17926 41064
rect 13688 40888 17448 40916
rect 13688 40876 13694 40888
rect 17494 40876 17500 40928
rect 17552 40916 17558 40928
rect 18708 40925 18736 41092
rect 19705 41089 19717 41092
rect 19751 41089 19763 41123
rect 19705 41083 19763 41089
rect 22649 41123 22707 41129
rect 22649 41089 22661 41123
rect 22695 41120 22707 41123
rect 23382 41120 23388 41132
rect 22695 41092 23388 41120
rect 22695 41089 22707 41092
rect 22649 41083 22707 41089
rect 23382 41080 23388 41092
rect 23440 41120 23446 41132
rect 23584 41120 23612 41151
rect 23934 41120 23940 41132
rect 23440 41092 23612 41120
rect 23676 41092 23940 41120
rect 23440 41080 23446 41092
rect 18782 41012 18788 41064
rect 18840 41052 18846 41064
rect 19610 41052 19616 41064
rect 18840 41024 19616 41052
rect 18840 41012 18846 41024
rect 19610 41012 19616 41024
rect 19668 41012 19674 41064
rect 23676 41061 23704 41092
rect 23934 41080 23940 41092
rect 23992 41080 23998 41132
rect 47762 41120 47768 41132
rect 31726 41092 47768 41120
rect 19889 41055 19947 41061
rect 19889 41021 19901 41055
rect 19935 41021 19947 41055
rect 19889 41015 19947 41021
rect 23661 41055 23719 41061
rect 23661 41021 23673 41055
rect 23707 41021 23719 41055
rect 23661 41015 23719 41021
rect 19518 40944 19524 40996
rect 19576 40984 19582 40996
rect 19904 40984 19932 41015
rect 23842 41012 23848 41064
rect 23900 41052 23906 41064
rect 25041 41055 25099 41061
rect 25041 41052 25053 41055
rect 23900 41024 25053 41052
rect 23900 41012 23906 41024
rect 25041 41021 25053 41024
rect 25087 41021 25099 41055
rect 25041 41015 25099 41021
rect 23474 40984 23480 40996
rect 19576 40956 19932 40984
rect 22066 40956 23480 40984
rect 19576 40944 19582 40956
rect 18693 40919 18751 40925
rect 18693 40916 18705 40919
rect 17552 40888 18705 40916
rect 17552 40876 17558 40888
rect 18693 40885 18705 40888
rect 18739 40916 18751 40919
rect 22066 40916 22094 40956
rect 23474 40944 23480 40956
rect 23532 40944 23538 40996
rect 18739 40888 22094 40916
rect 18739 40885 18751 40888
rect 18693 40879 18751 40885
rect 22646 40876 22652 40928
rect 22704 40916 22710 40928
rect 23109 40919 23167 40925
rect 23109 40916 23121 40919
rect 22704 40888 23121 40916
rect 22704 40876 22710 40888
rect 23109 40885 23121 40888
rect 23155 40885 23167 40919
rect 23109 40879 23167 40885
rect 23198 40876 23204 40928
rect 23256 40916 23262 40928
rect 24397 40919 24455 40925
rect 24397 40916 24409 40919
rect 23256 40888 24409 40916
rect 23256 40876 23262 40888
rect 24397 40885 24409 40888
rect 24443 40916 24455 40919
rect 31726 40916 31754 41092
rect 47762 41080 47768 41092
rect 47820 41080 47826 41132
rect 24443 40888 31754 40916
rect 24443 40885 24455 40888
rect 24397 40879 24455 40885
rect 1104 40826 49864 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 32950 40826
rect 33002 40774 33014 40826
rect 33066 40774 33078 40826
rect 33130 40774 33142 40826
rect 33194 40774 33206 40826
rect 33258 40774 42950 40826
rect 43002 40774 43014 40826
rect 43066 40774 43078 40826
rect 43130 40774 43142 40826
rect 43194 40774 43206 40826
rect 43258 40774 49864 40826
rect 1104 40752 49864 40774
rect 7742 40672 7748 40724
rect 7800 40712 7806 40724
rect 7837 40715 7895 40721
rect 7837 40712 7849 40715
rect 7800 40684 7849 40712
rect 7800 40672 7806 40684
rect 7837 40681 7849 40684
rect 7883 40681 7895 40715
rect 7837 40675 7895 40681
rect 9122 40672 9128 40724
rect 9180 40672 9186 40724
rect 10686 40672 10692 40724
rect 10744 40712 10750 40724
rect 10744 40684 11560 40712
rect 10744 40672 10750 40684
rect 7377 40647 7435 40653
rect 7377 40613 7389 40647
rect 7423 40644 7435 40647
rect 11532 40644 11560 40684
rect 11974 40672 11980 40724
rect 12032 40672 12038 40724
rect 12526 40672 12532 40724
rect 12584 40712 12590 40724
rect 12989 40715 13047 40721
rect 12989 40712 13001 40715
rect 12584 40684 13001 40712
rect 12584 40672 12590 40684
rect 12989 40681 13001 40684
rect 13035 40681 13047 40715
rect 17116 40715 17174 40721
rect 12989 40675 13047 40681
rect 14200 40684 16574 40712
rect 7423 40616 10364 40644
rect 11532 40616 12848 40644
rect 7423 40613 7435 40616
rect 7377 40607 7435 40613
rect 8389 40579 8447 40585
rect 8389 40545 8401 40579
rect 8435 40576 8447 40579
rect 9030 40576 9036 40588
rect 8435 40548 9036 40576
rect 8435 40545 8447 40548
rect 8389 40539 8447 40545
rect 9030 40536 9036 40548
rect 9088 40536 9094 40588
rect 9306 40536 9312 40588
rect 9364 40576 9370 40588
rect 9677 40579 9735 40585
rect 9677 40576 9689 40579
rect 9364 40548 9689 40576
rect 9364 40536 9370 40548
rect 9677 40545 9689 40548
rect 9723 40545 9735 40579
rect 10336 40576 10364 40616
rect 10336 40548 11744 40576
rect 9677 40539 9735 40545
rect 8205 40511 8263 40517
rect 8205 40477 8217 40511
rect 8251 40508 8263 40511
rect 8294 40508 8300 40520
rect 8251 40480 8300 40508
rect 8251 40477 8263 40480
rect 8205 40471 8263 40477
rect 8294 40468 8300 40480
rect 8352 40468 8358 40520
rect 8478 40468 8484 40520
rect 8536 40508 8542 40520
rect 10229 40511 10287 40517
rect 10229 40508 10241 40511
rect 8536 40480 10241 40508
rect 8536 40468 8542 40480
rect 10229 40477 10241 40480
rect 10275 40477 10287 40511
rect 11716 40508 11744 40548
rect 12710 40508 12716 40520
rect 11716 40480 12716 40508
rect 10229 40471 10287 40477
rect 8754 40400 8760 40452
rect 8812 40440 8818 40452
rect 9585 40443 9643 40449
rect 9585 40440 9597 40443
rect 8812 40412 9597 40440
rect 8812 40400 8818 40412
rect 9585 40409 9597 40412
rect 9631 40409 9643 40443
rect 10244 40440 10272 40471
rect 12710 40468 12716 40480
rect 12768 40468 12774 40520
rect 12820 40508 12848 40616
rect 12986 40536 12992 40588
rect 13044 40576 13050 40588
rect 13541 40579 13599 40585
rect 13541 40576 13553 40579
rect 13044 40548 13553 40576
rect 13044 40536 13050 40548
rect 13541 40545 13553 40548
rect 13587 40545 13599 40579
rect 13541 40539 13599 40545
rect 13357 40511 13415 40517
rect 13357 40508 13369 40511
rect 12820 40480 13369 40508
rect 13357 40477 13369 40480
rect 13403 40477 13415 40511
rect 13357 40471 13415 40477
rect 13449 40511 13507 40517
rect 13449 40477 13461 40511
rect 13495 40508 13507 40511
rect 14200 40508 14228 40684
rect 14277 40579 14335 40585
rect 14277 40545 14289 40579
rect 14323 40576 14335 40579
rect 14550 40576 14556 40588
rect 14323 40548 14556 40576
rect 14323 40545 14335 40548
rect 14277 40539 14335 40545
rect 14550 40536 14556 40548
rect 14608 40536 14614 40588
rect 13495 40480 14228 40508
rect 13495 40477 13507 40480
rect 13449 40471 13507 40477
rect 10410 40440 10416 40452
rect 10244 40412 10416 40440
rect 9585 40403 9643 40409
rect 10410 40400 10416 40412
rect 10468 40400 10474 40452
rect 10505 40443 10563 40449
rect 10505 40409 10517 40443
rect 10551 40409 10563 40443
rect 10505 40403 10563 40409
rect 7742 40332 7748 40384
rect 7800 40372 7806 40384
rect 8297 40375 8355 40381
rect 8297 40372 8309 40375
rect 7800 40344 8309 40372
rect 7800 40332 7806 40344
rect 8297 40341 8309 40344
rect 8343 40341 8355 40375
rect 8297 40335 8355 40341
rect 8386 40332 8392 40384
rect 8444 40372 8450 40384
rect 9493 40375 9551 40381
rect 9493 40372 9505 40375
rect 8444 40344 9505 40372
rect 8444 40332 8450 40344
rect 9493 40341 9505 40344
rect 9539 40341 9551 40375
rect 10520 40372 10548 40403
rect 11238 40400 11244 40452
rect 11296 40400 11302 40452
rect 13262 40440 13268 40452
rect 12406 40412 13268 40440
rect 12406 40372 12434 40412
rect 13262 40400 13268 40412
rect 13320 40400 13326 40452
rect 10520 40344 12434 40372
rect 12529 40375 12587 40381
rect 9493 40335 9551 40341
rect 12529 40341 12541 40375
rect 12575 40372 12587 40375
rect 13464 40372 13492 40471
rect 14090 40400 14096 40452
rect 14148 40440 14154 40452
rect 14553 40443 14611 40449
rect 14553 40440 14565 40443
rect 14148 40412 14565 40440
rect 14148 40400 14154 40412
rect 14553 40409 14565 40412
rect 14599 40409 14611 40443
rect 15930 40440 15936 40452
rect 15778 40412 15936 40440
rect 14553 40403 14611 40409
rect 15930 40400 15936 40412
rect 15988 40400 15994 40452
rect 12575 40344 13492 40372
rect 12575 40341 12587 40344
rect 12529 40335 12587 40341
rect 14182 40332 14188 40384
rect 14240 40372 14246 40384
rect 16025 40375 16083 40381
rect 16025 40372 16037 40375
rect 14240 40344 16037 40372
rect 14240 40332 14246 40344
rect 16025 40341 16037 40344
rect 16071 40372 16083 40375
rect 16114 40372 16120 40384
rect 16071 40344 16120 40372
rect 16071 40341 16083 40344
rect 16025 40335 16083 40341
rect 16114 40332 16120 40344
rect 16172 40332 16178 40384
rect 16546 40372 16574 40684
rect 17116 40681 17128 40715
rect 17162 40712 17174 40715
rect 19978 40712 19984 40724
rect 17162 40684 19984 40712
rect 17162 40681 17174 40684
rect 17116 40675 17174 40681
rect 19978 40672 19984 40684
rect 20036 40672 20042 40724
rect 20622 40672 20628 40724
rect 20680 40712 20686 40724
rect 23658 40712 23664 40724
rect 20680 40684 23664 40712
rect 20680 40672 20686 40684
rect 23658 40672 23664 40684
rect 23716 40672 23722 40724
rect 24394 40672 24400 40724
rect 24452 40712 24458 40724
rect 49050 40712 49056 40724
rect 24452 40684 49056 40712
rect 24452 40672 24458 40684
rect 49050 40672 49056 40684
rect 49108 40672 49114 40724
rect 19058 40604 19064 40656
rect 19116 40644 19122 40656
rect 19116 40616 20944 40644
rect 19116 40604 19122 40616
rect 16853 40579 16911 40585
rect 16853 40545 16865 40579
rect 16899 40576 16911 40579
rect 19702 40576 19708 40588
rect 16899 40548 19708 40576
rect 16899 40545 16911 40548
rect 16853 40539 16911 40545
rect 19702 40536 19708 40548
rect 19760 40536 19766 40588
rect 20916 40585 20944 40616
rect 20901 40579 20959 40585
rect 20901 40545 20913 40579
rect 20947 40545 20959 40579
rect 20901 40539 20959 40545
rect 21818 40536 21824 40588
rect 21876 40536 21882 40588
rect 24762 40536 24768 40588
rect 24820 40576 24826 40588
rect 25133 40579 25191 40585
rect 25133 40576 25145 40579
rect 24820 40548 25145 40576
rect 24820 40536 24826 40548
rect 25133 40545 25145 40548
rect 25179 40545 25191 40579
rect 25133 40539 25191 40545
rect 19150 40508 19156 40520
rect 18262 40480 19156 40508
rect 19150 40468 19156 40480
rect 19208 40468 19214 40520
rect 19720 40508 19748 40536
rect 21542 40508 21548 40520
rect 19720 40480 21548 40508
rect 21542 40468 21548 40480
rect 21600 40468 21606 40520
rect 23750 40468 23756 40520
rect 23808 40508 23814 40520
rect 23845 40511 23903 40517
rect 23845 40508 23857 40511
rect 23808 40480 23857 40508
rect 23808 40468 23814 40480
rect 23845 40477 23857 40480
rect 23891 40508 23903 40511
rect 25041 40511 25099 40517
rect 25041 40508 25053 40511
rect 23891 40480 25053 40508
rect 23891 40477 23903 40480
rect 23845 40471 23903 40477
rect 25041 40477 25053 40480
rect 25087 40508 25099 40511
rect 25087 40480 31754 40508
rect 25087 40477 25099 40480
rect 25041 40471 25099 40477
rect 18874 40400 18880 40452
rect 18932 40400 18938 40452
rect 20717 40443 20775 40449
rect 19812 40412 20484 40440
rect 19812 40384 19840 40412
rect 18782 40372 18788 40384
rect 16546 40344 18788 40372
rect 18782 40332 18788 40344
rect 18840 40332 18846 40384
rect 19794 40332 19800 40384
rect 19852 40332 19858 40384
rect 20346 40332 20352 40384
rect 20404 40332 20410 40384
rect 20456 40372 20484 40412
rect 20717 40409 20729 40443
rect 20763 40440 20775 40443
rect 20898 40440 20904 40452
rect 20763 40412 20904 40440
rect 20763 40409 20775 40412
rect 20717 40403 20775 40409
rect 20898 40400 20904 40412
rect 20956 40400 20962 40452
rect 21266 40400 21272 40452
rect 21324 40440 21330 40452
rect 22278 40440 22284 40452
rect 21324 40412 22284 40440
rect 21324 40400 21330 40412
rect 22278 40400 22284 40412
rect 22336 40400 22342 40452
rect 23474 40400 23480 40452
rect 23532 40440 23538 40452
rect 23658 40440 23664 40452
rect 23532 40412 23664 40440
rect 23532 40400 23538 40412
rect 23658 40400 23664 40412
rect 23716 40440 23722 40452
rect 24949 40443 25007 40449
rect 24949 40440 24961 40443
rect 23716 40412 24961 40440
rect 23716 40400 23722 40412
rect 24949 40409 24961 40412
rect 24995 40409 25007 40443
rect 31726 40440 31754 40480
rect 45278 40440 45284 40452
rect 31726 40412 45284 40440
rect 24949 40403 25007 40409
rect 20622 40372 20628 40384
rect 20456 40344 20628 40372
rect 20622 40332 20628 40344
rect 20680 40372 20686 40384
rect 20809 40375 20867 40381
rect 20809 40372 20821 40375
rect 20680 40344 20821 40372
rect 20680 40332 20686 40344
rect 20809 40341 20821 40344
rect 20855 40341 20867 40375
rect 20916 40372 20944 40400
rect 22830 40372 22836 40384
rect 20916 40344 22836 40372
rect 20809 40335 20867 40341
rect 22830 40332 22836 40344
rect 22888 40332 22894 40384
rect 23290 40332 23296 40384
rect 23348 40332 23354 40384
rect 24578 40332 24584 40384
rect 24636 40332 24642 40384
rect 24964 40372 24992 40403
rect 45278 40400 45284 40412
rect 45336 40400 45342 40452
rect 25869 40375 25927 40381
rect 25869 40372 25881 40375
rect 24964 40344 25881 40372
rect 25869 40341 25881 40344
rect 25915 40372 25927 40375
rect 46934 40372 46940 40384
rect 25915 40344 46940 40372
rect 25915 40341 25927 40344
rect 25869 40335 25927 40341
rect 46934 40332 46940 40344
rect 46992 40332 46998 40384
rect 1104 40282 49864 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 27950 40282
rect 28002 40230 28014 40282
rect 28066 40230 28078 40282
rect 28130 40230 28142 40282
rect 28194 40230 28206 40282
rect 28258 40230 37950 40282
rect 38002 40230 38014 40282
rect 38066 40230 38078 40282
rect 38130 40230 38142 40282
rect 38194 40230 38206 40282
rect 38258 40230 47950 40282
rect 48002 40230 48014 40282
rect 48066 40230 48078 40282
rect 48130 40230 48142 40282
rect 48194 40230 48206 40282
rect 48258 40230 49864 40282
rect 1104 40208 49864 40230
rect 8846 40128 8852 40180
rect 8904 40168 8910 40180
rect 10229 40171 10287 40177
rect 10229 40168 10241 40171
rect 8904 40140 10241 40168
rect 8904 40128 8910 40140
rect 10229 40137 10241 40140
rect 10275 40137 10287 40171
rect 11238 40168 11244 40180
rect 10229 40131 10287 40137
rect 10888 40140 11244 40168
rect 4338 40100 4344 40112
rect 1780 40072 4344 40100
rect 1780 40041 1808 40072
rect 4338 40060 4344 40072
rect 4396 40060 4402 40112
rect 7837 40103 7895 40109
rect 7837 40069 7849 40103
rect 7883 40100 7895 40103
rect 8294 40100 8300 40112
rect 7883 40072 8300 40100
rect 7883 40069 7895 40072
rect 7837 40063 7895 40069
rect 8294 40060 8300 40072
rect 8352 40060 8358 40112
rect 10134 40100 10140 40112
rect 9982 40072 10140 40100
rect 10134 40060 10140 40072
rect 10192 40100 10198 40112
rect 10888 40100 10916 40140
rect 11238 40128 11244 40140
rect 11296 40168 11302 40180
rect 11296 40140 12204 40168
rect 11296 40128 11302 40140
rect 10192 40072 10916 40100
rect 10965 40103 11023 40109
rect 10192 40060 10198 40072
rect 10965 40069 10977 40103
rect 11011 40100 11023 40103
rect 12066 40100 12072 40112
rect 11011 40072 12072 40100
rect 11011 40069 11023 40072
rect 10965 40063 11023 40069
rect 12066 40060 12072 40072
rect 12124 40060 12130 40112
rect 12176 40100 12204 40140
rect 12342 40128 12348 40180
rect 12400 40168 12406 40180
rect 17402 40168 17408 40180
rect 12400 40140 17408 40168
rect 12400 40128 12406 40140
rect 17402 40128 17408 40140
rect 17460 40168 17466 40180
rect 20714 40168 20720 40180
rect 17460 40140 20720 40168
rect 17460 40128 17466 40140
rect 15473 40103 15531 40109
rect 12176 40072 12466 40100
rect 15473 40069 15485 40103
rect 15519 40100 15531 40103
rect 17034 40100 17040 40112
rect 15519 40072 17040 40100
rect 15519 40069 15531 40072
rect 15473 40063 15531 40069
rect 17034 40060 17040 40072
rect 17092 40060 17098 40112
rect 17604 40109 17632 40140
rect 20714 40128 20720 40140
rect 20772 40168 20778 40180
rect 20772 40140 22048 40168
rect 20772 40128 20778 40140
rect 17589 40103 17647 40109
rect 17589 40069 17601 40103
rect 17635 40069 17647 40103
rect 17589 40063 17647 40069
rect 18322 40060 18328 40112
rect 18380 40100 18386 40112
rect 18506 40100 18512 40112
rect 18380 40072 18512 40100
rect 18380 40060 18386 40072
rect 18506 40060 18512 40072
rect 18564 40060 18570 40112
rect 19058 40100 19064 40112
rect 18892 40072 19064 40100
rect 1765 40035 1823 40041
rect 1765 40001 1777 40035
rect 1811 40001 1823 40035
rect 1765 39995 1823 40001
rect 8478 39992 8484 40044
rect 8536 39992 8542 40044
rect 11698 39992 11704 40044
rect 11756 39992 11762 40044
rect 13814 40032 13820 40044
rect 13188 40004 13820 40032
rect 2038 39924 2044 39976
rect 2096 39924 2102 39976
rect 7285 39967 7343 39973
rect 7285 39933 7297 39967
rect 7331 39964 7343 39967
rect 8386 39964 8392 39976
rect 7331 39936 8392 39964
rect 7331 39933 7343 39936
rect 7285 39927 7343 39933
rect 8386 39924 8392 39936
rect 8444 39924 8450 39976
rect 8757 39967 8815 39973
rect 8757 39933 8769 39967
rect 8803 39964 8815 39967
rect 10870 39964 10876 39976
rect 8803 39936 10876 39964
rect 8803 39933 8815 39936
rect 8757 39927 8815 39933
rect 10870 39924 10876 39936
rect 10928 39924 10934 39976
rect 11514 39924 11520 39976
rect 11572 39964 11578 39976
rect 11974 39964 11980 39976
rect 11572 39936 11980 39964
rect 11572 39924 11578 39936
rect 11974 39924 11980 39936
rect 12032 39924 12038 39976
rect 12434 39924 12440 39976
rect 12492 39964 12498 39976
rect 13188 39964 13216 40004
rect 13814 39992 13820 40004
rect 13872 39992 13878 40044
rect 13906 39992 13912 40044
rect 13964 40032 13970 40044
rect 13964 40004 15700 40032
rect 13964 39992 13970 40004
rect 12492 39936 13216 39964
rect 12492 39924 12498 39936
rect 13262 39924 13268 39976
rect 13320 39964 13326 39976
rect 13449 39967 13507 39973
rect 13449 39964 13461 39967
rect 13320 39936 13461 39964
rect 13320 39924 13326 39936
rect 13449 39933 13461 39936
rect 13495 39964 13507 39967
rect 13630 39964 13636 39976
rect 13495 39936 13636 39964
rect 13495 39933 13507 39936
rect 13449 39927 13507 39933
rect 13630 39924 13636 39936
rect 13688 39924 13694 39976
rect 15672 39973 15700 40004
rect 18892 39976 18920 40072
rect 19058 40060 19064 40072
rect 19116 40060 19122 40112
rect 19150 40060 19156 40112
rect 19208 40100 19214 40112
rect 19208 40072 19380 40100
rect 19208 40060 19214 40072
rect 15565 39967 15623 39973
rect 15565 39933 15577 39967
rect 15611 39933 15623 39967
rect 15565 39927 15623 39933
rect 15657 39967 15715 39973
rect 15657 39933 15669 39967
rect 15703 39933 15715 39967
rect 15657 39927 15715 39933
rect 3970 39856 3976 39908
rect 4028 39896 4034 39908
rect 14645 39899 14703 39905
rect 14645 39896 14657 39899
rect 4028 39868 8064 39896
rect 4028 39856 4034 39868
rect 4062 39788 4068 39840
rect 4120 39828 4126 39840
rect 7929 39831 7987 39837
rect 7929 39828 7941 39831
rect 4120 39800 7941 39828
rect 4120 39788 4126 39800
rect 7929 39797 7941 39800
rect 7975 39797 7987 39831
rect 8036 39828 8064 39868
rect 13372 39868 14657 39896
rect 11057 39831 11115 39837
rect 11057 39828 11069 39831
rect 8036 39800 11069 39828
rect 7929 39791 7987 39797
rect 11057 39797 11069 39800
rect 11103 39797 11115 39831
rect 11057 39791 11115 39797
rect 11698 39788 11704 39840
rect 11756 39828 11762 39840
rect 13372 39828 13400 39868
rect 14645 39865 14657 39868
rect 14691 39896 14703 39899
rect 15580 39896 15608 39927
rect 18322 39924 18328 39976
rect 18380 39924 18386 39976
rect 18874 39924 18880 39976
rect 18932 39924 18938 39976
rect 19352 39964 19380 40072
rect 19978 40060 19984 40112
rect 20036 40060 20042 40112
rect 21266 40100 21272 40112
rect 21206 40086 21272 40100
rect 21192 40072 21272 40086
rect 19702 39992 19708 40044
rect 19760 39992 19766 40044
rect 21192 39964 21220 40072
rect 21266 40060 21272 40072
rect 21324 40060 21330 40112
rect 21450 40060 21456 40112
rect 21508 40100 21514 40112
rect 22020 40109 22048 40140
rect 22005 40103 22063 40109
rect 21508 40072 21956 40100
rect 21508 40060 21514 40072
rect 21928 40032 21956 40072
rect 22005 40069 22017 40103
rect 22051 40069 22063 40103
rect 24762 40100 24768 40112
rect 22005 40063 22063 40069
rect 22112 40072 24768 40100
rect 22112 40032 22140 40072
rect 24762 40060 24768 40072
rect 24820 40100 24826 40112
rect 24820 40072 24900 40100
rect 24820 40060 24826 40072
rect 21928 40004 22140 40032
rect 23474 39992 23480 40044
rect 23532 40032 23538 40044
rect 24670 40032 24676 40044
rect 23532 40004 24676 40032
rect 23532 39992 23538 40004
rect 24670 39992 24676 40004
rect 24728 39992 24734 40044
rect 19352 39936 21220 39964
rect 21542 39924 21548 39976
rect 21600 39964 21606 39976
rect 22741 39967 22799 39973
rect 22741 39964 22753 39967
rect 21600 39936 22753 39964
rect 21600 39924 21606 39936
rect 22741 39933 22753 39936
rect 22787 39933 22799 39967
rect 22741 39927 22799 39933
rect 23842 39924 23848 39976
rect 23900 39964 23906 39976
rect 24872 39973 24900 40072
rect 24765 39967 24823 39973
rect 24765 39964 24777 39967
rect 23900 39936 24777 39964
rect 23900 39924 23906 39936
rect 24765 39933 24777 39936
rect 24811 39933 24823 39967
rect 24765 39927 24823 39933
rect 24857 39967 24915 39973
rect 24857 39933 24869 39967
rect 24903 39933 24915 39967
rect 24857 39927 24915 39933
rect 14691 39868 16068 39896
rect 14691 39865 14703 39868
rect 14645 39859 14703 39865
rect 11756 39800 13400 39828
rect 11756 39788 11762 39800
rect 15102 39788 15108 39840
rect 15160 39788 15166 39840
rect 16040 39828 16068 39868
rect 21008 39868 31754 39896
rect 21008 39828 21036 39868
rect 16040 39800 21036 39828
rect 21450 39788 21456 39840
rect 21508 39788 21514 39840
rect 21910 39788 21916 39840
rect 21968 39828 21974 39840
rect 23566 39828 23572 39840
rect 21968 39800 23572 39828
rect 21968 39788 21974 39800
rect 23566 39788 23572 39800
rect 23624 39788 23630 39840
rect 23842 39788 23848 39840
rect 23900 39788 23906 39840
rect 24302 39788 24308 39840
rect 24360 39788 24366 39840
rect 31726 39828 31754 39868
rect 38654 39828 38660 39840
rect 31726 39800 38660 39828
rect 38654 39788 38660 39800
rect 38712 39788 38718 39840
rect 1104 39738 49864 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 32950 39738
rect 33002 39686 33014 39738
rect 33066 39686 33078 39738
rect 33130 39686 33142 39738
rect 33194 39686 33206 39738
rect 33258 39686 42950 39738
rect 43002 39686 43014 39738
rect 43066 39686 43078 39738
rect 43130 39686 43142 39738
rect 43194 39686 43206 39738
rect 43258 39686 49864 39738
rect 1104 39664 49864 39686
rect 7558 39584 7564 39636
rect 7616 39624 7622 39636
rect 8202 39624 8208 39636
rect 7616 39596 8208 39624
rect 7616 39584 7622 39596
rect 8202 39584 8208 39596
rect 8260 39584 8266 39636
rect 8573 39627 8631 39633
rect 8573 39593 8585 39627
rect 8619 39624 8631 39627
rect 9030 39624 9036 39636
rect 8619 39596 9036 39624
rect 8619 39593 8631 39596
rect 8573 39587 8631 39593
rect 9030 39584 9036 39596
rect 9088 39584 9094 39636
rect 10597 39627 10655 39633
rect 10597 39593 10609 39627
rect 10643 39624 10655 39627
rect 10778 39624 10784 39636
rect 10643 39596 10784 39624
rect 10643 39593 10655 39596
rect 10597 39587 10655 39593
rect 10778 39584 10784 39596
rect 10836 39584 10842 39636
rect 11793 39627 11851 39633
rect 11793 39593 11805 39627
rect 11839 39624 11851 39627
rect 12250 39624 12256 39636
rect 11839 39596 12256 39624
rect 11839 39593 11851 39596
rect 11793 39587 11851 39593
rect 12250 39584 12256 39596
rect 12308 39584 12314 39636
rect 13173 39627 13231 39633
rect 13173 39593 13185 39627
rect 13219 39624 13231 39627
rect 13354 39624 13360 39636
rect 13219 39596 13360 39624
rect 13219 39593 13231 39596
rect 13173 39587 13231 39593
rect 13354 39584 13360 39596
rect 13412 39584 13418 39636
rect 14642 39584 14648 39636
rect 14700 39624 14706 39636
rect 14829 39627 14887 39633
rect 14829 39624 14841 39627
rect 14700 39596 14841 39624
rect 14700 39584 14706 39596
rect 14829 39593 14841 39596
rect 14875 39593 14887 39627
rect 14829 39587 14887 39593
rect 16482 39584 16488 39636
rect 16540 39584 16546 39636
rect 16942 39584 16948 39636
rect 17000 39584 17006 39636
rect 18141 39627 18199 39633
rect 18141 39593 18153 39627
rect 18187 39624 18199 39627
rect 18414 39624 18420 39636
rect 18187 39596 18420 39624
rect 18187 39593 18199 39596
rect 18141 39587 18199 39593
rect 18414 39584 18420 39596
rect 18472 39584 18478 39636
rect 37826 39624 37832 39636
rect 18524 39596 37832 39624
rect 1854 39516 1860 39568
rect 1912 39556 1918 39568
rect 14734 39556 14740 39568
rect 1912 39528 2544 39556
rect 1912 39516 1918 39528
rect 2516 39500 2544 39528
rect 12452 39528 14740 39556
rect 1302 39448 1308 39500
rect 1360 39488 1366 39500
rect 2041 39491 2099 39497
rect 2041 39488 2053 39491
rect 1360 39460 2053 39488
rect 1360 39448 1366 39460
rect 2041 39457 2053 39460
rect 2087 39457 2099 39491
rect 2041 39451 2099 39457
rect 2498 39448 2504 39500
rect 2556 39488 2562 39500
rect 5537 39491 5595 39497
rect 5537 39488 5549 39491
rect 2556 39460 5549 39488
rect 2556 39448 2562 39460
rect 5537 39457 5549 39460
rect 5583 39457 5595 39491
rect 5537 39451 5595 39457
rect 5721 39491 5779 39497
rect 5721 39457 5733 39491
rect 5767 39488 5779 39491
rect 6546 39488 6552 39500
rect 5767 39460 6552 39488
rect 5767 39457 5779 39460
rect 5721 39451 5779 39457
rect 6546 39448 6552 39460
rect 6604 39448 6610 39500
rect 6825 39491 6883 39497
rect 6825 39457 6837 39491
rect 6871 39488 6883 39491
rect 8478 39488 8484 39500
rect 6871 39460 8484 39488
rect 6871 39457 6883 39460
rect 6825 39451 6883 39457
rect 8478 39448 8484 39460
rect 8536 39448 8542 39500
rect 8662 39448 8668 39500
rect 8720 39488 8726 39500
rect 9677 39491 9735 39497
rect 9677 39488 9689 39491
rect 8720 39460 9689 39488
rect 8720 39448 8726 39460
rect 9677 39457 9689 39460
rect 9723 39457 9735 39491
rect 11057 39491 11115 39497
rect 11057 39488 11069 39491
rect 9677 39451 9735 39457
rect 9784 39460 11069 39488
rect 1765 39423 1823 39429
rect 1765 39389 1777 39423
rect 1811 39420 1823 39423
rect 4614 39420 4620 39432
rect 1811 39392 4620 39420
rect 1811 39389 1823 39392
rect 1765 39383 1823 39389
rect 4614 39380 4620 39392
rect 4672 39380 4678 39432
rect 5442 39380 5448 39432
rect 5500 39380 5506 39432
rect 8202 39380 8208 39432
rect 8260 39380 8266 39432
rect 9030 39380 9036 39432
rect 9088 39420 9094 39432
rect 9784 39420 9812 39460
rect 11057 39457 11069 39460
rect 11103 39457 11115 39491
rect 11057 39451 11115 39457
rect 11238 39448 11244 39500
rect 11296 39448 11302 39500
rect 12452 39497 12480 39528
rect 14734 39516 14740 39528
rect 14792 39516 14798 39568
rect 17770 39516 17776 39568
rect 17828 39556 17834 39568
rect 18524 39556 18552 39596
rect 37826 39584 37832 39596
rect 37884 39584 37890 39636
rect 19794 39556 19800 39568
rect 17828 39528 18552 39556
rect 18616 39528 19800 39556
rect 17828 39516 17834 39528
rect 12437 39491 12495 39497
rect 12437 39457 12449 39491
rect 12483 39457 12495 39491
rect 12437 39451 12495 39457
rect 13817 39491 13875 39497
rect 13817 39457 13829 39491
rect 13863 39457 13875 39491
rect 13817 39451 13875 39457
rect 9088 39392 9812 39420
rect 9088 39380 9094 39392
rect 11882 39380 11888 39432
rect 11940 39420 11946 39432
rect 12161 39423 12219 39429
rect 12161 39420 12173 39423
rect 11940 39392 12173 39420
rect 11940 39380 11946 39392
rect 12161 39389 12173 39392
rect 12207 39389 12219 39423
rect 12161 39383 12219 39389
rect 12250 39380 12256 39432
rect 12308 39380 12314 39432
rect 12894 39380 12900 39432
rect 12952 39420 12958 39432
rect 13832 39420 13860 39451
rect 13998 39448 14004 39500
rect 14056 39488 14062 39500
rect 15194 39488 15200 39500
rect 14056 39460 15200 39488
rect 14056 39448 14062 39460
rect 15194 39448 15200 39460
rect 15252 39448 15258 39500
rect 15473 39491 15531 39497
rect 15473 39457 15485 39491
rect 15519 39488 15531 39491
rect 15562 39488 15568 39500
rect 15519 39460 15568 39488
rect 15519 39457 15531 39460
rect 15473 39451 15531 39457
rect 15562 39448 15568 39460
rect 15620 39448 15626 39500
rect 17586 39448 17592 39500
rect 17644 39448 17650 39500
rect 18616 39420 18644 39528
rect 19794 39516 19800 39528
rect 19852 39516 19858 39568
rect 21726 39516 21732 39568
rect 21784 39556 21790 39568
rect 23201 39559 23259 39565
rect 23201 39556 23213 39559
rect 21784 39528 23213 39556
rect 21784 39516 21790 39528
rect 23201 39525 23213 39528
rect 23247 39525 23259 39559
rect 23201 39519 23259 39525
rect 18785 39491 18843 39497
rect 18785 39457 18797 39491
rect 18831 39457 18843 39491
rect 18785 39451 18843 39457
rect 12952 39392 13860 39420
rect 13924 39392 18644 39420
rect 18800 39420 18828 39451
rect 19702 39448 19708 39500
rect 19760 39488 19766 39500
rect 20349 39491 20407 39497
rect 20349 39488 20361 39491
rect 19760 39460 20361 39488
rect 19760 39448 19766 39460
rect 20349 39457 20361 39460
rect 20395 39457 20407 39491
rect 20349 39451 20407 39457
rect 20625 39491 20683 39497
rect 20625 39457 20637 39491
rect 20671 39488 20683 39491
rect 21910 39488 21916 39500
rect 20671 39460 21916 39488
rect 20671 39457 20683 39460
rect 20625 39451 20683 39457
rect 21910 39448 21916 39460
rect 21968 39448 21974 39500
rect 22094 39448 22100 39500
rect 22152 39448 22158 39500
rect 22738 39448 22744 39500
rect 22796 39448 22802 39500
rect 23290 39448 23296 39500
rect 23348 39488 23354 39500
rect 23753 39491 23811 39497
rect 23753 39488 23765 39491
rect 23348 39460 23765 39488
rect 23348 39448 23354 39460
rect 23753 39457 23765 39460
rect 23799 39457 23811 39491
rect 23753 39451 23811 39457
rect 19978 39420 19984 39432
rect 18800 39392 19984 39420
rect 12952 39380 12958 39392
rect 7101 39355 7159 39361
rect 7101 39321 7113 39355
rect 7147 39321 7159 39355
rect 7101 39315 7159 39321
rect 5077 39287 5135 39293
rect 5077 39253 5089 39287
rect 5123 39284 5135 39287
rect 5810 39284 5816 39296
rect 5123 39256 5816 39284
rect 5123 39253 5135 39256
rect 5077 39247 5135 39253
rect 5810 39244 5816 39256
rect 5868 39244 5874 39296
rect 7116 39284 7144 39315
rect 8662 39312 8668 39364
rect 8720 39352 8726 39364
rect 9585 39355 9643 39361
rect 9585 39352 9597 39355
rect 8720 39324 9597 39352
rect 8720 39312 8726 39324
rect 9585 39321 9597 39324
rect 9631 39321 9643 39355
rect 9585 39315 9643 39321
rect 10965 39355 11023 39361
rect 10965 39321 10977 39355
rect 11011 39352 11023 39355
rect 12066 39352 12072 39364
rect 11011 39324 12072 39352
rect 11011 39321 11023 39324
rect 10965 39315 11023 39321
rect 12066 39312 12072 39324
rect 12124 39312 12130 39364
rect 13633 39355 13691 39361
rect 13633 39321 13645 39355
rect 13679 39352 13691 39355
rect 13924 39352 13952 39392
rect 19978 39380 19984 39392
rect 20036 39380 20042 39432
rect 22557 39423 22615 39429
rect 22557 39389 22569 39423
rect 22603 39420 22615 39423
rect 24302 39420 24308 39432
rect 22603 39392 24308 39420
rect 22603 39389 22615 39392
rect 22557 39383 22615 39389
rect 24302 39380 24308 39392
rect 24360 39380 24366 39432
rect 13679 39324 13952 39352
rect 17405 39355 17463 39361
rect 13679 39321 13691 39324
rect 13633 39315 13691 39321
rect 17405 39321 17417 39355
rect 17451 39352 17463 39355
rect 20346 39352 20352 39364
rect 17451 39324 20352 39352
rect 17451 39321 17463 39324
rect 17405 39315 17463 39321
rect 20346 39312 20352 39324
rect 20404 39312 20410 39364
rect 21266 39312 21272 39364
rect 21324 39312 21330 39364
rect 22649 39355 22707 39361
rect 22649 39321 22661 39355
rect 22695 39352 22707 39355
rect 24578 39352 24584 39364
rect 22695 39324 24584 39352
rect 22695 39321 22707 39324
rect 22649 39315 22707 39321
rect 24578 39312 24584 39324
rect 24636 39312 24642 39364
rect 8570 39284 8576 39296
rect 7116 39256 8576 39284
rect 8570 39244 8576 39256
rect 8628 39244 8634 39296
rect 9122 39244 9128 39296
rect 9180 39244 9186 39296
rect 9490 39244 9496 39296
rect 9548 39244 9554 39296
rect 12618 39244 12624 39296
rect 12676 39284 12682 39296
rect 13541 39287 13599 39293
rect 13541 39284 13553 39287
rect 12676 39256 13553 39284
rect 12676 39244 12682 39256
rect 13541 39253 13553 39256
rect 13587 39253 13599 39287
rect 13541 39247 13599 39253
rect 14182 39244 14188 39296
rect 14240 39284 14246 39296
rect 14458 39284 14464 39296
rect 14240 39256 14464 39284
rect 14240 39244 14246 39256
rect 14458 39244 14464 39256
rect 14516 39244 14522 39296
rect 15194 39244 15200 39296
rect 15252 39244 15258 39296
rect 15286 39244 15292 39296
rect 15344 39244 15350 39296
rect 17218 39244 17224 39296
rect 17276 39284 17282 39296
rect 17313 39287 17371 39293
rect 17313 39284 17325 39287
rect 17276 39256 17325 39284
rect 17276 39244 17282 39256
rect 17313 39253 17325 39256
rect 17359 39253 17371 39287
rect 17313 39247 17371 39253
rect 18414 39244 18420 39296
rect 18472 39284 18478 39296
rect 18509 39287 18567 39293
rect 18509 39284 18521 39287
rect 18472 39256 18521 39284
rect 18472 39244 18478 39256
rect 18509 39253 18521 39256
rect 18555 39253 18567 39287
rect 18509 39247 18567 39253
rect 18601 39287 18659 39293
rect 18601 39253 18613 39287
rect 18647 39284 18659 39287
rect 21634 39284 21640 39296
rect 18647 39256 21640 39284
rect 18647 39253 18659 39256
rect 18601 39247 18659 39253
rect 21634 39244 21640 39256
rect 21692 39244 21698 39296
rect 22186 39244 22192 39296
rect 22244 39244 22250 39296
rect 23566 39244 23572 39296
rect 23624 39244 23630 39296
rect 23661 39287 23719 39293
rect 23661 39253 23673 39287
rect 23707 39284 23719 39287
rect 23750 39284 23756 39296
rect 23707 39256 23756 39284
rect 23707 39253 23719 39256
rect 23661 39247 23719 39253
rect 23750 39244 23756 39256
rect 23808 39244 23814 39296
rect 1104 39194 49864 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 27950 39194
rect 28002 39142 28014 39194
rect 28066 39142 28078 39194
rect 28130 39142 28142 39194
rect 28194 39142 28206 39194
rect 28258 39142 37950 39194
rect 38002 39142 38014 39194
rect 38066 39142 38078 39194
rect 38130 39142 38142 39194
rect 38194 39142 38206 39194
rect 38258 39142 47950 39194
rect 48002 39142 48014 39194
rect 48066 39142 48078 39194
rect 48130 39142 48142 39194
rect 48194 39142 48206 39194
rect 48258 39142 49864 39194
rect 1104 39120 49864 39142
rect 5629 39083 5687 39089
rect 5629 39049 5641 39083
rect 5675 39080 5687 39083
rect 5718 39080 5724 39092
rect 5675 39052 5724 39080
rect 5675 39049 5687 39052
rect 5629 39043 5687 39049
rect 5718 39040 5724 39052
rect 5776 39040 5782 39092
rect 10134 39080 10140 39092
rect 9140 39052 10140 39080
rect 6641 39015 6699 39021
rect 6641 38981 6653 39015
rect 6687 39012 6699 39015
rect 7282 39012 7288 39024
rect 6687 38984 7288 39012
rect 6687 38981 6699 38984
rect 6641 38975 6699 38981
rect 7282 38972 7288 38984
rect 7340 38972 7346 39024
rect 8202 38972 8208 39024
rect 8260 39012 8266 39024
rect 9140 39012 9168 39052
rect 10134 39040 10140 39052
rect 10192 39040 10198 39092
rect 12161 39083 12219 39089
rect 12161 39049 12173 39083
rect 12207 39080 12219 39083
rect 12526 39080 12532 39092
rect 12207 39052 12532 39080
rect 12207 39049 12219 39052
rect 12161 39043 12219 39049
rect 12526 39040 12532 39052
rect 12584 39040 12590 39092
rect 12989 39083 13047 39089
rect 12989 39049 13001 39083
rect 13035 39080 13047 39083
rect 13170 39080 13176 39092
rect 13035 39052 13176 39080
rect 13035 39049 13047 39052
rect 12989 39043 13047 39049
rect 13170 39040 13176 39052
rect 13228 39040 13234 39092
rect 13357 39083 13415 39089
rect 13357 39080 13369 39083
rect 13280 39052 13369 39080
rect 10965 39015 11023 39021
rect 8260 38984 9246 39012
rect 8260 38972 8266 38984
rect 10965 38981 10977 39015
rect 11011 39012 11023 39015
rect 11698 39012 11704 39024
rect 11011 38984 11704 39012
rect 11011 38981 11023 38984
rect 10965 38975 11023 38981
rect 11698 38972 11704 38984
rect 11756 38972 11762 39024
rect 12710 38972 12716 39024
rect 12768 39012 12774 39024
rect 13280 39012 13308 39052
rect 13357 39049 13369 39052
rect 13403 39049 13415 39083
rect 13357 39043 13415 39049
rect 14182 39040 14188 39092
rect 14240 39040 14246 39092
rect 15010 39040 15016 39092
rect 15068 39080 15074 39092
rect 16853 39083 16911 39089
rect 16853 39080 16865 39083
rect 15068 39052 16865 39080
rect 15068 39040 15074 39052
rect 16853 39049 16865 39052
rect 16899 39049 16911 39083
rect 16853 39043 16911 39049
rect 16942 39040 16948 39092
rect 17000 39080 17006 39092
rect 17313 39083 17371 39089
rect 17313 39080 17325 39083
rect 17000 39052 17325 39080
rect 17000 39040 17006 39052
rect 17313 39049 17325 39052
rect 17359 39080 17371 39083
rect 17770 39080 17776 39092
rect 17359 39052 17776 39080
rect 17359 39049 17371 39052
rect 17313 39043 17371 39049
rect 17770 39040 17776 39052
rect 17828 39080 17834 39092
rect 18049 39083 18107 39089
rect 18049 39080 18061 39083
rect 17828 39052 18061 39080
rect 17828 39040 17834 39052
rect 18049 39049 18061 39052
rect 18095 39049 18107 39083
rect 18049 39043 18107 39049
rect 19978 39040 19984 39092
rect 20036 39080 20042 39092
rect 20625 39083 20683 39089
rect 20625 39080 20637 39083
rect 20036 39052 20637 39080
rect 20036 39040 20042 39052
rect 20625 39049 20637 39052
rect 20671 39049 20683 39083
rect 22833 39083 22891 39089
rect 22833 39080 22845 39083
rect 20625 39043 20683 39049
rect 22066 39052 22845 39080
rect 12768 38984 13308 39012
rect 14553 39015 14611 39021
rect 12768 38972 12774 38984
rect 14553 38981 14565 39015
rect 14599 39012 14611 39015
rect 21266 39012 21272 39024
rect 14599 38984 16252 39012
rect 20378 38984 21272 39012
rect 14599 38981 14611 38984
rect 14553 38975 14611 38981
rect 5258 38904 5264 38956
rect 5316 38944 5322 38956
rect 7653 38947 7711 38953
rect 7653 38944 7665 38947
rect 5316 38916 7665 38944
rect 5316 38904 5322 38916
rect 7653 38913 7665 38916
rect 7699 38913 7711 38947
rect 7653 38907 7711 38913
rect 8478 38904 8484 38956
rect 8536 38904 8542 38956
rect 12526 38904 12532 38956
rect 12584 38904 12590 38956
rect 12621 38947 12679 38953
rect 12621 38913 12633 38947
rect 12667 38944 12679 38947
rect 13078 38944 13084 38956
rect 12667 38916 13084 38944
rect 12667 38913 12679 38916
rect 12621 38907 12679 38913
rect 13078 38904 13084 38916
rect 13136 38904 13142 38956
rect 13998 38904 14004 38956
rect 14056 38904 14062 38956
rect 14645 38947 14703 38953
rect 14645 38913 14657 38947
rect 14691 38944 14703 38947
rect 15470 38944 15476 38956
rect 14691 38916 15476 38944
rect 14691 38913 14703 38916
rect 14645 38907 14703 38913
rect 15470 38904 15476 38916
rect 15528 38904 15534 38956
rect 15565 38947 15623 38953
rect 15565 38913 15577 38947
rect 15611 38944 15623 38947
rect 16022 38944 16028 38956
rect 15611 38916 16028 38944
rect 15611 38913 15623 38916
rect 15565 38907 15623 38913
rect 16022 38904 16028 38916
rect 16080 38904 16086 38956
rect 16224 38953 16252 38984
rect 21266 38972 21272 38984
rect 21324 38972 21330 39024
rect 16209 38947 16267 38953
rect 16209 38913 16221 38947
rect 16255 38913 16267 38947
rect 16209 38907 16267 38913
rect 16850 38904 16856 38956
rect 16908 38944 16914 38956
rect 17221 38947 17279 38953
rect 17221 38944 17233 38947
rect 16908 38916 17233 38944
rect 16908 38904 16914 38916
rect 17221 38913 17233 38916
rect 17267 38913 17279 38947
rect 17221 38907 17279 38913
rect 18230 38904 18236 38956
rect 18288 38944 18294 38956
rect 18417 38947 18475 38953
rect 18417 38944 18429 38947
rect 18288 38916 18429 38944
rect 18288 38904 18294 38916
rect 18417 38913 18429 38916
rect 18463 38913 18475 38947
rect 18417 38907 18475 38913
rect 4982 38836 4988 38888
rect 5040 38876 5046 38888
rect 5721 38879 5779 38885
rect 5721 38876 5733 38879
rect 5040 38848 5733 38876
rect 5040 38836 5046 38848
rect 5721 38845 5733 38848
rect 5767 38845 5779 38879
rect 5721 38839 5779 38845
rect 5905 38879 5963 38885
rect 5905 38845 5917 38879
rect 5951 38876 5963 38879
rect 6454 38876 6460 38888
rect 5951 38848 6460 38876
rect 5951 38845 5963 38848
rect 5905 38839 5963 38845
rect 6454 38836 6460 38848
rect 6512 38836 6518 38888
rect 7190 38836 7196 38888
rect 7248 38876 7254 38888
rect 7745 38879 7803 38885
rect 7745 38876 7757 38879
rect 7248 38848 7757 38876
rect 7248 38836 7254 38848
rect 7745 38845 7757 38848
rect 7791 38845 7803 38879
rect 7745 38839 7803 38845
rect 7929 38879 7987 38885
rect 7929 38845 7941 38879
rect 7975 38876 7987 38879
rect 8757 38879 8815 38885
rect 8757 38876 8769 38879
rect 7975 38848 8769 38876
rect 7975 38845 7987 38848
rect 7929 38839 7987 38845
rect 8496 38820 8524 38848
rect 8757 38845 8769 38848
rect 8803 38845 8815 38879
rect 8757 38839 8815 38845
rect 9122 38836 9128 38888
rect 9180 38876 9186 38888
rect 11882 38876 11888 38888
rect 9180 38848 11888 38876
rect 9180 38836 9186 38848
rect 11882 38836 11888 38848
rect 11940 38836 11946 38888
rect 12805 38879 12863 38885
rect 12805 38845 12817 38879
rect 12851 38876 12863 38879
rect 12986 38876 12992 38888
rect 12851 38848 12992 38876
rect 12851 38845 12863 38848
rect 12805 38839 12863 38845
rect 12986 38836 12992 38848
rect 13044 38836 13050 38888
rect 13446 38836 13452 38888
rect 13504 38836 13510 38888
rect 13630 38836 13636 38888
rect 13688 38836 13694 38888
rect 14734 38836 14740 38888
rect 14792 38836 14798 38888
rect 17405 38879 17463 38885
rect 17405 38845 17417 38879
rect 17451 38845 17463 38879
rect 17405 38839 17463 38845
rect 5626 38768 5632 38820
rect 5684 38808 5690 38820
rect 7285 38811 7343 38817
rect 7285 38808 7297 38811
rect 5684 38780 7297 38808
rect 5684 38768 5690 38780
rect 7285 38777 7297 38780
rect 7331 38777 7343 38811
rect 7285 38771 7343 38777
rect 8478 38768 8484 38820
rect 8536 38768 8542 38820
rect 11146 38768 11152 38820
rect 11204 38768 11210 38820
rect 14274 38808 14280 38820
rect 13556 38780 14280 38808
rect 5261 38743 5319 38749
rect 5261 38709 5273 38743
rect 5307 38740 5319 38743
rect 5350 38740 5356 38752
rect 5307 38712 5356 38740
rect 5307 38709 5319 38712
rect 5261 38703 5319 38709
rect 5350 38700 5356 38712
rect 5408 38700 5414 38752
rect 6086 38700 6092 38752
rect 6144 38740 6150 38752
rect 6733 38743 6791 38749
rect 6733 38740 6745 38743
rect 6144 38712 6745 38740
rect 6144 38700 6150 38712
rect 6733 38709 6745 38712
rect 6779 38709 6791 38743
rect 6733 38703 6791 38709
rect 8938 38700 8944 38752
rect 8996 38740 9002 38752
rect 9766 38740 9772 38752
rect 8996 38712 9772 38740
rect 8996 38700 9002 38712
rect 9766 38700 9772 38712
rect 9824 38740 9830 38752
rect 10229 38743 10287 38749
rect 10229 38740 10241 38743
rect 9824 38712 10241 38740
rect 9824 38700 9830 38712
rect 10229 38709 10241 38712
rect 10275 38709 10287 38743
rect 10229 38703 10287 38709
rect 11238 38700 11244 38752
rect 11296 38740 11302 38752
rect 13556 38740 13584 38780
rect 14274 38768 14280 38780
rect 14332 38768 14338 38820
rect 11296 38712 13584 38740
rect 11296 38700 11302 38712
rect 13998 38700 14004 38752
rect 14056 38740 14062 38752
rect 15381 38743 15439 38749
rect 15381 38740 15393 38743
rect 14056 38712 15393 38740
rect 14056 38700 14062 38712
rect 15381 38709 15393 38712
rect 15427 38709 15439 38743
rect 15381 38703 15439 38709
rect 15654 38700 15660 38752
rect 15712 38740 15718 38752
rect 17420 38740 17448 38839
rect 18690 38836 18696 38888
rect 18748 38876 18754 38888
rect 18877 38879 18935 38885
rect 18877 38876 18889 38879
rect 18748 38848 18889 38876
rect 18748 38836 18754 38848
rect 18877 38845 18889 38848
rect 18923 38845 18935 38879
rect 18877 38839 18935 38845
rect 19153 38879 19211 38885
rect 19153 38845 19165 38879
rect 19199 38876 19211 38879
rect 19242 38876 19248 38888
rect 19199 38848 19248 38876
rect 19199 38845 19211 38848
rect 19153 38839 19211 38845
rect 19242 38836 19248 38848
rect 19300 38836 19306 38888
rect 19886 38836 19892 38888
rect 19944 38876 19950 38888
rect 20162 38876 20168 38888
rect 19944 38848 20168 38876
rect 19944 38836 19950 38848
rect 20162 38836 20168 38848
rect 20220 38876 20226 38888
rect 22066 38876 22094 39052
rect 22833 39049 22845 39052
rect 22879 39080 22891 39083
rect 23842 39080 23848 39092
rect 22879 39052 23848 39080
rect 22879 39049 22891 39052
rect 22833 39043 22891 39049
rect 23842 39040 23848 39052
rect 23900 39080 23906 39092
rect 23900 39052 31754 39080
rect 23900 39040 23906 39052
rect 23474 38904 23480 38956
rect 23532 38944 23538 38956
rect 23753 38947 23811 38953
rect 23753 38944 23765 38947
rect 23532 38916 23765 38944
rect 23532 38904 23538 38916
rect 23753 38913 23765 38916
rect 23799 38913 23811 38947
rect 23753 38907 23811 38913
rect 20220 38848 22094 38876
rect 20220 38836 20226 38848
rect 22554 38836 22560 38888
rect 22612 38876 22618 38888
rect 23290 38876 23296 38888
rect 22612 38848 23296 38876
rect 22612 38836 22618 38848
rect 23290 38836 23296 38848
rect 23348 38876 23354 38888
rect 23937 38879 23995 38885
rect 23937 38876 23949 38879
rect 23348 38848 23949 38876
rect 23348 38836 23354 38848
rect 23937 38845 23949 38848
rect 23983 38845 23995 38879
rect 31726 38876 31754 39052
rect 48866 38876 48872 38888
rect 31726 38848 48872 38876
rect 23937 38839 23995 38845
rect 48866 38836 48872 38848
rect 48924 38836 48930 38888
rect 21634 38768 21640 38820
rect 21692 38808 21698 38820
rect 23385 38811 23443 38817
rect 23385 38808 23397 38811
rect 21692 38780 23397 38808
rect 21692 38768 21698 38780
rect 23385 38777 23397 38780
rect 23431 38777 23443 38811
rect 23385 38771 23443 38777
rect 15712 38712 17448 38740
rect 15712 38700 15718 38712
rect 18414 38700 18420 38752
rect 18472 38740 18478 38752
rect 19150 38740 19156 38752
rect 18472 38712 19156 38740
rect 18472 38700 18478 38712
rect 19150 38700 19156 38712
rect 19208 38700 19214 38752
rect 19242 38700 19248 38752
rect 19300 38740 19306 38752
rect 22094 38740 22100 38752
rect 19300 38712 22100 38740
rect 19300 38700 19306 38712
rect 22094 38700 22100 38712
rect 22152 38700 22158 38752
rect 1104 38650 49864 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 32950 38650
rect 33002 38598 33014 38650
rect 33066 38598 33078 38650
rect 33130 38598 33142 38650
rect 33194 38598 33206 38650
rect 33258 38598 42950 38650
rect 43002 38598 43014 38650
rect 43066 38598 43078 38650
rect 43130 38598 43142 38650
rect 43194 38598 43206 38650
rect 43258 38598 49864 38650
rect 1104 38576 49864 38598
rect 4614 38496 4620 38548
rect 4672 38496 4678 38548
rect 5258 38496 5264 38548
rect 5316 38496 5322 38548
rect 5718 38496 5724 38548
rect 5776 38536 5782 38548
rect 6914 38536 6920 38548
rect 5776 38508 6920 38536
rect 5776 38496 5782 38508
rect 6914 38496 6920 38508
rect 6972 38496 6978 38548
rect 9217 38539 9275 38545
rect 9217 38505 9229 38539
rect 9263 38536 9275 38539
rect 9490 38536 9496 38548
rect 9263 38508 9496 38536
rect 9263 38505 9275 38508
rect 9217 38499 9275 38505
rect 9490 38496 9496 38508
rect 9548 38496 9554 38548
rect 11974 38496 11980 38548
rect 12032 38536 12038 38548
rect 13725 38539 13783 38545
rect 13725 38536 13737 38539
rect 12032 38508 13737 38536
rect 12032 38496 12038 38508
rect 13725 38505 13737 38508
rect 13771 38505 13783 38539
rect 15102 38536 15108 38548
rect 13725 38499 13783 38505
rect 13832 38508 15108 38536
rect 8294 38428 8300 38480
rect 8352 38468 8358 38480
rect 8573 38471 8631 38477
rect 8573 38468 8585 38471
rect 8352 38440 8585 38468
rect 8352 38428 8358 38440
rect 8573 38437 8585 38440
rect 8619 38468 8631 38471
rect 9306 38468 9312 38480
rect 8619 38440 9312 38468
rect 8619 38437 8631 38440
rect 8573 38431 8631 38437
rect 9306 38428 9312 38440
rect 9364 38428 9370 38480
rect 1302 38360 1308 38412
rect 1360 38400 1366 38412
rect 2041 38403 2099 38409
rect 2041 38400 2053 38403
rect 1360 38372 2053 38400
rect 1360 38360 1366 38372
rect 2041 38369 2053 38372
rect 2087 38369 2099 38403
rect 5534 38400 5540 38412
rect 2041 38363 2099 38369
rect 2746 38372 5540 38400
rect 1765 38335 1823 38341
rect 1765 38301 1777 38335
rect 1811 38332 1823 38335
rect 2746 38332 2774 38372
rect 5534 38360 5540 38372
rect 5592 38360 5598 38412
rect 5813 38403 5871 38409
rect 5813 38369 5825 38403
rect 5859 38400 5871 38403
rect 6730 38400 6736 38412
rect 5859 38372 6736 38400
rect 5859 38369 5871 38372
rect 5813 38363 5871 38369
rect 6730 38360 6736 38372
rect 6788 38360 6794 38412
rect 7101 38403 7159 38409
rect 7101 38369 7113 38403
rect 7147 38400 7159 38403
rect 8846 38400 8852 38412
rect 7147 38372 8852 38400
rect 7147 38369 7159 38372
rect 7101 38363 7159 38369
rect 8846 38360 8852 38372
rect 8904 38400 8910 38412
rect 9398 38400 9404 38412
rect 8904 38372 9404 38400
rect 8904 38360 8910 38372
rect 9398 38360 9404 38372
rect 9456 38360 9462 38412
rect 9490 38360 9496 38412
rect 9548 38400 9554 38412
rect 9766 38400 9772 38412
rect 9548 38372 9772 38400
rect 9548 38360 9554 38372
rect 9766 38360 9772 38372
rect 9824 38360 9830 38412
rect 10962 38360 10968 38412
rect 11020 38360 11026 38412
rect 13832 38400 13860 38508
rect 15102 38496 15108 38508
rect 15160 38496 15166 38548
rect 19058 38496 19064 38548
rect 19116 38536 19122 38548
rect 22281 38539 22339 38545
rect 22281 38536 22293 38539
rect 19116 38508 22293 38536
rect 19116 38496 19122 38508
rect 22281 38505 22293 38508
rect 22327 38536 22339 38539
rect 22738 38536 22744 38548
rect 22327 38508 22744 38536
rect 22327 38505 22339 38508
rect 22281 38499 22339 38505
rect 22738 38496 22744 38508
rect 22796 38496 22802 38548
rect 17862 38428 17868 38480
rect 17920 38468 17926 38480
rect 18233 38471 18291 38477
rect 18233 38468 18245 38471
rect 17920 38440 18245 38468
rect 17920 38428 17926 38440
rect 18233 38437 18245 38440
rect 18279 38437 18291 38471
rect 18233 38431 18291 38437
rect 11072 38372 13860 38400
rect 1811 38304 2774 38332
rect 4801 38335 4859 38341
rect 1811 38301 1823 38304
rect 1765 38295 1823 38301
rect 4801 38301 4813 38335
rect 4847 38301 4859 38335
rect 4801 38295 4859 38301
rect 5629 38335 5687 38341
rect 5629 38301 5641 38335
rect 5675 38332 5687 38335
rect 5902 38332 5908 38344
rect 5675 38304 5908 38332
rect 5675 38301 5687 38304
rect 5629 38295 5687 38301
rect 4816 38264 4844 38295
rect 5902 38292 5908 38304
rect 5960 38292 5966 38344
rect 6822 38292 6828 38344
rect 6880 38292 6886 38344
rect 8202 38292 8208 38344
rect 8260 38332 8266 38344
rect 8386 38332 8392 38344
rect 8260 38304 8392 38332
rect 8260 38292 8266 38304
rect 8386 38292 8392 38304
rect 8444 38292 8450 38344
rect 9585 38335 9643 38341
rect 9585 38301 9597 38335
rect 9631 38332 9643 38335
rect 11072 38332 11100 38372
rect 14550 38360 14556 38412
rect 14608 38400 14614 38412
rect 16482 38400 16488 38412
rect 14608 38372 16488 38400
rect 14608 38360 14614 38372
rect 16482 38360 16488 38372
rect 16540 38400 16546 38412
rect 18322 38400 18328 38412
rect 16540 38372 18328 38400
rect 16540 38360 16546 38372
rect 18322 38360 18328 38372
rect 18380 38360 18386 38412
rect 20809 38403 20867 38409
rect 20809 38369 20821 38403
rect 20855 38400 20867 38403
rect 21450 38400 21456 38412
rect 20855 38372 21456 38400
rect 20855 38369 20867 38372
rect 20809 38363 20867 38369
rect 21450 38360 21456 38372
rect 21508 38360 21514 38412
rect 23753 38403 23811 38409
rect 23753 38369 23765 38403
rect 23799 38400 23811 38403
rect 23934 38400 23940 38412
rect 23799 38372 23940 38400
rect 23799 38369 23811 38372
rect 23753 38363 23811 38369
rect 23934 38360 23940 38372
rect 23992 38360 23998 38412
rect 9631 38304 11100 38332
rect 9631 38301 9643 38304
rect 9585 38295 9643 38301
rect 11974 38292 11980 38344
rect 12032 38292 12038 38344
rect 14274 38292 14280 38344
rect 14332 38292 14338 38344
rect 20530 38292 20536 38344
rect 20588 38292 20594 38344
rect 22830 38292 22836 38344
rect 22888 38332 22894 38344
rect 23477 38335 23535 38341
rect 23477 38332 23489 38335
rect 22888 38304 23489 38332
rect 22888 38292 22894 38304
rect 23477 38301 23489 38304
rect 23523 38301 23535 38335
rect 23477 38295 23535 38301
rect 23566 38292 23572 38344
rect 23624 38332 23630 38344
rect 24394 38332 24400 38344
rect 23624 38304 24400 38332
rect 23624 38292 23630 38304
rect 24394 38292 24400 38304
rect 24452 38292 24458 38344
rect 7374 38264 7380 38276
rect 4816 38236 7380 38264
rect 7374 38224 7380 38236
rect 7432 38224 7438 38276
rect 9858 38264 9864 38276
rect 8404 38236 9864 38264
rect 5442 38156 5448 38208
rect 5500 38196 5506 38208
rect 5721 38199 5779 38205
rect 5721 38196 5733 38199
rect 5500 38168 5733 38196
rect 5500 38156 5506 38168
rect 5721 38165 5733 38168
rect 5767 38165 5779 38199
rect 5721 38159 5779 38165
rect 6638 38156 6644 38208
rect 6696 38196 6702 38208
rect 8404 38196 8432 38236
rect 9858 38224 9864 38236
rect 9916 38224 9922 38276
rect 9950 38224 9956 38276
rect 10008 38264 10014 38276
rect 10781 38267 10839 38273
rect 10781 38264 10793 38267
rect 10008 38236 10793 38264
rect 10008 38224 10014 38236
rect 10781 38233 10793 38236
rect 10827 38233 10839 38267
rect 10781 38227 10839 38233
rect 12253 38267 12311 38273
rect 12253 38233 12265 38267
rect 12299 38264 12311 38267
rect 12299 38236 12664 38264
rect 12299 38233 12311 38236
rect 12253 38227 12311 38233
rect 6696 38168 8432 38196
rect 6696 38156 6702 38168
rect 8846 38156 8852 38208
rect 8904 38196 8910 38208
rect 9677 38199 9735 38205
rect 9677 38196 9689 38199
rect 8904 38168 9689 38196
rect 8904 38156 8910 38168
rect 9677 38165 9689 38168
rect 9723 38165 9735 38199
rect 9677 38159 9735 38165
rect 9766 38156 9772 38208
rect 9824 38196 9830 38208
rect 10413 38199 10471 38205
rect 10413 38196 10425 38199
rect 9824 38168 10425 38196
rect 9824 38156 9830 38168
rect 10413 38165 10425 38168
rect 10459 38165 10471 38199
rect 10413 38159 10471 38165
rect 10870 38156 10876 38208
rect 10928 38156 10934 38208
rect 11054 38156 11060 38208
rect 11112 38196 11118 38208
rect 12526 38196 12532 38208
rect 11112 38168 12532 38196
rect 11112 38156 11118 38168
rect 12526 38156 12532 38168
rect 12584 38156 12590 38208
rect 12636 38196 12664 38236
rect 12710 38224 12716 38276
rect 12768 38224 12774 38276
rect 14553 38267 14611 38273
rect 14553 38233 14565 38267
rect 14599 38264 14611 38267
rect 14826 38264 14832 38276
rect 14599 38236 14832 38264
rect 14599 38233 14611 38236
rect 14553 38227 14611 38233
rect 14826 38224 14832 38236
rect 14884 38224 14890 38276
rect 14936 38236 15042 38264
rect 13078 38196 13084 38208
rect 12636 38168 13084 38196
rect 13078 38156 13084 38168
rect 13136 38156 13142 38208
rect 14458 38156 14464 38208
rect 14516 38196 14522 38208
rect 14936 38196 14964 38236
rect 16666 38224 16672 38276
rect 16724 38264 16730 38276
rect 16761 38267 16819 38273
rect 16761 38264 16773 38267
rect 16724 38236 16773 38264
rect 16724 38224 16730 38236
rect 16761 38233 16773 38236
rect 16807 38233 16819 38267
rect 16761 38227 16819 38233
rect 17218 38224 17224 38276
rect 17276 38224 17282 38276
rect 18064 38236 18368 38264
rect 14516 38168 14964 38196
rect 14516 38156 14522 38168
rect 15562 38156 15568 38208
rect 15620 38196 15626 38208
rect 16025 38199 16083 38205
rect 16025 38196 16037 38199
rect 15620 38168 16037 38196
rect 15620 38156 15626 38168
rect 16025 38165 16037 38168
rect 16071 38165 16083 38199
rect 16025 38159 16083 38165
rect 16114 38156 16120 38208
rect 16172 38196 16178 38208
rect 18064 38196 18092 38236
rect 16172 38168 18092 38196
rect 18340 38196 18368 38236
rect 21266 38224 21272 38276
rect 21324 38224 21330 38276
rect 22278 38196 22284 38208
rect 18340 38168 22284 38196
rect 16172 38156 16178 38168
rect 22278 38156 22284 38168
rect 22336 38156 22342 38208
rect 22370 38156 22376 38208
rect 22428 38196 22434 38208
rect 23109 38199 23167 38205
rect 23109 38196 23121 38199
rect 22428 38168 23121 38196
rect 22428 38156 22434 38168
rect 23109 38165 23121 38168
rect 23155 38165 23167 38199
rect 23109 38159 23167 38165
rect 1104 38106 49864 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 27950 38106
rect 28002 38054 28014 38106
rect 28066 38054 28078 38106
rect 28130 38054 28142 38106
rect 28194 38054 28206 38106
rect 28258 38054 37950 38106
rect 38002 38054 38014 38106
rect 38066 38054 38078 38106
rect 38130 38054 38142 38106
rect 38194 38054 38206 38106
rect 38258 38054 47950 38106
rect 48002 38054 48014 38106
rect 48066 38054 48078 38106
rect 48130 38054 48142 38106
rect 48194 38054 48206 38106
rect 48258 38054 49864 38106
rect 1104 38032 49864 38054
rect 4338 37952 4344 38004
rect 4396 37952 4402 38004
rect 5629 37995 5687 38001
rect 5629 37961 5641 37995
rect 5675 37992 5687 37995
rect 5902 37992 5908 38004
rect 5675 37964 5908 37992
rect 5675 37961 5687 37964
rect 5629 37955 5687 37961
rect 5902 37952 5908 37964
rect 5960 37952 5966 38004
rect 7282 37992 7288 38004
rect 6564 37964 7288 37992
rect 5718 37924 5724 37936
rect 2746 37896 5724 37924
rect 1765 37859 1823 37865
rect 1765 37825 1777 37859
rect 1811 37856 1823 37859
rect 2746 37856 2774 37896
rect 5718 37884 5724 37896
rect 5776 37884 5782 37936
rect 1811 37828 2774 37856
rect 4249 37859 4307 37865
rect 1811 37825 1823 37828
rect 1765 37819 1823 37825
rect 4249 37825 4261 37859
rect 4295 37856 4307 37859
rect 6564 37856 6592 37964
rect 7282 37952 7288 37964
rect 7340 37992 7346 38004
rect 7466 37992 7472 38004
rect 7340 37964 7472 37992
rect 7340 37952 7346 37964
rect 7466 37952 7472 37964
rect 7524 37952 7530 38004
rect 8570 37952 8576 38004
rect 8628 37952 8634 38004
rect 8938 37952 8944 38004
rect 8996 37992 9002 38004
rect 9582 37992 9588 38004
rect 8996 37964 9588 37992
rect 8996 37952 9002 37964
rect 9582 37952 9588 37964
rect 9640 37952 9646 38004
rect 9677 37995 9735 38001
rect 9677 37961 9689 37995
rect 9723 37992 9735 37995
rect 9858 37992 9864 38004
rect 9723 37964 9864 37992
rect 9723 37961 9735 37964
rect 9677 37955 9735 37961
rect 9858 37952 9864 37964
rect 9916 37952 9922 38004
rect 10413 37995 10471 38001
rect 10413 37961 10425 37995
rect 10459 37992 10471 37995
rect 11606 37992 11612 38004
rect 10459 37964 11612 37992
rect 10459 37961 10471 37964
rect 10413 37955 10471 37961
rect 11606 37952 11612 37964
rect 11664 37952 11670 38004
rect 12158 37952 12164 38004
rect 12216 37992 12222 38004
rect 12529 37995 12587 38001
rect 12529 37992 12541 37995
rect 12216 37964 12541 37992
rect 12216 37952 12222 37964
rect 12529 37961 12541 37964
rect 12575 37961 12587 37995
rect 12529 37955 12587 37961
rect 12710 37952 12716 38004
rect 12768 37992 12774 38004
rect 14458 37992 14464 38004
rect 12768 37964 14464 37992
rect 12768 37952 12774 37964
rect 14458 37952 14464 37964
rect 14516 37952 14522 38004
rect 17862 37992 17868 38004
rect 14844 37964 17868 37992
rect 10962 37924 10968 37936
rect 9968 37896 10968 37924
rect 4295 37828 6592 37856
rect 4295 37825 4307 37828
rect 4249 37819 4307 37825
rect 8202 37816 8208 37868
rect 8260 37856 8266 37868
rect 8386 37856 8392 37868
rect 8260 37828 8392 37856
rect 8260 37816 8266 37828
rect 8386 37816 8392 37828
rect 8444 37816 8450 37868
rect 1302 37748 1308 37800
rect 1360 37788 1366 37800
rect 2041 37791 2099 37797
rect 2041 37788 2053 37791
rect 1360 37760 2053 37788
rect 1360 37748 1366 37760
rect 2041 37757 2053 37760
rect 2087 37757 2099 37791
rect 2041 37751 2099 37757
rect 4522 37748 4528 37800
rect 4580 37788 4586 37800
rect 4890 37788 4896 37800
rect 4580 37760 4896 37788
rect 4580 37748 4586 37760
rect 4890 37748 4896 37760
rect 4948 37788 4954 37800
rect 5442 37788 5448 37800
rect 4948 37760 5448 37788
rect 4948 37748 4954 37760
rect 5442 37748 5448 37760
rect 5500 37788 5506 37800
rect 5721 37791 5779 37797
rect 5721 37788 5733 37791
rect 5500 37760 5733 37788
rect 5500 37748 5506 37760
rect 5721 37757 5733 37760
rect 5767 37757 5779 37791
rect 5721 37751 5779 37757
rect 5902 37748 5908 37800
rect 5960 37748 5966 37800
rect 6822 37748 6828 37800
rect 6880 37748 6886 37800
rect 7101 37791 7159 37797
rect 7101 37757 7113 37791
rect 7147 37788 7159 37791
rect 8294 37788 8300 37800
rect 7147 37760 8300 37788
rect 7147 37757 7159 37760
rect 7101 37751 7159 37757
rect 8294 37748 8300 37760
rect 8352 37748 8358 37800
rect 9858 37748 9864 37800
rect 9916 37788 9922 37800
rect 9968 37788 9996 37896
rect 10962 37884 10968 37896
rect 11020 37884 11026 37936
rect 13814 37884 13820 37936
rect 13872 37884 13878 37936
rect 14844 37933 14872 37964
rect 17862 37952 17868 37964
rect 17920 37952 17926 38004
rect 22278 37952 22284 38004
rect 22336 37992 22342 38004
rect 23109 37995 23167 38001
rect 23109 37992 23121 37995
rect 22336 37964 23121 37992
rect 22336 37952 22342 37964
rect 23109 37961 23121 37964
rect 23155 37961 23167 37995
rect 23109 37955 23167 37961
rect 23201 37995 23259 38001
rect 23201 37961 23213 37995
rect 23247 37992 23259 37995
rect 23382 37992 23388 38004
rect 23247 37964 23388 37992
rect 23247 37961 23259 37964
rect 23201 37955 23259 37961
rect 23382 37952 23388 37964
rect 23440 37952 23446 38004
rect 14829 37927 14887 37933
rect 14829 37893 14841 37927
rect 14875 37893 14887 37927
rect 14829 37887 14887 37893
rect 15378 37884 15384 37936
rect 15436 37884 15442 37936
rect 17218 37884 17224 37936
rect 17276 37924 17282 37936
rect 17276 37896 17710 37924
rect 17276 37884 17282 37896
rect 18598 37884 18604 37936
rect 18656 37924 18662 37936
rect 18782 37924 18788 37936
rect 18656 37896 18788 37924
rect 18656 37884 18662 37896
rect 18782 37884 18788 37896
rect 18840 37884 18846 37936
rect 20073 37927 20131 37933
rect 20073 37893 20085 37927
rect 20119 37924 20131 37927
rect 20714 37924 20720 37936
rect 20119 37896 20720 37924
rect 20119 37893 20131 37896
rect 20073 37887 20131 37893
rect 20714 37884 20720 37896
rect 20772 37924 20778 37936
rect 22002 37924 22008 37936
rect 20772 37896 22008 37924
rect 20772 37884 20778 37896
rect 22002 37884 22008 37896
rect 22060 37884 22066 37936
rect 10781 37859 10839 37865
rect 10781 37825 10793 37859
rect 10827 37856 10839 37859
rect 11885 37859 11943 37865
rect 11885 37856 11897 37859
rect 10827 37828 11897 37856
rect 10827 37825 10839 37828
rect 10781 37819 10839 37825
rect 11885 37825 11897 37828
rect 11931 37825 11943 37859
rect 11885 37819 11943 37825
rect 12618 37816 12624 37868
rect 12676 37856 12682 37868
rect 12897 37859 12955 37865
rect 12897 37856 12909 37859
rect 12676 37828 12909 37856
rect 12676 37816 12682 37828
rect 12897 37825 12909 37828
rect 12943 37825 12955 37859
rect 12897 37819 12955 37825
rect 14550 37816 14556 37868
rect 14608 37816 14614 37868
rect 16482 37816 16488 37868
rect 16540 37856 16546 37868
rect 16945 37859 17003 37865
rect 16945 37856 16957 37859
rect 16540 37828 16957 37856
rect 16540 37816 16546 37828
rect 16945 37825 16957 37828
rect 16991 37825 17003 37859
rect 16945 37819 17003 37825
rect 9916 37760 9996 37788
rect 9916 37748 9922 37760
rect 10134 37748 10140 37800
rect 10192 37788 10198 37800
rect 10873 37791 10931 37797
rect 10873 37788 10885 37791
rect 10192 37760 10885 37788
rect 10192 37748 10198 37760
rect 10873 37757 10885 37760
rect 10919 37757 10931 37791
rect 10873 37751 10931 37757
rect 10965 37791 11023 37797
rect 10965 37757 10977 37791
rect 11011 37757 11023 37791
rect 10965 37751 11023 37757
rect 8110 37680 8116 37732
rect 8168 37720 8174 37732
rect 9490 37720 9496 37732
rect 8168 37692 9496 37720
rect 8168 37680 8174 37692
rect 9490 37680 9496 37692
rect 9548 37680 9554 37732
rect 10980 37720 11008 37751
rect 12986 37748 12992 37800
rect 13044 37748 13050 37800
rect 13078 37748 13084 37800
rect 13136 37788 13142 37800
rect 13722 37788 13728 37800
rect 13136 37760 13728 37788
rect 13136 37748 13142 37760
rect 13722 37748 13728 37760
rect 13780 37748 13786 37800
rect 14090 37788 14096 37800
rect 13924 37760 14096 37788
rect 13924 37720 13952 37760
rect 14090 37748 14096 37760
rect 14148 37748 14154 37800
rect 15194 37748 15200 37800
rect 15252 37788 15258 37800
rect 16114 37788 16120 37800
rect 15252 37760 16120 37788
rect 15252 37748 15258 37760
rect 16114 37748 16120 37760
rect 16172 37748 16178 37800
rect 17221 37791 17279 37797
rect 17221 37757 17233 37791
rect 17267 37788 17279 37791
rect 17586 37788 17592 37800
rect 17267 37760 17592 37788
rect 17267 37757 17279 37760
rect 17221 37751 17279 37757
rect 17586 37748 17592 37760
rect 17644 37788 17650 37800
rect 18782 37788 18788 37800
rect 17644 37760 18788 37788
rect 17644 37748 17650 37760
rect 18782 37748 18788 37760
rect 18840 37748 18846 37800
rect 20162 37748 20168 37800
rect 20220 37788 20226 37800
rect 20530 37788 20536 37800
rect 20220 37760 20536 37788
rect 20220 37748 20226 37760
rect 20530 37748 20536 37760
rect 20588 37788 20594 37800
rect 20809 37791 20867 37797
rect 20809 37788 20821 37791
rect 20588 37760 20821 37788
rect 20588 37748 20594 37760
rect 20809 37757 20821 37760
rect 20855 37757 20867 37791
rect 20809 37751 20867 37757
rect 23290 37748 23296 37800
rect 23348 37748 23354 37800
rect 10980 37692 13952 37720
rect 14001 37723 14059 37729
rect 14001 37689 14013 37723
rect 14047 37720 14059 37723
rect 14550 37720 14556 37732
rect 14047 37692 14556 37720
rect 14047 37689 14059 37692
rect 14001 37683 14059 37689
rect 14550 37680 14556 37692
rect 14608 37680 14614 37732
rect 5261 37655 5319 37661
rect 5261 37621 5273 37655
rect 5307 37652 5319 37655
rect 8386 37652 8392 37664
rect 5307 37624 8392 37652
rect 5307 37621 5319 37624
rect 5261 37615 5319 37621
rect 8386 37612 8392 37624
rect 8444 37612 8450 37664
rect 9214 37612 9220 37664
rect 9272 37612 9278 37664
rect 14826 37612 14832 37664
rect 14884 37652 14890 37664
rect 16301 37655 16359 37661
rect 16301 37652 16313 37655
rect 14884 37624 16313 37652
rect 14884 37612 14890 37624
rect 16301 37621 16313 37624
rect 16347 37621 16359 37655
rect 16301 37615 16359 37621
rect 16666 37612 16672 37664
rect 16724 37652 16730 37664
rect 18693 37655 18751 37661
rect 18693 37652 18705 37655
rect 16724 37624 18705 37652
rect 16724 37612 16730 37624
rect 18693 37621 18705 37624
rect 18739 37621 18751 37655
rect 18693 37615 18751 37621
rect 21358 37612 21364 37664
rect 21416 37652 21422 37664
rect 22741 37655 22799 37661
rect 22741 37652 22753 37655
rect 21416 37624 22753 37652
rect 21416 37612 21422 37624
rect 22741 37621 22753 37624
rect 22787 37621 22799 37655
rect 22741 37615 22799 37621
rect 1104 37562 49864 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 32950 37562
rect 33002 37510 33014 37562
rect 33066 37510 33078 37562
rect 33130 37510 33142 37562
rect 33194 37510 33206 37562
rect 33258 37510 42950 37562
rect 43002 37510 43014 37562
rect 43066 37510 43078 37562
rect 43130 37510 43142 37562
rect 43194 37510 43206 37562
rect 43258 37510 49864 37562
rect 1104 37488 49864 37510
rect 5902 37408 5908 37460
rect 5960 37448 5966 37460
rect 5960 37420 8248 37448
rect 5960 37408 5966 37420
rect 8018 37380 8024 37392
rect 5828 37352 8024 37380
rect 5626 37272 5632 37324
rect 5684 37272 5690 37324
rect 5828 37321 5856 37352
rect 8018 37340 8024 37352
rect 8076 37340 8082 37392
rect 5813 37315 5871 37321
rect 5813 37281 5825 37315
rect 5859 37281 5871 37315
rect 5813 37275 5871 37281
rect 6638 37272 6644 37324
rect 6696 37312 6702 37324
rect 6825 37315 6883 37321
rect 6825 37312 6837 37315
rect 6696 37284 6837 37312
rect 6696 37272 6702 37284
rect 6825 37281 6837 37284
rect 6871 37281 6883 37315
rect 6825 37275 6883 37281
rect 7009 37315 7067 37321
rect 7009 37281 7021 37315
rect 7055 37312 7067 37315
rect 7374 37312 7380 37324
rect 7055 37284 7380 37312
rect 7055 37281 7067 37284
rect 7009 37275 7067 37281
rect 7374 37272 7380 37284
rect 7432 37272 7438 37324
rect 8220 37321 8248 37420
rect 8294 37408 8300 37460
rect 8352 37448 8358 37460
rect 11054 37448 11060 37460
rect 8352 37420 11060 37448
rect 8352 37408 8358 37420
rect 11054 37408 11060 37420
rect 11112 37408 11118 37460
rect 13722 37408 13728 37460
rect 13780 37408 13786 37460
rect 18782 37408 18788 37460
rect 18840 37408 18846 37460
rect 22278 37408 22284 37460
rect 22336 37448 22342 37460
rect 23934 37448 23940 37460
rect 22336 37420 23940 37448
rect 22336 37408 22342 37420
rect 23934 37408 23940 37420
rect 23992 37408 23998 37460
rect 9858 37380 9864 37392
rect 9600 37352 9864 37380
rect 8205 37315 8263 37321
rect 7576 37284 8064 37312
rect 7576 37244 7604 37284
rect 6288 37216 7604 37244
rect 6288 37176 6316 37216
rect 7650 37204 7656 37256
rect 7708 37244 7714 37256
rect 7929 37247 7987 37253
rect 7929 37244 7941 37247
rect 7708 37216 7941 37244
rect 7708 37204 7714 37216
rect 7929 37213 7941 37216
rect 7975 37213 7987 37247
rect 8036 37244 8064 37284
rect 8205 37281 8217 37315
rect 8251 37312 8263 37315
rect 9600 37312 9628 37352
rect 9858 37340 9864 37352
rect 9916 37380 9922 37392
rect 10226 37380 10232 37392
rect 9916 37352 10232 37380
rect 9916 37340 9922 37352
rect 10226 37340 10232 37352
rect 10284 37340 10290 37392
rect 8251 37284 9628 37312
rect 8251 37281 8263 37284
rect 8205 37275 8263 37281
rect 9674 37272 9680 37324
rect 9732 37312 9738 37324
rect 11241 37315 11299 37321
rect 11241 37312 11253 37315
rect 9732 37284 11253 37312
rect 9732 37272 9738 37284
rect 11241 37281 11253 37284
rect 11287 37281 11299 37315
rect 11241 37275 11299 37281
rect 12253 37315 12311 37321
rect 12253 37281 12265 37315
rect 12299 37312 12311 37315
rect 13538 37312 13544 37324
rect 12299 37284 13544 37312
rect 12299 37281 12311 37284
rect 12253 37275 12311 37281
rect 13538 37272 13544 37284
rect 13596 37272 13602 37324
rect 14274 37272 14280 37324
rect 14332 37312 14338 37324
rect 14645 37315 14703 37321
rect 14645 37312 14657 37315
rect 14332 37284 14657 37312
rect 14332 37272 14338 37284
rect 14645 37281 14657 37284
rect 14691 37281 14703 37315
rect 14645 37275 14703 37281
rect 14921 37315 14979 37321
rect 14921 37281 14933 37315
rect 14967 37312 14979 37315
rect 15562 37312 15568 37324
rect 14967 37284 15568 37312
rect 14967 37281 14979 37284
rect 14921 37275 14979 37281
rect 15562 37272 15568 37284
rect 15620 37272 15626 37324
rect 16114 37272 16120 37324
rect 16172 37312 16178 37324
rect 17313 37315 17371 37321
rect 17313 37312 17325 37315
rect 16172 37284 17325 37312
rect 16172 37272 16178 37284
rect 17313 37281 17325 37284
rect 17359 37312 17371 37315
rect 18874 37312 18880 37324
rect 17359 37284 18880 37312
rect 17359 37281 17371 37284
rect 17313 37275 17371 37281
rect 18874 37272 18880 37284
rect 18932 37272 18938 37324
rect 21450 37272 21456 37324
rect 21508 37312 21514 37324
rect 23290 37312 23296 37324
rect 21508 37284 23296 37312
rect 21508 37272 21514 37284
rect 23290 37272 23296 37284
rect 23348 37272 23354 37324
rect 8662 37244 8668 37256
rect 8036 37216 8668 37244
rect 7929 37207 7987 37213
rect 8662 37204 8668 37216
rect 8720 37204 8726 37256
rect 9030 37204 9036 37256
rect 9088 37244 9094 37256
rect 10321 37247 10379 37253
rect 10321 37244 10333 37247
rect 9088 37216 10333 37244
rect 9088 37204 9094 37216
rect 10321 37213 10333 37216
rect 10367 37213 10379 37247
rect 10321 37207 10379 37213
rect 11054 37204 11060 37256
rect 11112 37204 11118 37256
rect 11974 37204 11980 37256
rect 12032 37204 12038 37256
rect 17037 37247 17095 37253
rect 17037 37213 17049 37247
rect 17083 37213 17095 37247
rect 17037 37207 17095 37213
rect 7190 37176 7196 37188
rect 5184 37148 6316 37176
rect 6380 37148 7196 37176
rect 5184 37117 5212 37148
rect 5169 37111 5227 37117
rect 5169 37077 5181 37111
rect 5215 37077 5227 37111
rect 5169 37071 5227 37077
rect 5534 37068 5540 37120
rect 5592 37068 5598 37120
rect 6380 37117 6408 37148
rect 7190 37136 7196 37148
rect 7248 37136 7254 37188
rect 7466 37136 7472 37188
rect 7524 37176 7530 37188
rect 7524 37148 7788 37176
rect 7524 37136 7530 37148
rect 6365 37111 6423 37117
rect 6365 37077 6377 37111
rect 6411 37077 6423 37111
rect 6365 37071 6423 37077
rect 6730 37068 6736 37120
rect 6788 37068 6794 37120
rect 7558 37068 7564 37120
rect 7616 37068 7622 37120
rect 7760 37108 7788 37148
rect 7834 37136 7840 37188
rect 7892 37176 7898 37188
rect 9490 37176 9496 37188
rect 7892 37148 9496 37176
rect 7892 37136 7898 37148
rect 9490 37136 9496 37148
rect 9548 37176 9554 37188
rect 9585 37179 9643 37185
rect 9585 37176 9597 37179
rect 9548 37148 9597 37176
rect 9548 37136 9554 37148
rect 9585 37145 9597 37148
rect 9631 37145 9643 37179
rect 9585 37139 9643 37145
rect 12710 37136 12716 37188
rect 12768 37136 12774 37188
rect 14458 37136 14464 37188
rect 14516 37176 14522 37188
rect 15378 37176 15384 37188
rect 14516 37148 15384 37176
rect 14516 37136 14522 37148
rect 15378 37136 15384 37148
rect 15436 37136 15442 37188
rect 8021 37111 8079 37117
rect 8021 37108 8033 37111
rect 7760 37080 8033 37108
rect 8021 37077 8033 37080
rect 8067 37077 8079 37111
rect 8021 37071 8079 37077
rect 8202 37068 8208 37120
rect 8260 37108 8266 37120
rect 10410 37108 10416 37120
rect 8260 37080 10416 37108
rect 8260 37068 8266 37080
rect 10410 37068 10416 37080
rect 10468 37068 10474 37120
rect 15930 37068 15936 37120
rect 15988 37108 15994 37120
rect 16393 37111 16451 37117
rect 16393 37108 16405 37111
rect 15988 37080 16405 37108
rect 15988 37068 15994 37080
rect 16393 37077 16405 37080
rect 16439 37077 16451 37111
rect 17052 37108 17080 37207
rect 18690 37204 18696 37256
rect 18748 37244 18754 37256
rect 20162 37244 20168 37256
rect 18748 37216 20168 37244
rect 18748 37204 18754 37216
rect 20162 37204 20168 37216
rect 20220 37244 20226 37256
rect 20533 37247 20591 37253
rect 20533 37244 20545 37247
rect 20220 37216 20545 37244
rect 20220 37204 20226 37216
rect 20533 37213 20545 37216
rect 20579 37213 20591 37247
rect 20533 37207 20591 37213
rect 22830 37204 22836 37256
rect 22888 37244 22894 37256
rect 23109 37247 23167 37253
rect 23109 37244 23121 37247
rect 22888 37216 23121 37244
rect 22888 37204 22894 37216
rect 23109 37213 23121 37216
rect 23155 37213 23167 37247
rect 23109 37207 23167 37213
rect 23201 37247 23259 37253
rect 23201 37213 23213 37247
rect 23247 37244 23259 37247
rect 23566 37244 23572 37256
rect 23247 37216 23572 37244
rect 23247 37213 23259 37216
rect 23201 37207 23259 37213
rect 23566 37204 23572 37216
rect 23624 37204 23630 37256
rect 17218 37136 17224 37188
rect 17276 37176 17282 37188
rect 17402 37176 17408 37188
rect 17276 37148 17408 37176
rect 17276 37136 17282 37148
rect 17402 37136 17408 37148
rect 17460 37136 17466 37188
rect 17770 37136 17776 37188
rect 17828 37136 17834 37188
rect 18782 37136 18788 37188
rect 18840 37176 18846 37188
rect 18840 37148 20760 37176
rect 18840 37136 18846 37148
rect 20732 37120 20760 37148
rect 20806 37136 20812 37188
rect 20864 37136 20870 37188
rect 21266 37176 21272 37188
rect 20916 37148 21272 37176
rect 18690 37108 18696 37120
rect 17052 37080 18696 37108
rect 16393 37071 16451 37077
rect 18690 37068 18696 37080
rect 18748 37068 18754 37120
rect 20714 37068 20720 37120
rect 20772 37108 20778 37120
rect 20916 37108 20944 37148
rect 21266 37136 21272 37148
rect 21324 37136 21330 37188
rect 22204 37148 22784 37176
rect 20772 37080 20944 37108
rect 20772 37068 20778 37080
rect 21174 37068 21180 37120
rect 21232 37108 21238 37120
rect 22204 37108 22232 37148
rect 22756 37117 22784 37148
rect 21232 37080 22232 37108
rect 22741 37111 22799 37117
rect 21232 37068 21238 37080
rect 22741 37077 22753 37111
rect 22787 37077 22799 37111
rect 22741 37071 22799 37077
rect 1104 37018 49864 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 27950 37018
rect 28002 36966 28014 37018
rect 28066 36966 28078 37018
rect 28130 36966 28142 37018
rect 28194 36966 28206 37018
rect 28258 36966 37950 37018
rect 38002 36966 38014 37018
rect 38066 36966 38078 37018
rect 38130 36966 38142 37018
rect 38194 36966 38206 37018
rect 38258 36966 47950 37018
rect 48002 36966 48014 37018
rect 48066 36966 48078 37018
rect 48130 36966 48142 37018
rect 48194 36966 48206 37018
rect 48258 36966 49864 37018
rect 1104 36944 49864 36966
rect 5629 36907 5687 36913
rect 5629 36873 5641 36907
rect 5675 36904 5687 36907
rect 6178 36904 6184 36916
rect 5675 36876 6184 36904
rect 5675 36873 5687 36876
rect 5629 36867 5687 36873
rect 6178 36864 6184 36876
rect 6236 36864 6242 36916
rect 7009 36907 7067 36913
rect 7009 36873 7021 36907
rect 7055 36904 7067 36907
rect 7098 36904 7104 36916
rect 7055 36876 7104 36904
rect 7055 36873 7067 36876
rect 7009 36867 7067 36873
rect 7098 36864 7104 36876
rect 7156 36864 7162 36916
rect 7374 36864 7380 36916
rect 7432 36904 7438 36916
rect 7650 36904 7656 36916
rect 7432 36876 7656 36904
rect 7432 36864 7438 36876
rect 7650 36864 7656 36876
rect 7708 36864 7714 36916
rect 8386 36864 8392 36916
rect 8444 36864 8450 36916
rect 8481 36907 8539 36913
rect 8481 36873 8493 36907
rect 8527 36904 8539 36907
rect 9214 36904 9220 36916
rect 8527 36876 9220 36904
rect 8527 36873 8539 36876
rect 8481 36867 8539 36873
rect 9214 36864 9220 36876
rect 9272 36864 9278 36916
rect 9582 36864 9588 36916
rect 9640 36864 9646 36916
rect 10413 36907 10471 36913
rect 10413 36873 10425 36907
rect 10459 36904 10471 36907
rect 10594 36904 10600 36916
rect 10459 36876 10600 36904
rect 10459 36873 10471 36876
rect 10413 36867 10471 36873
rect 10594 36864 10600 36876
rect 10652 36864 10658 36916
rect 12618 36904 12624 36916
rect 11900 36876 12624 36904
rect 4617 36839 4675 36845
rect 4617 36805 4629 36839
rect 4663 36836 4675 36839
rect 5074 36836 5080 36848
rect 4663 36808 5080 36836
rect 4663 36805 4675 36808
rect 4617 36799 4675 36805
rect 5074 36796 5080 36808
rect 5132 36796 5138 36848
rect 6730 36796 6736 36848
rect 6788 36836 6794 36848
rect 8938 36836 8944 36848
rect 6788 36808 8944 36836
rect 6788 36796 6794 36808
rect 8938 36796 8944 36808
rect 8996 36796 9002 36848
rect 10873 36839 10931 36845
rect 10873 36836 10885 36839
rect 9048 36808 10885 36836
rect 1762 36728 1768 36780
rect 1820 36728 1826 36780
rect 6822 36728 6828 36780
rect 6880 36768 6886 36780
rect 6880 36740 7328 36768
rect 6880 36728 6886 36740
rect 1302 36660 1308 36712
rect 1360 36700 1366 36712
rect 2041 36703 2099 36709
rect 2041 36700 2053 36703
rect 1360 36672 2053 36700
rect 1360 36660 1366 36672
rect 2041 36669 2053 36672
rect 2087 36669 2099 36703
rect 2041 36663 2099 36669
rect 3510 36660 3516 36712
rect 3568 36700 3574 36712
rect 5721 36703 5779 36709
rect 5721 36700 5733 36703
rect 3568 36672 5733 36700
rect 3568 36660 3574 36672
rect 5721 36669 5733 36672
rect 5767 36669 5779 36703
rect 5721 36663 5779 36669
rect 5905 36703 5963 36709
rect 5905 36669 5917 36703
rect 5951 36700 5963 36703
rect 6546 36700 6552 36712
rect 5951 36672 6552 36700
rect 5951 36669 5963 36672
rect 5905 36663 5963 36669
rect 6546 36660 6552 36672
rect 6604 36660 6610 36712
rect 7098 36660 7104 36712
rect 7156 36660 7162 36712
rect 7300 36709 7328 36740
rect 7374 36728 7380 36780
rect 7432 36768 7438 36780
rect 9048 36768 9076 36808
rect 10873 36805 10885 36808
rect 10919 36805 10931 36839
rect 10873 36799 10931 36805
rect 7432 36740 9076 36768
rect 10781 36771 10839 36777
rect 7432 36728 7438 36740
rect 10781 36737 10793 36771
rect 10827 36768 10839 36771
rect 11790 36768 11796 36780
rect 10827 36740 11796 36768
rect 10827 36737 10839 36740
rect 10781 36731 10839 36737
rect 11790 36728 11796 36740
rect 11848 36728 11854 36780
rect 7285 36703 7343 36709
rect 7285 36669 7297 36703
rect 7331 36700 7343 36703
rect 7650 36700 7656 36712
rect 7331 36672 7656 36700
rect 7331 36669 7343 36672
rect 7285 36663 7343 36669
rect 7650 36660 7656 36672
rect 7708 36660 7714 36712
rect 8662 36660 8668 36712
rect 8720 36660 8726 36712
rect 9122 36660 9128 36712
rect 9180 36700 9186 36712
rect 9582 36700 9588 36712
rect 9180 36672 9588 36700
rect 9180 36660 9186 36672
rect 9582 36660 9588 36672
rect 9640 36700 9646 36712
rect 9677 36703 9735 36709
rect 9677 36700 9689 36703
rect 9640 36672 9689 36700
rect 9640 36660 9646 36672
rect 9677 36669 9689 36672
rect 9723 36669 9735 36703
rect 9677 36663 9735 36669
rect 9769 36703 9827 36709
rect 9769 36669 9781 36703
rect 9815 36700 9827 36703
rect 10594 36700 10600 36712
rect 9815 36672 10600 36700
rect 9815 36669 9827 36672
rect 9769 36663 9827 36669
rect 10594 36660 10600 36672
rect 10652 36660 10658 36712
rect 10965 36703 11023 36709
rect 10965 36669 10977 36703
rect 11011 36700 11023 36703
rect 11330 36700 11336 36712
rect 11011 36672 11336 36700
rect 11011 36669 11023 36672
rect 10965 36663 11023 36669
rect 11330 36660 11336 36672
rect 11388 36660 11394 36712
rect 3418 36592 3424 36644
rect 3476 36632 3482 36644
rect 7466 36632 7472 36644
rect 3476 36604 7472 36632
rect 3476 36592 3482 36604
rect 7466 36592 7472 36604
rect 7524 36592 7530 36644
rect 8021 36635 8079 36641
rect 8021 36601 8033 36635
rect 8067 36632 8079 36635
rect 9858 36632 9864 36644
rect 8067 36604 9864 36632
rect 8067 36601 8079 36604
rect 8021 36595 8079 36601
rect 9858 36592 9864 36604
rect 9916 36592 9922 36644
rect 9950 36592 9956 36644
rect 10008 36632 10014 36644
rect 11900 36632 11928 36876
rect 12618 36864 12624 36876
rect 12676 36864 12682 36916
rect 14737 36907 14795 36913
rect 14737 36873 14749 36907
rect 14783 36904 14795 36907
rect 15102 36904 15108 36916
rect 14783 36876 15108 36904
rect 14783 36873 14795 36876
rect 14737 36867 14795 36873
rect 15102 36864 15108 36876
rect 15160 36864 15166 36916
rect 15470 36864 15476 36916
rect 15528 36864 15534 36916
rect 15933 36907 15991 36913
rect 15933 36873 15945 36907
rect 15979 36904 15991 36907
rect 16390 36904 16396 36916
rect 15979 36876 16396 36904
rect 15979 36873 15991 36876
rect 15933 36867 15991 36873
rect 16390 36864 16396 36876
rect 16448 36864 16454 36916
rect 16574 36864 16580 36916
rect 16632 36904 16638 36916
rect 22005 36907 22063 36913
rect 22005 36904 22017 36907
rect 16632 36876 22017 36904
rect 16632 36864 16638 36876
rect 22005 36873 22017 36876
rect 22051 36873 22063 36907
rect 22005 36867 22063 36873
rect 22370 36864 22376 36916
rect 22428 36864 22434 36916
rect 22465 36907 22523 36913
rect 22465 36873 22477 36907
rect 22511 36904 22523 36907
rect 22646 36904 22652 36916
rect 22511 36876 22652 36904
rect 22511 36873 22523 36876
rect 22465 36867 22523 36873
rect 22646 36864 22652 36876
rect 22704 36864 22710 36916
rect 12066 36796 12072 36848
rect 12124 36836 12130 36848
rect 12989 36839 13047 36845
rect 12989 36836 13001 36839
rect 12124 36808 13001 36836
rect 12124 36796 12130 36808
rect 12989 36805 13001 36808
rect 13035 36836 13047 36839
rect 14274 36836 14280 36848
rect 13035 36808 14280 36836
rect 13035 36805 13047 36808
rect 12989 36799 13047 36805
rect 14274 36796 14280 36808
rect 14332 36796 14338 36848
rect 18046 36836 18052 36848
rect 14752 36808 18052 36836
rect 12161 36771 12219 36777
rect 12161 36737 12173 36771
rect 12207 36768 12219 36771
rect 12342 36768 12348 36780
rect 12207 36740 12348 36768
rect 12207 36737 12219 36740
rect 12161 36731 12219 36737
rect 12342 36728 12348 36740
rect 12400 36728 12406 36780
rect 13725 36771 13783 36777
rect 13725 36737 13737 36771
rect 13771 36737 13783 36771
rect 13725 36731 13783 36737
rect 13740 36700 13768 36731
rect 13814 36728 13820 36780
rect 13872 36768 13878 36780
rect 14645 36771 14703 36777
rect 14645 36768 14657 36771
rect 13872 36740 14657 36768
rect 13872 36728 13878 36740
rect 14645 36737 14657 36740
rect 14691 36737 14703 36771
rect 14645 36731 14703 36737
rect 14752 36700 14780 36808
rect 18046 36796 18052 36808
rect 18104 36796 18110 36848
rect 18141 36839 18199 36845
rect 18141 36805 18153 36839
rect 18187 36836 18199 36839
rect 18874 36836 18880 36848
rect 18187 36808 18880 36836
rect 18187 36805 18199 36808
rect 18141 36799 18199 36805
rect 18874 36796 18880 36808
rect 18932 36796 18938 36848
rect 19245 36839 19303 36845
rect 19245 36805 19257 36839
rect 19291 36836 19303 36839
rect 19334 36836 19340 36848
rect 19291 36808 19340 36836
rect 19291 36805 19303 36808
rect 19245 36799 19303 36805
rect 19334 36796 19340 36808
rect 19392 36796 19398 36848
rect 20714 36836 20720 36848
rect 20470 36808 20720 36836
rect 20714 36796 20720 36808
rect 20772 36796 20778 36848
rect 15194 36728 15200 36780
rect 15252 36768 15258 36780
rect 15841 36771 15899 36777
rect 15841 36768 15853 36771
rect 15252 36740 15853 36768
rect 15252 36728 15258 36740
rect 15841 36737 15853 36740
rect 15887 36737 15899 36771
rect 15841 36731 15899 36737
rect 16850 36728 16856 36780
rect 16908 36728 16914 36780
rect 16942 36728 16948 36780
rect 17000 36768 17006 36780
rect 17313 36771 17371 36777
rect 17313 36768 17325 36771
rect 17000 36740 17325 36768
rect 17000 36728 17006 36740
rect 17313 36737 17325 36740
rect 17359 36737 17371 36771
rect 17313 36731 17371 36737
rect 18233 36771 18291 36777
rect 18233 36737 18245 36771
rect 18279 36768 18291 36771
rect 18598 36768 18604 36780
rect 18279 36740 18604 36768
rect 18279 36737 18291 36740
rect 18233 36731 18291 36737
rect 18598 36728 18604 36740
rect 18656 36728 18662 36780
rect 18690 36728 18696 36780
rect 18748 36768 18754 36780
rect 18969 36771 19027 36777
rect 18969 36768 18981 36771
rect 18748 36740 18981 36768
rect 18748 36728 18754 36740
rect 18969 36737 18981 36740
rect 19015 36737 19027 36771
rect 23566 36768 23572 36780
rect 18969 36731 19027 36737
rect 22066 36740 23572 36768
rect 13740 36672 14780 36700
rect 14826 36660 14832 36712
rect 14884 36660 14890 36712
rect 16022 36660 16028 36712
rect 16080 36660 16086 36712
rect 17402 36660 17408 36712
rect 17460 36660 17466 36712
rect 17589 36703 17647 36709
rect 17589 36669 17601 36703
rect 17635 36669 17647 36703
rect 17589 36663 17647 36669
rect 18417 36703 18475 36709
rect 18417 36669 18429 36703
rect 18463 36700 18475 36703
rect 18782 36700 18788 36712
rect 18463 36672 18788 36700
rect 18463 36669 18475 36672
rect 18417 36663 18475 36669
rect 10008 36604 11928 36632
rect 14277 36635 14335 36641
rect 10008 36592 10014 36604
rect 14277 36601 14289 36635
rect 14323 36632 14335 36635
rect 15286 36632 15292 36644
rect 14323 36604 15292 36632
rect 14323 36601 14335 36604
rect 14277 36595 14335 36601
rect 15286 36592 15292 36604
rect 15344 36592 15350 36644
rect 17604 36632 17632 36663
rect 18782 36660 18788 36672
rect 18840 36660 18846 36712
rect 18874 36660 18880 36712
rect 18932 36700 18938 36712
rect 22066 36700 22094 36740
rect 23566 36728 23572 36740
rect 23624 36728 23630 36780
rect 18932 36672 22094 36700
rect 22557 36703 22615 36709
rect 18932 36660 18938 36672
rect 22557 36669 22569 36703
rect 22603 36669 22615 36703
rect 22557 36663 22615 36669
rect 17604 36604 19104 36632
rect 4706 36524 4712 36576
rect 4764 36524 4770 36576
rect 5261 36567 5319 36573
rect 5261 36533 5273 36567
rect 5307 36564 5319 36567
rect 5810 36564 5816 36576
rect 5307 36536 5816 36564
rect 5307 36533 5319 36536
rect 5261 36527 5319 36533
rect 5810 36524 5816 36536
rect 5868 36524 5874 36576
rect 6641 36567 6699 36573
rect 6641 36533 6653 36567
rect 6687 36564 6699 36567
rect 7926 36564 7932 36576
rect 6687 36536 7932 36564
rect 6687 36533 6699 36536
rect 6641 36527 6699 36533
rect 7926 36524 7932 36536
rect 7984 36524 7990 36576
rect 8294 36524 8300 36576
rect 8352 36564 8358 36576
rect 9217 36567 9275 36573
rect 9217 36564 9229 36567
rect 8352 36536 9229 36564
rect 8352 36524 8358 36536
rect 9217 36533 9229 36536
rect 9263 36533 9275 36567
rect 9217 36527 9275 36533
rect 11330 36524 11336 36576
rect 11388 36564 11394 36576
rect 13541 36567 13599 36573
rect 13541 36564 13553 36567
rect 11388 36536 13553 36564
rect 11388 36524 11394 36536
rect 13541 36533 13553 36536
rect 13587 36533 13599 36567
rect 13541 36527 13599 36533
rect 16945 36567 17003 36573
rect 16945 36533 16957 36567
rect 16991 36564 17003 36567
rect 17678 36564 17684 36576
rect 16991 36536 17684 36564
rect 16991 36533 17003 36536
rect 16945 36527 17003 36533
rect 17678 36524 17684 36536
rect 17736 36524 17742 36576
rect 17770 36524 17776 36576
rect 17828 36524 17834 36576
rect 18046 36524 18052 36576
rect 18104 36564 18110 36576
rect 18966 36564 18972 36576
rect 18104 36536 18972 36564
rect 18104 36524 18110 36536
rect 18966 36524 18972 36536
rect 19024 36524 19030 36576
rect 19076 36564 19104 36604
rect 21542 36592 21548 36644
rect 21600 36632 21606 36644
rect 22572 36632 22600 36663
rect 21600 36604 22600 36632
rect 21600 36592 21606 36604
rect 20717 36567 20775 36573
rect 20717 36564 20729 36567
rect 19076 36536 20729 36564
rect 20717 36533 20729 36536
rect 20763 36564 20775 36567
rect 20806 36564 20812 36576
rect 20763 36536 20812 36564
rect 20763 36533 20775 36536
rect 20717 36527 20775 36533
rect 20806 36524 20812 36536
rect 20864 36524 20870 36576
rect 1104 36474 49864 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 32950 36474
rect 33002 36422 33014 36474
rect 33066 36422 33078 36474
rect 33130 36422 33142 36474
rect 33194 36422 33206 36474
rect 33258 36422 42950 36474
rect 43002 36422 43014 36474
rect 43066 36422 43078 36474
rect 43130 36422 43142 36474
rect 43194 36422 43206 36474
rect 43258 36422 49864 36474
rect 1104 36400 49864 36422
rect 5534 36320 5540 36372
rect 5592 36360 5598 36372
rect 7837 36363 7895 36369
rect 7837 36360 7849 36363
rect 5592 36332 7849 36360
rect 5592 36320 5598 36332
rect 7837 36329 7849 36332
rect 7883 36329 7895 36363
rect 10594 36360 10600 36372
rect 7837 36323 7895 36329
rect 7944 36332 10600 36360
rect 6546 36252 6552 36304
rect 6604 36292 6610 36304
rect 7944 36292 7972 36332
rect 10594 36320 10600 36332
rect 10652 36320 10658 36372
rect 11790 36320 11796 36372
rect 11848 36320 11854 36372
rect 12437 36363 12495 36369
rect 12437 36329 12449 36363
rect 12483 36360 12495 36363
rect 12802 36360 12808 36372
rect 12483 36332 12808 36360
rect 12483 36329 12495 36332
rect 12437 36323 12495 36329
rect 12802 36320 12808 36332
rect 12860 36320 12866 36372
rect 14734 36320 14740 36372
rect 14792 36360 14798 36372
rect 16117 36363 16175 36369
rect 16117 36360 16129 36363
rect 14792 36332 16129 36360
rect 14792 36320 14798 36332
rect 16117 36329 16129 36332
rect 16163 36329 16175 36363
rect 16117 36323 16175 36329
rect 17402 36320 17408 36372
rect 17460 36360 17466 36372
rect 22186 36360 22192 36372
rect 17460 36332 22192 36360
rect 17460 36320 17466 36332
rect 22186 36320 22192 36332
rect 22244 36320 22250 36372
rect 6604 36264 7972 36292
rect 6604 36252 6610 36264
rect 19058 36252 19064 36304
rect 19116 36292 19122 36304
rect 19334 36292 19340 36304
rect 19116 36264 19340 36292
rect 19116 36252 19122 36264
rect 19334 36252 19340 36264
rect 19392 36252 19398 36304
rect 21910 36252 21916 36304
rect 21968 36252 21974 36304
rect 6089 36227 6147 36233
rect 6089 36193 6101 36227
rect 6135 36224 6147 36227
rect 6454 36224 6460 36236
rect 6135 36196 6460 36224
rect 6135 36193 6147 36196
rect 6089 36187 6147 36193
rect 6454 36184 6460 36196
rect 6512 36224 6518 36236
rect 7098 36224 7104 36236
rect 6512 36196 7104 36224
rect 6512 36184 6518 36196
rect 7098 36184 7104 36196
rect 7156 36224 7162 36236
rect 7193 36227 7251 36233
rect 7193 36224 7205 36227
rect 7156 36196 7205 36224
rect 7156 36184 7162 36196
rect 7193 36193 7205 36196
rect 7239 36193 7251 36227
rect 7193 36187 7251 36193
rect 7926 36184 7932 36236
rect 7984 36224 7990 36236
rect 8297 36227 8355 36233
rect 8297 36224 8309 36227
rect 7984 36196 8309 36224
rect 7984 36184 7990 36196
rect 8297 36193 8309 36196
rect 8343 36193 8355 36227
rect 8297 36187 8355 36193
rect 8478 36184 8484 36236
rect 8536 36224 8542 36236
rect 8938 36224 8944 36236
rect 8536 36196 8944 36224
rect 8536 36184 8542 36196
rect 8938 36184 8944 36196
rect 8996 36224 9002 36236
rect 11149 36227 11207 36233
rect 11149 36224 11161 36227
rect 8996 36196 11161 36224
rect 8996 36184 9002 36196
rect 11149 36193 11161 36196
rect 11195 36224 11207 36227
rect 13081 36227 13139 36233
rect 11195 36196 12434 36224
rect 11195 36193 11207 36196
rect 11149 36187 11207 36193
rect 1765 36159 1823 36165
rect 1765 36125 1777 36159
rect 1811 36156 1823 36159
rect 4062 36156 4068 36168
rect 1811 36128 4068 36156
rect 1811 36125 1823 36128
rect 1765 36119 1823 36125
rect 4062 36116 4068 36128
rect 4120 36116 4126 36168
rect 5813 36159 5871 36165
rect 5813 36125 5825 36159
rect 5859 36156 5871 36159
rect 6362 36156 6368 36168
rect 5859 36128 6368 36156
rect 5859 36125 5871 36128
rect 5813 36119 5871 36125
rect 6362 36116 6368 36128
rect 6420 36116 6426 36168
rect 6638 36156 6644 36168
rect 6472 36128 6644 36156
rect 6472 36100 6500 36128
rect 6638 36116 6644 36128
rect 6696 36116 6702 36168
rect 6914 36116 6920 36168
rect 6972 36156 6978 36168
rect 9030 36156 9036 36168
rect 6972 36128 9036 36156
rect 6972 36116 6978 36128
rect 9030 36116 9036 36128
rect 9088 36156 9094 36168
rect 9125 36159 9183 36165
rect 9125 36156 9137 36159
rect 9088 36128 9137 36156
rect 9088 36116 9094 36128
rect 9125 36125 9137 36128
rect 9171 36125 9183 36159
rect 12406 36156 12434 36196
rect 13081 36193 13093 36227
rect 13127 36224 13139 36227
rect 13722 36224 13728 36236
rect 13127 36196 13728 36224
rect 13127 36193 13139 36196
rect 13081 36187 13139 36193
rect 13722 36184 13728 36196
rect 13780 36184 13786 36236
rect 14645 36227 14703 36233
rect 14645 36193 14657 36227
rect 14691 36224 14703 36227
rect 16022 36224 16028 36236
rect 14691 36196 16028 36224
rect 14691 36193 14703 36196
rect 14645 36187 14703 36193
rect 16022 36184 16028 36196
rect 16080 36184 16086 36236
rect 16850 36184 16856 36236
rect 16908 36224 16914 36236
rect 18693 36227 18751 36233
rect 18693 36224 18705 36227
rect 16908 36196 18705 36224
rect 16908 36184 16914 36196
rect 18693 36193 18705 36196
rect 18739 36193 18751 36227
rect 18693 36187 18751 36193
rect 20162 36184 20168 36236
rect 20220 36184 20226 36236
rect 13906 36156 13912 36168
rect 12406 36128 13912 36156
rect 9125 36119 9183 36125
rect 13906 36116 13912 36128
rect 13964 36116 13970 36168
rect 14274 36116 14280 36168
rect 14332 36156 14338 36168
rect 14369 36159 14427 36165
rect 14369 36156 14381 36159
rect 14332 36128 14381 36156
rect 14332 36116 14338 36128
rect 14369 36125 14381 36128
rect 14415 36125 14427 36159
rect 14369 36119 14427 36125
rect 18414 36116 18420 36168
rect 18472 36156 18478 36168
rect 18509 36159 18567 36165
rect 18509 36156 18521 36159
rect 18472 36128 18521 36156
rect 18472 36116 18478 36128
rect 18509 36125 18521 36128
rect 18555 36125 18567 36159
rect 18509 36119 18567 36125
rect 2774 36048 2780 36100
rect 2832 36048 2838 36100
rect 5905 36091 5963 36097
rect 5905 36057 5917 36091
rect 5951 36088 5963 36091
rect 6270 36088 6276 36100
rect 5951 36060 6276 36088
rect 5951 36057 5963 36060
rect 5905 36051 5963 36057
rect 6270 36048 6276 36060
rect 6328 36048 6334 36100
rect 6454 36048 6460 36100
rect 6512 36048 6518 36100
rect 7006 36048 7012 36100
rect 7064 36048 7070 36100
rect 7101 36091 7159 36097
rect 7101 36057 7113 36091
rect 7147 36088 7159 36091
rect 7374 36088 7380 36100
rect 7147 36060 7380 36088
rect 7147 36057 7159 36060
rect 7101 36051 7159 36057
rect 7374 36048 7380 36060
rect 7432 36048 7438 36100
rect 7650 36048 7656 36100
rect 7708 36088 7714 36100
rect 9401 36091 9459 36097
rect 9401 36088 9413 36091
rect 7708 36060 9413 36088
rect 7708 36048 7714 36060
rect 9401 36057 9413 36060
rect 9447 36057 9459 36091
rect 9401 36051 9459 36057
rect 10410 36048 10416 36100
rect 10468 36048 10474 36100
rect 11238 36048 11244 36100
rect 11296 36088 11302 36100
rect 11296 36060 15056 36088
rect 11296 36048 11302 36060
rect 5445 36023 5503 36029
rect 5445 35989 5457 36023
rect 5491 36020 5503 36023
rect 5718 36020 5724 36032
rect 5491 35992 5724 36020
rect 5491 35989 5503 35992
rect 5445 35983 5503 35989
rect 5718 35980 5724 35992
rect 5776 35980 5782 36032
rect 6641 36023 6699 36029
rect 6641 35989 6653 36023
rect 6687 36020 6699 36023
rect 6822 36020 6828 36032
rect 6687 35992 6828 36020
rect 6687 35989 6699 35992
rect 6641 35983 6699 35989
rect 6822 35980 6828 35992
rect 6880 35980 6886 36032
rect 7926 35980 7932 36032
rect 7984 36020 7990 36032
rect 8205 36023 8263 36029
rect 8205 36020 8217 36023
rect 7984 35992 8217 36020
rect 7984 35980 7990 35992
rect 8205 35989 8217 35992
rect 8251 35989 8263 36023
rect 8205 35983 8263 35989
rect 12802 35980 12808 36032
rect 12860 35980 12866 36032
rect 12897 36023 12955 36029
rect 12897 35989 12909 36023
rect 12943 36020 12955 36023
rect 13354 36020 13360 36032
rect 12943 35992 13360 36020
rect 12943 35989 12955 35992
rect 12897 35983 12955 35989
rect 13354 35980 13360 35992
rect 13412 35980 13418 36032
rect 15028 36020 15056 36060
rect 15378 36048 15384 36100
rect 15436 36048 15442 36100
rect 17589 36091 17647 36097
rect 17589 36088 17601 36091
rect 16040 36060 17601 36088
rect 16040 36020 16068 36060
rect 17589 36057 17601 36060
rect 17635 36088 17647 36091
rect 18601 36091 18659 36097
rect 18601 36088 18613 36091
rect 17635 36060 18613 36088
rect 17635 36057 17647 36060
rect 17589 36051 17647 36057
rect 18601 36057 18613 36060
rect 18647 36057 18659 36091
rect 18601 36051 18659 36057
rect 15028 35992 16068 36020
rect 16206 35980 16212 36032
rect 16264 36020 16270 36032
rect 18141 36023 18199 36029
rect 18141 36020 18153 36023
rect 16264 35992 18153 36020
rect 16264 35980 16270 35992
rect 18141 35989 18153 35992
rect 18187 35989 18199 36023
rect 18616 36020 18644 36051
rect 20438 36048 20444 36100
rect 20496 36048 20502 36100
rect 20714 36048 20720 36100
rect 20772 36088 20778 36100
rect 23382 36088 23388 36100
rect 20772 36060 20930 36088
rect 21836 36060 23388 36088
rect 20772 36048 20778 36060
rect 21836 36020 21864 36060
rect 23382 36048 23388 36060
rect 23440 36048 23446 36100
rect 18616 35992 21864 36020
rect 18141 35983 18199 35989
rect 1104 35930 49864 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 27950 35930
rect 28002 35878 28014 35930
rect 28066 35878 28078 35930
rect 28130 35878 28142 35930
rect 28194 35878 28206 35930
rect 28258 35878 37950 35930
rect 38002 35878 38014 35930
rect 38066 35878 38078 35930
rect 38130 35878 38142 35930
rect 38194 35878 38206 35930
rect 38258 35878 47950 35930
rect 48002 35878 48014 35930
rect 48066 35878 48078 35930
rect 48130 35878 48142 35930
rect 48194 35878 48206 35930
rect 48258 35878 49864 35930
rect 1104 35856 49864 35878
rect 5718 35776 5724 35828
rect 5776 35816 5782 35828
rect 7193 35819 7251 35825
rect 7193 35816 7205 35819
rect 5776 35788 7205 35816
rect 5776 35776 5782 35788
rect 7193 35785 7205 35788
rect 7239 35785 7251 35819
rect 7193 35779 7251 35785
rect 7742 35776 7748 35828
rect 7800 35816 7806 35828
rect 8021 35819 8079 35825
rect 8021 35816 8033 35819
rect 7800 35788 8033 35816
rect 7800 35776 7806 35788
rect 8021 35785 8033 35788
rect 8067 35785 8079 35819
rect 9585 35819 9643 35825
rect 8021 35779 8079 35785
rect 8128 35788 8616 35816
rect 5629 35751 5687 35757
rect 5629 35717 5641 35751
rect 5675 35748 5687 35751
rect 5994 35748 6000 35760
rect 5675 35720 6000 35748
rect 5675 35717 5687 35720
rect 5629 35711 5687 35717
rect 5994 35708 6000 35720
rect 6052 35708 6058 35760
rect 8128 35748 8156 35788
rect 7392 35720 8156 35748
rect 8389 35751 8447 35757
rect 5350 35640 5356 35692
rect 5408 35680 5414 35692
rect 7285 35683 7343 35689
rect 7285 35680 7297 35683
rect 5408 35652 7297 35680
rect 5408 35640 5414 35652
rect 7285 35649 7297 35652
rect 7331 35649 7343 35683
rect 7285 35643 7343 35649
rect 5721 35615 5779 35621
rect 5721 35581 5733 35615
rect 5767 35581 5779 35615
rect 5721 35575 5779 35581
rect 5905 35615 5963 35621
rect 5905 35581 5917 35615
rect 5951 35612 5963 35615
rect 6546 35612 6552 35624
rect 5951 35584 6552 35612
rect 5951 35581 5963 35584
rect 5905 35575 5963 35581
rect 4798 35504 4804 35556
rect 4856 35544 4862 35556
rect 5736 35544 5764 35575
rect 6546 35572 6552 35584
rect 6604 35572 6610 35624
rect 7392 35544 7420 35720
rect 8389 35717 8401 35751
rect 8435 35748 8447 35751
rect 8478 35748 8484 35760
rect 8435 35720 8484 35748
rect 8435 35717 8447 35720
rect 8389 35711 8447 35717
rect 8478 35708 8484 35720
rect 8536 35708 8542 35760
rect 8588 35748 8616 35788
rect 9585 35785 9597 35819
rect 9631 35816 9643 35819
rect 9766 35816 9772 35828
rect 9631 35788 9772 35816
rect 9631 35785 9643 35788
rect 9585 35779 9643 35785
rect 9766 35776 9772 35788
rect 9824 35776 9830 35828
rect 10042 35776 10048 35828
rect 10100 35816 10106 35828
rect 10413 35819 10471 35825
rect 10413 35816 10425 35819
rect 10100 35788 10425 35816
rect 10100 35776 10106 35788
rect 10413 35785 10425 35788
rect 10459 35785 10471 35819
rect 10413 35779 10471 35785
rect 13538 35776 13544 35828
rect 13596 35816 13602 35828
rect 14277 35819 14335 35825
rect 14277 35816 14289 35819
rect 13596 35788 14289 35816
rect 13596 35776 13602 35788
rect 14277 35785 14289 35788
rect 14323 35785 14335 35819
rect 14277 35779 14335 35785
rect 16025 35819 16083 35825
rect 16025 35785 16037 35819
rect 16071 35816 16083 35819
rect 16574 35816 16580 35828
rect 16071 35788 16580 35816
rect 16071 35785 16083 35788
rect 16025 35779 16083 35785
rect 16574 35776 16580 35788
rect 16632 35776 16638 35828
rect 17405 35819 17463 35825
rect 17405 35785 17417 35819
rect 17451 35816 17463 35819
rect 17770 35816 17776 35828
rect 17451 35788 17776 35816
rect 17451 35785 17463 35788
rect 17405 35779 17463 35785
rect 17770 35776 17776 35788
rect 17828 35776 17834 35828
rect 18877 35819 18935 35825
rect 18877 35785 18889 35819
rect 18923 35816 18935 35819
rect 19426 35816 19432 35828
rect 18923 35788 19432 35816
rect 18923 35785 18935 35788
rect 18877 35779 18935 35785
rect 10134 35748 10140 35760
rect 8588 35720 10140 35748
rect 10134 35708 10140 35720
rect 10192 35708 10198 35760
rect 10873 35751 10931 35757
rect 10873 35717 10885 35751
rect 10919 35748 10931 35751
rect 11514 35748 11520 35760
rect 10919 35720 11520 35748
rect 10919 35717 10931 35720
rect 10873 35711 10931 35717
rect 11514 35708 11520 35720
rect 11572 35708 11578 35760
rect 12710 35708 12716 35760
rect 12768 35748 12774 35760
rect 12768 35720 13294 35748
rect 12768 35708 12774 35720
rect 14458 35708 14464 35760
rect 14516 35748 14522 35760
rect 17313 35751 17371 35757
rect 17313 35748 17325 35751
rect 14516 35720 17325 35748
rect 14516 35708 14522 35720
rect 17313 35717 17325 35720
rect 17359 35717 17371 35751
rect 17313 35711 17371 35717
rect 7558 35640 7564 35692
rect 7616 35680 7622 35692
rect 9677 35683 9735 35689
rect 9677 35680 9689 35683
rect 7616 35652 9689 35680
rect 7616 35640 7622 35652
rect 9677 35649 9689 35652
rect 9723 35649 9735 35683
rect 9677 35643 9735 35649
rect 10781 35683 10839 35689
rect 10781 35649 10793 35683
rect 10827 35680 10839 35683
rect 11977 35683 12035 35689
rect 11977 35680 11989 35683
rect 10827 35652 11989 35680
rect 10827 35649 10839 35652
rect 10781 35643 10839 35649
rect 11977 35649 11989 35652
rect 12023 35649 12035 35683
rect 11977 35643 12035 35649
rect 14090 35640 14096 35692
rect 14148 35680 14154 35692
rect 15933 35683 15991 35689
rect 15933 35680 15945 35683
rect 14148 35652 15945 35680
rect 14148 35640 14154 35652
rect 15933 35649 15945 35652
rect 15979 35649 15991 35683
rect 18892 35680 18920 35779
rect 19426 35776 19432 35788
rect 19484 35776 19490 35828
rect 22278 35816 22284 35828
rect 19996 35788 22284 35816
rect 19996 35757 20024 35788
rect 22278 35776 22284 35788
rect 22336 35776 22342 35828
rect 18969 35751 19027 35757
rect 18969 35717 18981 35751
rect 19015 35748 19027 35751
rect 19981 35751 20039 35757
rect 19015 35720 19196 35748
rect 19015 35717 19027 35720
rect 18969 35711 19027 35717
rect 15933 35643 15991 35649
rect 16132 35652 18920 35680
rect 7466 35572 7472 35624
rect 7524 35572 7530 35624
rect 8481 35615 8539 35621
rect 8481 35581 8493 35615
rect 8527 35581 8539 35615
rect 8481 35575 8539 35581
rect 4856 35516 7420 35544
rect 8496 35544 8524 35575
rect 8570 35572 8576 35624
rect 8628 35572 8634 35624
rect 8662 35572 8668 35624
rect 8720 35612 8726 35624
rect 9769 35615 9827 35621
rect 9769 35612 9781 35615
rect 8720 35584 9781 35612
rect 8720 35572 8726 35584
rect 9769 35581 9781 35584
rect 9815 35612 9827 35615
rect 10502 35612 10508 35624
rect 9815 35584 10508 35612
rect 9815 35581 9827 35584
rect 9769 35575 9827 35581
rect 10502 35572 10508 35584
rect 10560 35572 10566 35624
rect 11057 35615 11115 35621
rect 11057 35581 11069 35615
rect 11103 35612 11115 35615
rect 12342 35612 12348 35624
rect 11103 35584 12348 35612
rect 11103 35581 11115 35584
rect 11057 35575 11115 35581
rect 12342 35572 12348 35584
rect 12400 35572 12406 35624
rect 12529 35615 12587 35621
rect 12529 35581 12541 35615
rect 12575 35612 12587 35615
rect 12805 35615 12863 35621
rect 12575 35584 12664 35612
rect 12575 35581 12587 35584
rect 12529 35575 12587 35581
rect 11238 35544 11244 35556
rect 8496 35516 11244 35544
rect 4856 35504 4862 35516
rect 11238 35504 11244 35516
rect 11296 35504 11302 35556
rect 5261 35479 5319 35485
rect 5261 35445 5273 35479
rect 5307 35476 5319 35479
rect 6730 35476 6736 35488
rect 5307 35448 6736 35476
rect 5307 35445 5319 35448
rect 5261 35439 5319 35445
rect 6730 35436 6736 35448
rect 6788 35436 6794 35488
rect 6825 35479 6883 35485
rect 6825 35445 6837 35479
rect 6871 35476 6883 35479
rect 9122 35476 9128 35488
rect 6871 35448 9128 35476
rect 6871 35445 6883 35448
rect 6825 35439 6883 35445
rect 9122 35436 9128 35448
rect 9180 35436 9186 35488
rect 9214 35436 9220 35488
rect 9272 35436 9278 35488
rect 12636 35476 12664 35584
rect 12805 35581 12817 35615
rect 12851 35612 12863 35615
rect 13538 35612 13544 35624
rect 12851 35584 13544 35612
rect 12851 35581 12863 35584
rect 12805 35575 12863 35581
rect 13538 35572 13544 35584
rect 13596 35572 13602 35624
rect 14642 35572 14648 35624
rect 14700 35612 14706 35624
rect 16132 35612 16160 35652
rect 14700 35584 16160 35612
rect 16209 35615 16267 35621
rect 14700 35572 14706 35584
rect 16209 35581 16221 35615
rect 16255 35612 16267 35615
rect 17402 35612 17408 35624
rect 16255 35584 17408 35612
rect 16255 35581 16267 35584
rect 16209 35575 16267 35581
rect 17402 35572 17408 35584
rect 17460 35572 17466 35624
rect 17589 35615 17647 35621
rect 17589 35581 17601 35615
rect 17635 35612 17647 35615
rect 17770 35612 17776 35624
rect 17635 35584 17776 35612
rect 17635 35581 17647 35584
rect 17589 35575 17647 35581
rect 17770 35572 17776 35584
rect 17828 35572 17834 35624
rect 17862 35572 17868 35624
rect 17920 35612 17926 35624
rect 19061 35615 19119 35621
rect 19061 35612 19073 35615
rect 17920 35584 19073 35612
rect 17920 35572 17926 35584
rect 19061 35581 19073 35584
rect 19107 35581 19119 35615
rect 19061 35575 19119 35581
rect 15838 35504 15844 35556
rect 15896 35544 15902 35556
rect 16945 35547 17003 35553
rect 16945 35544 16957 35547
rect 15896 35516 16957 35544
rect 15896 35504 15902 35516
rect 16945 35513 16957 35516
rect 16991 35513 17003 35547
rect 16945 35507 17003 35513
rect 17034 35504 17040 35556
rect 17092 35544 17098 35556
rect 19168 35544 19196 35720
rect 19981 35717 19993 35751
rect 20027 35717 20039 35751
rect 19981 35711 20039 35717
rect 20714 35708 20720 35760
rect 20772 35708 20778 35760
rect 22002 35708 22008 35760
rect 22060 35708 22066 35760
rect 19705 35615 19763 35621
rect 19705 35581 19717 35615
rect 19751 35581 19763 35615
rect 22833 35615 22891 35621
rect 22833 35612 22845 35615
rect 19705 35575 19763 35581
rect 22066 35584 22845 35612
rect 19334 35544 19340 35556
rect 17092 35516 19340 35544
rect 17092 35504 17098 35516
rect 19334 35504 19340 35516
rect 19392 35504 19398 35556
rect 19720 35488 19748 35575
rect 22066 35544 22094 35584
rect 22833 35581 22845 35584
rect 22879 35612 22891 35615
rect 24118 35612 24124 35624
rect 22879 35584 24124 35612
rect 22879 35581 22891 35584
rect 22833 35575 22891 35581
rect 24118 35572 24124 35584
rect 24176 35572 24182 35624
rect 21008 35516 22094 35544
rect 14274 35476 14280 35488
rect 12636 35448 14280 35476
rect 14274 35436 14280 35448
rect 14332 35436 14338 35488
rect 15565 35479 15623 35485
rect 15565 35445 15577 35479
rect 15611 35476 15623 35479
rect 17310 35476 17316 35488
rect 15611 35448 17316 35476
rect 15611 35445 15623 35448
rect 15565 35439 15623 35445
rect 17310 35436 17316 35448
rect 17368 35436 17374 35488
rect 18414 35436 18420 35488
rect 18472 35476 18478 35488
rect 18509 35479 18567 35485
rect 18509 35476 18521 35479
rect 18472 35448 18521 35476
rect 18472 35436 18478 35448
rect 18509 35445 18521 35448
rect 18555 35445 18567 35479
rect 18509 35439 18567 35445
rect 19702 35436 19708 35488
rect 19760 35476 19766 35488
rect 21008 35476 21036 35516
rect 19760 35448 21036 35476
rect 21453 35479 21511 35485
rect 19760 35436 19766 35448
rect 21453 35445 21465 35479
rect 21499 35476 21511 35479
rect 21542 35476 21548 35488
rect 21499 35448 21548 35476
rect 21499 35445 21511 35448
rect 21453 35439 21511 35445
rect 21542 35436 21548 35448
rect 21600 35436 21606 35488
rect 1104 35386 49864 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 32950 35386
rect 33002 35334 33014 35386
rect 33066 35334 33078 35386
rect 33130 35334 33142 35386
rect 33194 35334 33206 35386
rect 33258 35334 42950 35386
rect 43002 35334 43014 35386
rect 43066 35334 43078 35386
rect 43130 35334 43142 35386
rect 43194 35334 43206 35386
rect 43258 35334 49864 35386
rect 1104 35312 49864 35334
rect 7834 35232 7840 35284
rect 7892 35232 7898 35284
rect 10502 35232 10508 35284
rect 10560 35272 10566 35284
rect 11425 35275 11483 35281
rect 11425 35272 11437 35275
rect 10560 35244 11437 35272
rect 10560 35232 10566 35244
rect 11425 35241 11437 35244
rect 11471 35241 11483 35275
rect 11425 35235 11483 35241
rect 12529 35275 12587 35281
rect 12529 35241 12541 35275
rect 12575 35272 12587 35275
rect 12802 35272 12808 35284
rect 12575 35244 12808 35272
rect 12575 35241 12587 35244
rect 12529 35235 12587 35241
rect 12802 35232 12808 35244
rect 12860 35232 12866 35284
rect 12989 35275 13047 35281
rect 12989 35241 13001 35275
rect 13035 35272 13047 35275
rect 13446 35272 13452 35284
rect 13035 35244 13452 35272
rect 13035 35241 13047 35244
rect 12989 35235 13047 35241
rect 13446 35232 13452 35244
rect 13504 35232 13510 35284
rect 15565 35275 15623 35281
rect 15565 35241 15577 35275
rect 15611 35272 15623 35275
rect 16298 35272 16304 35284
rect 15611 35244 16304 35272
rect 15611 35241 15623 35244
rect 15565 35235 15623 35241
rect 16298 35232 16304 35244
rect 16356 35232 16362 35284
rect 17402 35232 17408 35284
rect 17460 35272 17466 35284
rect 18877 35275 18935 35281
rect 18877 35272 18889 35275
rect 17460 35244 18889 35272
rect 17460 35232 17466 35244
rect 18877 35241 18889 35244
rect 18923 35241 18935 35275
rect 18877 35235 18935 35241
rect 5445 35207 5503 35213
rect 5445 35173 5457 35207
rect 5491 35204 5503 35207
rect 7650 35204 7656 35216
rect 5491 35176 7656 35204
rect 5491 35173 5503 35176
rect 5445 35167 5503 35173
rect 7650 35164 7656 35176
rect 7708 35164 7714 35216
rect 8202 35164 8208 35216
rect 8260 35204 8266 35216
rect 9306 35204 9312 35216
rect 8260 35176 9312 35204
rect 8260 35164 8266 35176
rect 9306 35164 9312 35176
rect 9364 35164 9370 35216
rect 10962 35164 10968 35216
rect 11020 35204 11026 35216
rect 17034 35204 17040 35216
rect 11020 35176 17040 35204
rect 11020 35164 11026 35176
rect 17034 35164 17040 35176
rect 17092 35164 17098 35216
rect 19334 35164 19340 35216
rect 19392 35204 19398 35216
rect 23750 35204 23756 35216
rect 19392 35176 23756 35204
rect 19392 35164 19398 35176
rect 23750 35164 23756 35176
rect 23808 35164 23814 35216
rect 1302 35096 1308 35148
rect 1360 35136 1366 35148
rect 2041 35139 2099 35145
rect 2041 35136 2053 35139
rect 1360 35108 2053 35136
rect 1360 35096 1366 35108
rect 2041 35105 2053 35108
rect 2087 35105 2099 35139
rect 2041 35099 2099 35105
rect 5902 35096 5908 35148
rect 5960 35096 5966 35148
rect 6089 35139 6147 35145
rect 6089 35105 6101 35139
rect 6135 35105 6147 35139
rect 6089 35099 6147 35105
rect 1765 35071 1823 35077
rect 1765 35037 1777 35071
rect 1811 35068 1823 35071
rect 3970 35068 3976 35080
rect 1811 35040 3976 35068
rect 1811 35037 1823 35040
rect 1765 35031 1823 35037
rect 3970 35028 3976 35040
rect 4028 35028 4034 35080
rect 5810 35028 5816 35080
rect 5868 35028 5874 35080
rect 6104 35000 6132 35099
rect 6730 35096 6736 35148
rect 6788 35136 6794 35148
rect 7101 35139 7159 35145
rect 7101 35136 7113 35139
rect 6788 35108 7113 35136
rect 6788 35096 6794 35108
rect 7101 35105 7113 35108
rect 7147 35105 7159 35139
rect 7101 35099 7159 35105
rect 7190 35096 7196 35148
rect 7248 35096 7254 35148
rect 7742 35096 7748 35148
rect 7800 35136 7806 35148
rect 8389 35139 8447 35145
rect 8389 35136 8401 35139
rect 7800 35108 8401 35136
rect 7800 35096 7806 35108
rect 8389 35105 8401 35108
rect 8435 35105 8447 35139
rect 8389 35099 8447 35105
rect 9677 35139 9735 35145
rect 9677 35105 9689 35139
rect 9723 35136 9735 35139
rect 12066 35136 12072 35148
rect 9723 35108 12072 35136
rect 9723 35105 9735 35108
rect 9677 35099 9735 35105
rect 12066 35096 12072 35108
rect 12124 35096 12130 35148
rect 13538 35096 13544 35148
rect 13596 35096 13602 35148
rect 14918 35096 14924 35148
rect 14976 35096 14982 35148
rect 16117 35139 16175 35145
rect 16117 35105 16129 35139
rect 16163 35136 16175 35139
rect 16666 35136 16672 35148
rect 16163 35108 16672 35136
rect 16163 35105 16175 35108
rect 16117 35099 16175 35105
rect 16666 35096 16672 35108
rect 16724 35096 16730 35148
rect 17129 35139 17187 35145
rect 17129 35105 17141 35139
rect 17175 35136 17187 35139
rect 19702 35136 19708 35148
rect 17175 35108 19708 35136
rect 17175 35105 17187 35108
rect 17129 35099 17187 35105
rect 19702 35096 19708 35108
rect 19760 35096 19766 35148
rect 20622 35096 20628 35148
rect 20680 35096 20686 35148
rect 21726 35096 21732 35148
rect 21784 35096 21790 35148
rect 21818 35096 21824 35148
rect 21876 35096 21882 35148
rect 7009 35071 7067 35077
rect 7009 35037 7021 35071
rect 7055 35068 7067 35071
rect 8294 35068 8300 35080
rect 7055 35040 8300 35068
rect 7055 35037 7067 35040
rect 7009 35031 7067 35037
rect 8294 35028 8300 35040
rect 8352 35028 8358 35080
rect 13354 35028 13360 35080
rect 13412 35028 13418 35080
rect 13449 35071 13507 35077
rect 13449 35037 13461 35071
rect 13495 35068 13507 35071
rect 14642 35068 14648 35080
rect 13495 35040 14648 35068
rect 13495 35037 13507 35040
rect 13449 35031 13507 35037
rect 14642 35028 14648 35040
rect 14700 35028 14706 35080
rect 14829 35071 14887 35077
rect 14829 35037 14841 35071
rect 14875 35068 14887 35071
rect 16206 35068 16212 35080
rect 14875 35040 16212 35068
rect 14875 35037 14887 35040
rect 14829 35031 14887 35037
rect 16206 35028 16212 35040
rect 16264 35028 16270 35080
rect 20441 35071 20499 35077
rect 20441 35037 20453 35071
rect 20487 35068 20499 35071
rect 21174 35068 21180 35080
rect 20487 35040 21180 35068
rect 20487 35037 20499 35040
rect 20441 35031 20499 35037
rect 21174 35028 21180 35040
rect 21232 35028 21238 35080
rect 21634 35028 21640 35080
rect 21692 35028 21698 35080
rect 7190 35000 7196 35012
rect 6104 34972 7196 35000
rect 7190 34960 7196 34972
rect 7248 34960 7254 35012
rect 8110 34960 8116 35012
rect 8168 35000 8174 35012
rect 9953 35003 10011 35009
rect 8168 34972 8340 35000
rect 8168 34960 8174 34972
rect 6641 34935 6699 34941
rect 6641 34901 6653 34935
rect 6687 34932 6699 34935
rect 6914 34932 6920 34944
rect 6687 34904 6920 34932
rect 6687 34901 6699 34904
rect 6641 34895 6699 34901
rect 6914 34892 6920 34904
rect 6972 34892 6978 34944
rect 7006 34892 7012 34944
rect 7064 34932 7070 34944
rect 8128 34932 8156 34960
rect 7064 34904 8156 34932
rect 7064 34892 7070 34904
rect 8202 34892 8208 34944
rect 8260 34892 8266 34944
rect 8312 34941 8340 34972
rect 9953 34969 9965 35003
rect 9999 35000 10011 35003
rect 10226 35000 10232 35012
rect 9999 34972 10232 35000
rect 9999 34969 10011 34972
rect 9953 34963 10011 34969
rect 10226 34960 10232 34972
rect 10284 34960 10290 35012
rect 10410 34960 10416 35012
rect 10468 34960 10474 35012
rect 12802 34960 12808 35012
rect 12860 35000 12866 35012
rect 14737 35003 14795 35009
rect 14737 35000 14749 35003
rect 12860 34972 14749 35000
rect 12860 34960 12866 34972
rect 14737 34969 14749 34972
rect 14783 34969 14795 35003
rect 14737 34963 14795 34969
rect 15856 34972 16436 35000
rect 8297 34935 8355 34941
rect 8297 34901 8309 34935
rect 8343 34901 8355 34935
rect 8297 34895 8355 34901
rect 8386 34892 8392 34944
rect 8444 34932 8450 34944
rect 9674 34932 9680 34944
rect 8444 34904 9680 34932
rect 8444 34892 8450 34904
rect 9674 34892 9680 34904
rect 9732 34892 9738 34944
rect 14369 34935 14427 34941
rect 14369 34901 14381 34935
rect 14415 34932 14427 34935
rect 15856 34932 15884 34972
rect 14415 34904 15884 34932
rect 14415 34901 14427 34904
rect 14369 34895 14427 34901
rect 15930 34892 15936 34944
rect 15988 34892 15994 34944
rect 16025 34935 16083 34941
rect 16025 34901 16037 34935
rect 16071 34932 16083 34935
rect 16206 34932 16212 34944
rect 16071 34904 16212 34932
rect 16071 34901 16083 34904
rect 16025 34895 16083 34901
rect 16206 34892 16212 34904
rect 16264 34892 16270 34944
rect 16408 34932 16436 34972
rect 17310 34960 17316 35012
rect 17368 35000 17374 35012
rect 17405 35003 17463 35009
rect 17405 35000 17417 35003
rect 17368 34972 17417 35000
rect 17368 34960 17374 34972
rect 17405 34969 17417 34972
rect 17451 34969 17463 35003
rect 17405 34963 17463 34969
rect 17862 34960 17868 35012
rect 17920 34960 17926 35012
rect 20533 35003 20591 35009
rect 20533 34969 20545 35003
rect 20579 35000 20591 35003
rect 21358 35000 21364 35012
rect 20579 34972 21364 35000
rect 20579 34969 20591 34972
rect 20533 34963 20591 34969
rect 21358 34960 21364 34972
rect 21416 34960 21422 35012
rect 17494 34932 17500 34944
rect 16408 34904 17500 34932
rect 17494 34892 17500 34904
rect 17552 34892 17558 34944
rect 18322 34892 18328 34944
rect 18380 34932 18386 34944
rect 20073 34935 20131 34941
rect 20073 34932 20085 34935
rect 18380 34904 20085 34932
rect 18380 34892 18386 34904
rect 20073 34901 20085 34904
rect 20119 34901 20131 34935
rect 20073 34895 20131 34901
rect 21266 34892 21272 34944
rect 21324 34892 21330 34944
rect 1104 34842 49864 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 27950 34842
rect 28002 34790 28014 34842
rect 28066 34790 28078 34842
rect 28130 34790 28142 34842
rect 28194 34790 28206 34842
rect 28258 34790 37950 34842
rect 38002 34790 38014 34842
rect 38066 34790 38078 34842
rect 38130 34790 38142 34842
rect 38194 34790 38206 34842
rect 38258 34790 47950 34842
rect 48002 34790 48014 34842
rect 48066 34790 48078 34842
rect 48130 34790 48142 34842
rect 48194 34790 48206 34842
rect 48258 34790 49864 34842
rect 1104 34768 49864 34790
rect 8386 34728 8392 34740
rect 2746 34700 8392 34728
rect 2746 34660 2774 34700
rect 8386 34688 8392 34700
rect 8444 34688 8450 34740
rect 8754 34688 8760 34740
rect 8812 34688 8818 34740
rect 9217 34731 9275 34737
rect 9217 34697 9229 34731
rect 9263 34728 9275 34731
rect 10962 34728 10968 34740
rect 9263 34700 10968 34728
rect 9263 34697 9275 34700
rect 9217 34691 9275 34697
rect 10962 34688 10968 34700
rect 11020 34688 11026 34740
rect 16114 34728 16120 34740
rect 11072 34700 13676 34728
rect 1780 34632 2774 34660
rect 1780 34601 1808 34632
rect 6638 34620 6644 34672
rect 6696 34660 6702 34672
rect 10413 34663 10471 34669
rect 10413 34660 10425 34663
rect 6696 34632 10425 34660
rect 6696 34620 6702 34632
rect 10413 34629 10425 34632
rect 10459 34660 10471 34663
rect 11072 34660 11100 34700
rect 10459 34632 11100 34660
rect 10459 34629 10471 34632
rect 10413 34623 10471 34629
rect 12342 34620 12348 34672
rect 12400 34620 12406 34672
rect 12618 34620 12624 34672
rect 12676 34660 12682 34672
rect 13648 34660 13676 34700
rect 14108 34700 16120 34728
rect 13998 34660 14004 34672
rect 12676 34632 12834 34660
rect 13648 34632 14004 34660
rect 12676 34620 12682 34632
rect 13998 34620 14004 34632
rect 14056 34620 14062 34672
rect 1765 34595 1823 34601
rect 1765 34561 1777 34595
rect 1811 34561 1823 34595
rect 1765 34555 1823 34561
rect 7282 34552 7288 34604
rect 7340 34592 7346 34604
rect 7929 34595 7987 34601
rect 7929 34592 7941 34595
rect 7340 34564 7941 34592
rect 7340 34552 7346 34564
rect 7929 34561 7941 34564
rect 7975 34561 7987 34595
rect 7929 34555 7987 34561
rect 8021 34595 8079 34601
rect 8021 34561 8033 34595
rect 8067 34592 8079 34595
rect 8067 34564 8616 34592
rect 8067 34561 8079 34564
rect 8021 34555 8079 34561
rect 2038 34484 2044 34536
rect 2096 34484 2102 34536
rect 8036 34524 8064 34555
rect 7300 34496 8064 34524
rect 8113 34527 8171 34533
rect 7300 34468 7328 34496
rect 8113 34493 8125 34527
rect 8159 34493 8171 34527
rect 8588 34524 8616 34564
rect 8662 34552 8668 34604
rect 8720 34592 8726 34604
rect 9125 34595 9183 34601
rect 9125 34592 9137 34595
rect 8720 34564 9137 34592
rect 8720 34552 8726 34564
rect 9125 34561 9137 34564
rect 9171 34561 9183 34595
rect 9950 34592 9956 34604
rect 9125 34555 9183 34561
rect 9232 34564 9956 34592
rect 9232 34524 9260 34564
rect 9950 34552 9956 34564
rect 10008 34552 10014 34604
rect 10321 34595 10379 34601
rect 10321 34561 10333 34595
rect 10367 34592 10379 34595
rect 11882 34592 11888 34604
rect 10367 34564 11888 34592
rect 10367 34561 10379 34564
rect 10321 34555 10379 34561
rect 11882 34552 11888 34564
rect 11940 34552 11946 34604
rect 12066 34552 12072 34604
rect 12124 34552 12130 34604
rect 13630 34552 13636 34604
rect 13688 34592 13694 34604
rect 14108 34592 14136 34700
rect 16114 34688 16120 34700
rect 16172 34728 16178 34740
rect 16301 34731 16359 34737
rect 16301 34728 16313 34731
rect 16172 34700 16313 34728
rect 16172 34688 16178 34700
rect 16301 34697 16313 34700
rect 16347 34697 16359 34731
rect 16301 34691 16359 34697
rect 17494 34688 17500 34740
rect 17552 34728 17558 34740
rect 21453 34731 21511 34737
rect 21453 34728 21465 34731
rect 17552 34700 21465 34728
rect 17552 34688 17558 34700
rect 21453 34697 21465 34700
rect 21499 34728 21511 34731
rect 21818 34728 21824 34740
rect 21499 34700 21824 34728
rect 21499 34697 21511 34700
rect 21453 34691 21511 34697
rect 21818 34688 21824 34700
rect 21876 34688 21882 34740
rect 15378 34620 15384 34672
rect 15436 34620 15442 34672
rect 16206 34620 16212 34672
rect 16264 34660 16270 34672
rect 17218 34660 17224 34672
rect 16264 34632 17224 34660
rect 16264 34620 16270 34632
rect 17218 34620 17224 34632
rect 17276 34620 17282 34672
rect 17402 34620 17408 34672
rect 17460 34660 17466 34672
rect 17681 34663 17739 34669
rect 17681 34660 17693 34663
rect 17460 34632 17693 34660
rect 17460 34620 17466 34632
rect 17681 34629 17693 34632
rect 17727 34629 17739 34663
rect 17681 34623 17739 34629
rect 17954 34620 17960 34672
rect 18012 34660 18018 34672
rect 18012 34632 18170 34660
rect 18012 34620 18018 34632
rect 20714 34620 20720 34672
rect 20772 34620 20778 34672
rect 13688 34564 14136 34592
rect 13688 34552 13694 34564
rect 19702 34552 19708 34604
rect 19760 34552 19766 34604
rect 8588 34496 9260 34524
rect 9309 34527 9367 34533
rect 8113 34487 8171 34493
rect 9309 34493 9321 34527
rect 9355 34493 9367 34527
rect 9309 34487 9367 34493
rect 7282 34416 7288 34468
rect 7340 34416 7346 34468
rect 8128 34456 8156 34487
rect 8202 34456 8208 34468
rect 7484 34428 8208 34456
rect 7098 34348 7104 34400
rect 7156 34388 7162 34400
rect 7484 34388 7512 34428
rect 8202 34416 8208 34428
rect 8260 34416 8266 34468
rect 9324 34456 9352 34487
rect 10226 34484 10232 34536
rect 10284 34524 10290 34536
rect 10502 34524 10508 34536
rect 10284 34496 10508 34524
rect 10284 34484 10290 34496
rect 10502 34484 10508 34496
rect 10560 34484 10566 34536
rect 13538 34484 13544 34536
rect 13596 34524 13602 34536
rect 13817 34527 13875 34533
rect 13817 34524 13829 34527
rect 13596 34496 13829 34524
rect 13596 34484 13602 34496
rect 13817 34493 13829 34496
rect 13863 34493 13875 34527
rect 13817 34487 13875 34493
rect 14274 34484 14280 34536
rect 14332 34524 14338 34536
rect 14553 34527 14611 34533
rect 14553 34524 14565 34527
rect 14332 34496 14565 34524
rect 14332 34484 14338 34496
rect 14553 34493 14565 34496
rect 14599 34493 14611 34527
rect 14553 34487 14611 34493
rect 14826 34484 14832 34536
rect 14884 34484 14890 34536
rect 16666 34484 16672 34536
rect 16724 34524 16730 34536
rect 17405 34527 17463 34533
rect 17405 34524 17417 34527
rect 16724 34496 17417 34524
rect 16724 34484 16730 34496
rect 17405 34493 17417 34496
rect 17451 34493 17463 34527
rect 21542 34524 21548 34536
rect 17405 34487 17463 34493
rect 17512 34496 21548 34524
rect 9398 34456 9404 34468
rect 9324 34428 9404 34456
rect 9398 34416 9404 34428
rect 9456 34416 9462 34468
rect 13998 34416 14004 34468
rect 14056 34456 14062 34468
rect 14366 34456 14372 34468
rect 14056 34428 14372 34456
rect 14056 34416 14062 34428
rect 14366 34416 14372 34428
rect 14424 34416 14430 34468
rect 17310 34416 17316 34468
rect 17368 34456 17374 34468
rect 17512 34456 17540 34496
rect 21542 34484 21548 34496
rect 21600 34484 21606 34536
rect 22554 34456 22560 34468
rect 17368 34428 17540 34456
rect 21008 34428 22560 34456
rect 17368 34416 17374 34428
rect 7156 34360 7512 34388
rect 7156 34348 7162 34360
rect 7558 34348 7564 34400
rect 7616 34348 7622 34400
rect 9950 34348 9956 34400
rect 10008 34348 10014 34400
rect 10042 34348 10048 34400
rect 10100 34388 10106 34400
rect 12066 34388 12072 34400
rect 10100 34360 12072 34388
rect 10100 34348 10106 34360
rect 12066 34348 12072 34360
rect 12124 34348 12130 34400
rect 12158 34348 12164 34400
rect 12216 34388 12222 34400
rect 15194 34388 15200 34400
rect 12216 34360 15200 34388
rect 12216 34348 12222 34360
rect 15194 34348 15200 34360
rect 15252 34348 15258 34400
rect 16482 34348 16488 34400
rect 16540 34388 16546 34400
rect 18782 34388 18788 34400
rect 16540 34360 18788 34388
rect 16540 34348 16546 34360
rect 18782 34348 18788 34360
rect 18840 34388 18846 34400
rect 19153 34391 19211 34397
rect 19153 34388 19165 34391
rect 18840 34360 19165 34388
rect 18840 34348 18846 34360
rect 19153 34357 19165 34360
rect 19199 34357 19211 34391
rect 19153 34351 19211 34357
rect 19968 34391 20026 34397
rect 19968 34357 19980 34391
rect 20014 34388 20026 34391
rect 21008 34388 21036 34428
rect 22554 34416 22560 34428
rect 22612 34416 22618 34468
rect 20014 34360 21036 34388
rect 20014 34357 20026 34360
rect 19968 34351 20026 34357
rect 1104 34298 49864 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 32950 34298
rect 33002 34246 33014 34298
rect 33066 34246 33078 34298
rect 33130 34246 33142 34298
rect 33194 34246 33206 34298
rect 33258 34246 42950 34298
rect 43002 34246 43014 34298
rect 43066 34246 43078 34298
rect 43130 34246 43142 34298
rect 43194 34246 43206 34298
rect 43258 34246 49864 34298
rect 1104 34224 49864 34246
rect 7190 34144 7196 34196
rect 7248 34184 7254 34196
rect 7834 34184 7840 34196
rect 7248 34156 7840 34184
rect 7248 34144 7254 34156
rect 7834 34144 7840 34156
rect 7892 34184 7898 34196
rect 8113 34187 8171 34193
rect 8113 34184 8125 34187
rect 7892 34156 8125 34184
rect 7892 34144 7898 34156
rect 8113 34153 8125 34156
rect 8159 34153 8171 34187
rect 8113 34147 8171 34153
rect 10318 34144 10324 34196
rect 10376 34184 10382 34196
rect 10376 34156 12020 34184
rect 10376 34144 10382 34156
rect 7742 34076 7748 34128
rect 7800 34116 7806 34128
rect 7800 34088 10916 34116
rect 7800 34076 7806 34088
rect 6365 34051 6423 34057
rect 6365 34017 6377 34051
rect 6411 34048 6423 34051
rect 9030 34048 9036 34060
rect 6411 34020 9036 34048
rect 6411 34017 6423 34020
rect 6365 34011 6423 34017
rect 9030 34008 9036 34020
rect 9088 34008 9094 34060
rect 10888 34057 10916 34088
rect 11992 34057 12020 34156
rect 12066 34144 12072 34196
rect 12124 34184 12130 34196
rect 12124 34156 13216 34184
rect 12124 34144 12130 34156
rect 10873 34051 10931 34057
rect 10873 34017 10885 34051
rect 10919 34048 10931 34051
rect 11977 34051 12035 34057
rect 10919 34020 11928 34048
rect 10919 34017 10931 34020
rect 10873 34011 10931 34017
rect 10597 33983 10655 33989
rect 10597 33949 10609 33983
rect 10643 33980 10655 33983
rect 11054 33980 11060 33992
rect 10643 33952 11060 33980
rect 10643 33949 10655 33952
rect 10597 33943 10655 33949
rect 11054 33940 11060 33952
rect 11112 33940 11118 33992
rect 11422 33940 11428 33992
rect 11480 33980 11486 33992
rect 11793 33983 11851 33989
rect 11793 33980 11805 33983
rect 11480 33952 11805 33980
rect 11480 33940 11486 33952
rect 11793 33949 11805 33952
rect 11839 33949 11851 33983
rect 11900 33980 11928 34020
rect 11977 34017 11989 34051
rect 12023 34017 12035 34051
rect 11977 34011 12035 34017
rect 12434 34008 12440 34060
rect 12492 34048 12498 34060
rect 12986 34048 12992 34060
rect 12492 34020 12992 34048
rect 12492 34008 12498 34020
rect 12986 34008 12992 34020
rect 13044 34008 13050 34060
rect 13188 34057 13216 34156
rect 13906 34144 13912 34196
rect 13964 34184 13970 34196
rect 15930 34184 15936 34196
rect 13964 34156 15936 34184
rect 13964 34144 13970 34156
rect 15930 34144 15936 34156
rect 15988 34144 15994 34196
rect 21269 34187 21327 34193
rect 21269 34153 21281 34187
rect 21315 34184 21327 34187
rect 21450 34184 21456 34196
rect 21315 34156 21456 34184
rect 21315 34153 21327 34156
rect 21269 34147 21327 34153
rect 21450 34144 21456 34156
rect 21508 34144 21514 34196
rect 13173 34051 13231 34057
rect 13173 34017 13185 34051
rect 13219 34017 13231 34051
rect 13173 34011 13231 34017
rect 14553 34051 14611 34057
rect 14553 34017 14565 34051
rect 14599 34048 14611 34051
rect 14642 34048 14648 34060
rect 14599 34020 14648 34048
rect 14599 34017 14611 34020
rect 14553 34011 14611 34017
rect 14642 34008 14648 34020
rect 14700 34008 14706 34060
rect 19058 34008 19064 34060
rect 19116 34048 19122 34060
rect 19797 34051 19855 34057
rect 19797 34048 19809 34051
rect 19116 34020 19809 34048
rect 19116 34008 19122 34020
rect 19797 34017 19809 34020
rect 19843 34017 19855 34051
rect 19797 34011 19855 34017
rect 13538 33980 13544 33992
rect 11900 33952 13544 33980
rect 11793 33943 11851 33949
rect 13538 33940 13544 33952
rect 13596 33940 13602 33992
rect 14274 33940 14280 33992
rect 14332 33940 14338 33992
rect 16666 33940 16672 33992
rect 16724 33940 16730 33992
rect 19521 33983 19579 33989
rect 19521 33949 19533 33983
rect 19567 33949 19579 33983
rect 19521 33943 19579 33949
rect 6546 33872 6552 33924
rect 6604 33912 6610 33924
rect 6641 33915 6699 33921
rect 6641 33912 6653 33915
rect 6604 33884 6653 33912
rect 6604 33872 6610 33884
rect 6641 33881 6653 33884
rect 6687 33881 6699 33915
rect 7098 33912 7104 33924
rect 6641 33875 6699 33881
rect 7024 33884 7104 33912
rect 7024 33844 7052 33884
rect 7098 33872 7104 33884
rect 7156 33872 7162 33924
rect 10318 33912 10324 33924
rect 9600 33884 10324 33912
rect 9600 33844 9628 33884
rect 10318 33872 10324 33884
rect 10376 33872 10382 33924
rect 11885 33915 11943 33921
rect 11885 33881 11897 33915
rect 11931 33912 11943 33915
rect 12158 33912 12164 33924
rect 11931 33884 12164 33912
rect 11931 33881 11943 33884
rect 11885 33875 11943 33881
rect 12158 33872 12164 33884
rect 12216 33872 12222 33924
rect 12250 33872 12256 33924
rect 12308 33912 12314 33924
rect 12894 33912 12900 33924
rect 12308 33884 12900 33912
rect 12308 33872 12314 33884
rect 12894 33872 12900 33884
rect 12952 33872 12958 33924
rect 12986 33872 12992 33924
rect 13044 33872 13050 33924
rect 13081 33915 13139 33921
rect 13081 33881 13093 33915
rect 13127 33912 13139 33915
rect 13906 33912 13912 33924
rect 13127 33884 13912 33912
rect 13127 33881 13139 33884
rect 13081 33875 13139 33881
rect 13906 33872 13912 33884
rect 13964 33872 13970 33924
rect 14642 33872 14648 33924
rect 14700 33912 14706 33924
rect 14700 33884 15042 33912
rect 14700 33872 14706 33884
rect 16114 33872 16120 33924
rect 16172 33912 16178 33924
rect 16482 33912 16488 33924
rect 16172 33884 16488 33912
rect 16172 33872 16178 33884
rect 16482 33872 16488 33884
rect 16540 33912 16546 33924
rect 16945 33915 17003 33921
rect 16945 33912 16957 33915
rect 16540 33884 16957 33912
rect 16540 33872 16546 33884
rect 16945 33881 16957 33884
rect 16991 33881 17003 33915
rect 16945 33875 17003 33881
rect 17402 33872 17408 33924
rect 17460 33872 17466 33924
rect 19536 33912 19564 33943
rect 19702 33912 19708 33924
rect 19536 33884 19708 33912
rect 19702 33872 19708 33884
rect 19760 33872 19766 33924
rect 20806 33872 20812 33924
rect 20864 33872 20870 33924
rect 7024 33816 9628 33844
rect 9674 33804 9680 33856
rect 9732 33844 9738 33856
rect 10229 33847 10287 33853
rect 10229 33844 10241 33847
rect 9732 33816 10241 33844
rect 9732 33804 9738 33816
rect 10229 33813 10241 33816
rect 10275 33813 10287 33847
rect 10229 33807 10287 33813
rect 10689 33847 10747 33853
rect 10689 33813 10701 33847
rect 10735 33844 10747 33847
rect 10778 33844 10784 33856
rect 10735 33816 10784 33844
rect 10735 33813 10747 33816
rect 10689 33807 10747 33813
rect 10778 33804 10784 33816
rect 10836 33804 10842 33856
rect 11422 33804 11428 33856
rect 11480 33804 11486 33856
rect 12066 33804 12072 33856
rect 12124 33844 12130 33856
rect 12621 33847 12679 33853
rect 12621 33844 12633 33847
rect 12124 33816 12633 33844
rect 12124 33804 12130 33816
rect 12621 33813 12633 33816
rect 12667 33813 12679 33847
rect 12621 33807 12679 33813
rect 13354 33804 13360 33856
rect 13412 33844 13418 33856
rect 16025 33847 16083 33853
rect 16025 33844 16037 33847
rect 13412 33816 16037 33844
rect 13412 33804 13418 33816
rect 16025 33813 16037 33816
rect 16071 33813 16083 33847
rect 16025 33807 16083 33813
rect 17770 33804 17776 33856
rect 17828 33844 17834 33856
rect 18417 33847 18475 33853
rect 18417 33844 18429 33847
rect 17828 33816 18429 33844
rect 17828 33804 17834 33816
rect 18417 33813 18429 33816
rect 18463 33813 18475 33847
rect 18417 33807 18475 33813
rect 1104 33754 49864 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 27950 33754
rect 28002 33702 28014 33754
rect 28066 33702 28078 33754
rect 28130 33702 28142 33754
rect 28194 33702 28206 33754
rect 28258 33702 37950 33754
rect 38002 33702 38014 33754
rect 38066 33702 38078 33754
rect 38130 33702 38142 33754
rect 38194 33702 38206 33754
rect 38258 33702 47950 33754
rect 48002 33702 48014 33754
rect 48066 33702 48078 33754
rect 48130 33702 48142 33754
rect 48194 33702 48206 33754
rect 48258 33702 49864 33754
rect 1104 33680 49864 33702
rect 7190 33600 7196 33652
rect 7248 33640 7254 33652
rect 7374 33640 7380 33652
rect 7248 33612 7380 33640
rect 7248 33600 7254 33612
rect 7374 33600 7380 33612
rect 7432 33600 7438 33652
rect 7558 33600 7564 33652
rect 7616 33640 7622 33652
rect 8205 33643 8263 33649
rect 8205 33640 8217 33643
rect 7616 33612 8217 33640
rect 7616 33600 7622 33612
rect 8205 33609 8217 33612
rect 8251 33609 8263 33643
rect 8205 33603 8263 33609
rect 8404 33612 10640 33640
rect 6638 33532 6644 33584
rect 6696 33532 6702 33584
rect 6822 33532 6828 33584
rect 6880 33572 6886 33584
rect 8297 33575 8355 33581
rect 8297 33572 8309 33575
rect 6880 33544 8309 33572
rect 6880 33532 6886 33544
rect 8297 33541 8309 33544
rect 8343 33541 8355 33575
rect 8297 33535 8355 33541
rect 1765 33507 1823 33513
rect 1765 33473 1777 33507
rect 1811 33504 1823 33507
rect 6086 33504 6092 33516
rect 1811 33476 6092 33504
rect 1811 33473 1823 33476
rect 1765 33467 1823 33473
rect 6086 33464 6092 33476
rect 6144 33464 6150 33516
rect 1302 33396 1308 33448
rect 1360 33436 1366 33448
rect 2041 33439 2099 33445
rect 2041 33436 2053 33439
rect 1360 33408 2053 33436
rect 1360 33396 1366 33408
rect 2041 33405 2053 33408
rect 2087 33405 2099 33439
rect 2041 33399 2099 33405
rect 7466 33396 7472 33448
rect 7524 33436 7530 33448
rect 8404 33445 8432 33612
rect 10318 33532 10324 33584
rect 10376 33532 10382 33584
rect 9030 33464 9036 33516
rect 9088 33464 9094 33516
rect 10612 33504 10640 33612
rect 12894 33600 12900 33652
rect 12952 33640 12958 33652
rect 15654 33640 15660 33652
rect 12952 33612 15660 33640
rect 12952 33600 12958 33612
rect 15654 33600 15660 33612
rect 15712 33600 15718 33652
rect 16758 33600 16764 33652
rect 16816 33640 16822 33652
rect 17221 33643 17279 33649
rect 17221 33640 17233 33643
rect 16816 33612 17233 33640
rect 16816 33600 16822 33612
rect 17221 33609 17233 33612
rect 17267 33609 17279 33643
rect 17221 33603 17279 33609
rect 17681 33643 17739 33649
rect 17681 33609 17693 33643
rect 17727 33640 17739 33643
rect 18322 33640 18328 33652
rect 17727 33612 18328 33640
rect 17727 33609 17739 33612
rect 17681 33603 17739 33609
rect 18322 33600 18328 33612
rect 18380 33600 18386 33652
rect 18417 33643 18475 33649
rect 18417 33609 18429 33643
rect 18463 33640 18475 33643
rect 18506 33640 18512 33652
rect 18463 33612 18512 33640
rect 18463 33609 18475 33612
rect 18417 33603 18475 33609
rect 18506 33600 18512 33612
rect 18564 33600 18570 33652
rect 18877 33643 18935 33649
rect 18877 33609 18889 33643
rect 18923 33640 18935 33643
rect 21266 33640 21272 33652
rect 18923 33612 21272 33640
rect 18923 33609 18935 33612
rect 18877 33603 18935 33609
rect 21266 33600 21272 33612
rect 21324 33600 21330 33652
rect 10778 33532 10784 33584
rect 10836 33572 10842 33584
rect 13449 33575 13507 33581
rect 13449 33572 13461 33575
rect 10836 33544 13461 33572
rect 10836 33532 10842 33544
rect 13449 33541 13461 33544
rect 13495 33541 13507 33575
rect 13630 33572 13636 33584
rect 13449 33535 13507 33541
rect 13556 33544 13636 33572
rect 11054 33504 11060 33516
rect 10612 33476 11060 33504
rect 11054 33464 11060 33476
rect 11112 33504 11118 33516
rect 12250 33504 12256 33516
rect 11112 33476 12256 33504
rect 11112 33464 11118 33476
rect 12250 33464 12256 33476
rect 12308 33464 12314 33516
rect 13357 33507 13415 33513
rect 13357 33473 13369 33507
rect 13403 33473 13415 33507
rect 13357 33467 13415 33473
rect 8389 33439 8447 33445
rect 8389 33436 8401 33439
rect 7524 33408 8401 33436
rect 7524 33396 7530 33408
rect 8389 33405 8401 33408
rect 8435 33405 8447 33439
rect 9309 33439 9367 33445
rect 9309 33436 9321 33439
rect 8389 33399 8447 33405
rect 8496 33408 9321 33436
rect 8294 33328 8300 33380
rect 8352 33368 8358 33380
rect 8496 33368 8524 33408
rect 9309 33405 9321 33408
rect 9355 33436 9367 33439
rect 10042 33436 10048 33448
rect 9355 33408 10048 33436
rect 9355 33405 9367 33408
rect 9309 33399 9367 33405
rect 10042 33396 10048 33408
rect 10100 33396 10106 33448
rect 8352 33340 8524 33368
rect 13372 33368 13400 33467
rect 13556 33445 13584 33544
rect 13630 33532 13636 33544
rect 13688 33532 13694 33584
rect 14274 33532 14280 33584
rect 14332 33572 14338 33584
rect 16117 33575 16175 33581
rect 16117 33572 16129 33575
rect 14332 33544 16129 33572
rect 14332 33532 14338 33544
rect 16117 33541 16129 33544
rect 16163 33572 16175 33575
rect 16666 33572 16672 33584
rect 16163 33544 16672 33572
rect 16163 33541 16175 33544
rect 16117 33535 16175 33541
rect 16666 33532 16672 33544
rect 16724 33532 16730 33584
rect 13998 33464 14004 33516
rect 14056 33504 14062 33516
rect 14553 33507 14611 33513
rect 14056 33476 14136 33504
rect 14056 33464 14062 33476
rect 13541 33439 13599 33445
rect 13541 33405 13553 33439
rect 13587 33405 13599 33439
rect 13541 33399 13599 33405
rect 13998 33368 14004 33380
rect 13372 33340 14004 33368
rect 8352 33328 8358 33340
rect 13998 33328 14004 33340
rect 14056 33328 14062 33380
rect 14108 33368 14136 33476
rect 14553 33473 14565 33507
rect 14599 33504 14611 33507
rect 14734 33504 14740 33516
rect 14599 33476 14740 33504
rect 14599 33473 14611 33476
rect 14553 33467 14611 33473
rect 14734 33464 14740 33476
rect 14792 33464 14798 33516
rect 15378 33464 15384 33516
rect 15436 33504 15442 33516
rect 16482 33504 16488 33516
rect 15436 33476 16488 33504
rect 15436 33464 15442 33476
rect 16482 33464 16488 33476
rect 16540 33464 16546 33516
rect 17586 33464 17592 33516
rect 17644 33464 17650 33516
rect 18782 33464 18788 33516
rect 18840 33464 18846 33516
rect 19426 33504 19432 33516
rect 18984 33476 19432 33504
rect 14645 33439 14703 33445
rect 14645 33405 14657 33439
rect 14691 33405 14703 33439
rect 14645 33399 14703 33405
rect 14829 33439 14887 33445
rect 14829 33405 14841 33439
rect 14875 33436 14887 33439
rect 15102 33436 15108 33448
rect 14875 33408 15108 33436
rect 14875 33405 14887 33408
rect 14829 33399 14887 33405
rect 14185 33371 14243 33377
rect 14185 33368 14197 33371
rect 14108 33340 14197 33368
rect 14185 33337 14197 33340
rect 14231 33337 14243 33371
rect 14660 33368 14688 33399
rect 15102 33396 15108 33408
rect 15160 33396 15166 33448
rect 17865 33439 17923 33445
rect 17865 33405 17877 33439
rect 17911 33436 17923 33439
rect 18984 33436 19012 33476
rect 19426 33464 19432 33476
rect 19484 33504 19490 33516
rect 20438 33504 20444 33516
rect 19484 33476 20444 33504
rect 19484 33464 19490 33476
rect 20438 33464 20444 33476
rect 20496 33464 20502 33516
rect 17911 33408 19012 33436
rect 17911 33405 17923 33408
rect 17865 33399 17923 33405
rect 19058 33396 19064 33448
rect 19116 33396 19122 33448
rect 18414 33368 18420 33380
rect 14660 33340 18420 33368
rect 14185 33331 14243 33337
rect 18414 33328 18420 33340
rect 18472 33328 18478 33380
rect 5626 33260 5632 33312
rect 5684 33300 5690 33312
rect 6733 33303 6791 33309
rect 6733 33300 6745 33303
rect 5684 33272 6745 33300
rect 5684 33260 5690 33272
rect 6733 33269 6745 33272
rect 6779 33269 6791 33303
rect 6733 33263 6791 33269
rect 7837 33303 7895 33309
rect 7837 33269 7849 33303
rect 7883 33300 7895 33303
rect 10410 33300 10416 33312
rect 7883 33272 10416 33300
rect 7883 33269 7895 33272
rect 7837 33263 7895 33269
rect 10410 33260 10416 33272
rect 10468 33260 10474 33312
rect 12989 33303 13047 33309
rect 12989 33269 13001 33303
rect 13035 33300 13047 33303
rect 17126 33300 17132 33312
rect 13035 33272 17132 33300
rect 13035 33269 13047 33272
rect 12989 33263 13047 33269
rect 17126 33260 17132 33272
rect 17184 33260 17190 33312
rect 1104 33210 49864 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 32950 33210
rect 33002 33158 33014 33210
rect 33066 33158 33078 33210
rect 33130 33158 33142 33210
rect 33194 33158 33206 33210
rect 33258 33158 42950 33210
rect 43002 33158 43014 33210
rect 43066 33158 43078 33210
rect 43130 33158 43142 33210
rect 43194 33158 43206 33210
rect 43258 33158 49864 33210
rect 1104 33136 49864 33158
rect 7558 33056 7564 33108
rect 7616 33096 7622 33108
rect 10505 33099 10563 33105
rect 10505 33096 10517 33099
rect 7616 33068 10517 33096
rect 7616 33056 7622 33068
rect 10505 33065 10517 33068
rect 10551 33065 10563 33099
rect 10505 33059 10563 33065
rect 12342 33056 12348 33108
rect 12400 33096 12406 33108
rect 13449 33099 13507 33105
rect 13449 33096 13461 33099
rect 12400 33068 13461 33096
rect 12400 33056 12406 33068
rect 13449 33065 13461 33068
rect 13495 33065 13507 33099
rect 13449 33059 13507 33065
rect 13998 33056 14004 33108
rect 14056 33096 14062 33108
rect 14553 33099 14611 33105
rect 14553 33096 14565 33099
rect 14056 33068 14565 33096
rect 14056 33056 14062 33068
rect 14553 33065 14565 33068
rect 14599 33065 14611 33099
rect 14553 33059 14611 33065
rect 15013 33099 15071 33105
rect 15013 33065 15025 33099
rect 15059 33096 15071 33099
rect 19150 33096 19156 33108
rect 15059 33068 19156 33096
rect 15059 33065 15071 33068
rect 15013 33059 15071 33065
rect 19150 33056 19156 33068
rect 19208 33056 19214 33108
rect 20809 33099 20867 33105
rect 20809 33065 20821 33099
rect 20855 33096 20867 33099
rect 22002 33096 22008 33108
rect 20855 33068 22008 33096
rect 20855 33065 20867 33068
rect 20809 33059 20867 33065
rect 7469 33031 7527 33037
rect 7469 32997 7481 33031
rect 7515 33028 7527 33031
rect 9766 33028 9772 33040
rect 7515 33000 9772 33028
rect 7515 32997 7527 33000
rect 7469 32991 7527 32997
rect 9766 32988 9772 33000
rect 9824 32988 9830 33040
rect 1302 32920 1308 32972
rect 1360 32960 1366 32972
rect 2041 32963 2099 32969
rect 2041 32960 2053 32963
rect 1360 32932 2053 32960
rect 1360 32920 1366 32932
rect 2041 32929 2053 32932
rect 2087 32929 2099 32963
rect 2041 32923 2099 32929
rect 7742 32920 7748 32972
rect 7800 32960 7806 32972
rect 8021 32963 8079 32969
rect 8021 32960 8033 32963
rect 7800 32932 8033 32960
rect 7800 32920 7806 32932
rect 8021 32929 8033 32932
rect 8067 32929 8079 32963
rect 8021 32923 8079 32929
rect 9953 32963 10011 32969
rect 9953 32929 9965 32963
rect 9999 32960 10011 32963
rect 10870 32960 10876 32972
rect 9999 32932 10876 32960
rect 9999 32929 10011 32932
rect 9953 32923 10011 32929
rect 10870 32920 10876 32932
rect 10928 32920 10934 32972
rect 11057 32963 11115 32969
rect 11057 32960 11069 32963
rect 10980 32932 11069 32960
rect 1765 32895 1823 32901
rect 1765 32861 1777 32895
rect 1811 32892 1823 32895
rect 4706 32892 4712 32904
rect 1811 32864 4712 32892
rect 1811 32861 1823 32864
rect 1765 32855 1823 32861
rect 4706 32852 4712 32864
rect 4764 32852 4770 32904
rect 6914 32852 6920 32904
rect 6972 32892 6978 32904
rect 7837 32895 7895 32901
rect 7837 32892 7849 32895
rect 6972 32864 7849 32892
rect 6972 32852 6978 32864
rect 7837 32861 7849 32864
rect 7883 32861 7895 32895
rect 7837 32855 7895 32861
rect 9214 32852 9220 32904
rect 9272 32892 9278 32904
rect 9677 32895 9735 32901
rect 9677 32892 9689 32895
rect 9272 32864 9689 32892
rect 9272 32852 9278 32864
rect 9677 32861 9689 32864
rect 9723 32861 9735 32895
rect 9677 32855 9735 32861
rect 9769 32895 9827 32901
rect 9769 32861 9781 32895
rect 9815 32892 9827 32895
rect 9858 32892 9864 32904
rect 9815 32864 9864 32892
rect 9815 32861 9827 32864
rect 9769 32855 9827 32861
rect 9858 32852 9864 32864
rect 9916 32852 9922 32904
rect 10594 32852 10600 32904
rect 10652 32892 10658 32904
rect 10980 32892 11008 32932
rect 11057 32929 11069 32932
rect 11103 32929 11115 32963
rect 11057 32923 11115 32929
rect 15657 32963 15715 32969
rect 15657 32929 15669 32963
rect 15703 32960 15715 32963
rect 19242 32960 19248 32972
rect 15703 32932 19248 32960
rect 15703 32929 15715 32932
rect 15657 32923 15715 32929
rect 19242 32920 19248 32932
rect 19300 32920 19306 32972
rect 10652 32864 11008 32892
rect 10652 32852 10658 32864
rect 11698 32852 11704 32904
rect 11756 32852 11762 32904
rect 15381 32895 15439 32901
rect 15381 32861 15393 32895
rect 15427 32892 15439 32895
rect 16393 32895 16451 32901
rect 16393 32892 16405 32895
rect 15427 32864 16405 32892
rect 15427 32861 15439 32864
rect 15381 32855 15439 32861
rect 16393 32861 16405 32864
rect 16439 32861 16451 32895
rect 16393 32855 16451 32861
rect 16482 32852 16488 32904
rect 16540 32892 16546 32904
rect 16945 32895 17003 32901
rect 16945 32892 16957 32895
rect 16540 32864 16957 32892
rect 16540 32852 16546 32864
rect 16945 32861 16957 32864
rect 16991 32892 17003 32895
rect 20824 32892 20852 33059
rect 22002 33056 22008 33068
rect 22060 33056 22066 33108
rect 16991 32864 20852 32892
rect 16991 32861 17003 32864
rect 16945 32855 17003 32861
rect 5442 32784 5448 32836
rect 5500 32784 5506 32836
rect 7650 32784 7656 32836
rect 7708 32824 7714 32836
rect 7929 32827 7987 32833
rect 7929 32824 7941 32827
rect 7708 32796 7941 32824
rect 7708 32784 7714 32796
rect 7929 32793 7941 32796
rect 7975 32793 7987 32827
rect 7929 32787 7987 32793
rect 10686 32784 10692 32836
rect 10744 32824 10750 32836
rect 10873 32827 10931 32833
rect 10873 32824 10885 32827
rect 10744 32796 10885 32824
rect 10744 32784 10750 32796
rect 10873 32793 10885 32796
rect 10919 32793 10931 32827
rect 10873 32787 10931 32793
rect 11974 32784 11980 32836
rect 12032 32784 12038 32836
rect 12710 32784 12716 32836
rect 12768 32784 12774 32836
rect 16850 32824 16856 32836
rect 15396 32796 16856 32824
rect 5534 32716 5540 32768
rect 5592 32716 5598 32768
rect 9306 32716 9312 32768
rect 9364 32716 9370 32768
rect 10962 32716 10968 32768
rect 11020 32756 11026 32768
rect 13814 32756 13820 32768
rect 11020 32728 13820 32756
rect 11020 32716 11026 32728
rect 13814 32716 13820 32728
rect 13872 32716 13878 32768
rect 14918 32716 14924 32768
rect 14976 32756 14982 32768
rect 15396 32756 15424 32796
rect 16850 32784 16856 32796
rect 16908 32784 16914 32836
rect 17773 32827 17831 32833
rect 17773 32793 17785 32827
rect 17819 32824 17831 32827
rect 17862 32824 17868 32836
rect 17819 32796 17868 32824
rect 17819 32793 17831 32796
rect 17773 32787 17831 32793
rect 17862 32784 17868 32796
rect 17920 32784 17926 32836
rect 19518 32784 19524 32836
rect 19576 32784 19582 32836
rect 14976 32728 15424 32756
rect 14976 32716 14982 32728
rect 15470 32716 15476 32768
rect 15528 32716 15534 32768
rect 16022 32716 16028 32768
rect 16080 32756 16086 32768
rect 18966 32756 18972 32768
rect 16080 32728 18972 32756
rect 16080 32716 16086 32728
rect 18966 32716 18972 32728
rect 19024 32716 19030 32768
rect 1104 32666 49864 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 27950 32666
rect 28002 32614 28014 32666
rect 28066 32614 28078 32666
rect 28130 32614 28142 32666
rect 28194 32614 28206 32666
rect 28258 32614 37950 32666
rect 38002 32614 38014 32666
rect 38066 32614 38078 32666
rect 38130 32614 38142 32666
rect 38194 32614 38206 32666
rect 38258 32614 47950 32666
rect 48002 32614 48014 32666
rect 48066 32614 48078 32666
rect 48130 32614 48142 32666
rect 48194 32614 48206 32666
rect 48258 32614 49864 32666
rect 1104 32592 49864 32614
rect 8846 32512 8852 32564
rect 8904 32512 8910 32564
rect 9214 32512 9220 32564
rect 9272 32512 9278 32564
rect 9309 32555 9367 32561
rect 9309 32521 9321 32555
rect 9355 32552 9367 32555
rect 9674 32552 9680 32564
rect 9355 32524 9680 32552
rect 9355 32521 9367 32524
rect 9309 32515 9367 32521
rect 9674 32512 9680 32524
rect 9732 32512 9738 32564
rect 10410 32512 10416 32564
rect 10468 32512 10474 32564
rect 11698 32512 11704 32564
rect 11756 32552 11762 32564
rect 14274 32552 14280 32564
rect 11756 32524 14280 32552
rect 11756 32512 11762 32524
rect 5442 32444 5448 32496
rect 5500 32484 5506 32496
rect 5500 32456 8156 32484
rect 5500 32444 5506 32456
rect 8128 32425 8156 32456
rect 7193 32419 7251 32425
rect 7193 32385 7205 32419
rect 7239 32416 7251 32419
rect 8021 32419 8079 32425
rect 8021 32416 8033 32419
rect 7239 32388 8033 32416
rect 7239 32385 7251 32388
rect 7193 32379 7251 32385
rect 8021 32385 8033 32388
rect 8067 32385 8079 32419
rect 8021 32379 8079 32385
rect 8113 32419 8171 32425
rect 8113 32385 8125 32419
rect 8159 32416 8171 32419
rect 8159 32388 8708 32416
rect 8159 32385 8171 32388
rect 8113 32379 8171 32385
rect 8205 32351 8263 32357
rect 8205 32317 8217 32351
rect 8251 32317 8263 32351
rect 8205 32311 8263 32317
rect 6914 32240 6920 32292
rect 6972 32280 6978 32292
rect 7466 32280 7472 32292
rect 6972 32252 7472 32280
rect 6972 32240 6978 32252
rect 7466 32240 7472 32252
rect 7524 32280 7530 32292
rect 7834 32280 7840 32292
rect 7524 32252 7840 32280
rect 7524 32240 7530 32252
rect 7834 32240 7840 32252
rect 7892 32280 7898 32292
rect 8220 32280 8248 32311
rect 7892 32252 8248 32280
rect 8680 32280 8708 32388
rect 9122 32376 9128 32428
rect 9180 32416 9186 32428
rect 10505 32419 10563 32425
rect 10505 32416 10517 32419
rect 9180 32388 10517 32416
rect 9180 32376 9186 32388
rect 10505 32385 10517 32388
rect 10551 32385 10563 32419
rect 10505 32379 10563 32385
rect 11882 32376 11888 32428
rect 11940 32376 11946 32428
rect 12268 32416 12296 32524
rect 14274 32512 14280 32524
rect 14332 32552 14338 32564
rect 14458 32552 14464 32564
rect 14332 32524 14464 32552
rect 14332 32512 14338 32524
rect 14458 32512 14464 32524
rect 14516 32512 14522 32564
rect 14642 32512 14648 32564
rect 14700 32512 14706 32564
rect 14826 32512 14832 32564
rect 14884 32552 14890 32564
rect 16301 32555 16359 32561
rect 16301 32552 16313 32555
rect 14884 32524 16313 32552
rect 14884 32512 14890 32524
rect 16301 32521 16313 32524
rect 16347 32521 16359 32555
rect 18414 32552 18420 32564
rect 16301 32515 16359 32521
rect 17788 32524 18420 32552
rect 12710 32444 12716 32496
rect 12768 32484 12774 32496
rect 14660 32484 14688 32512
rect 12768 32456 13110 32484
rect 14660 32456 15318 32484
rect 12768 32444 12774 32456
rect 17402 32444 17408 32496
rect 17460 32484 17466 32496
rect 17788 32484 17816 32524
rect 18414 32512 18420 32524
rect 18472 32512 18478 32564
rect 18877 32555 18935 32561
rect 18877 32521 18889 32555
rect 18923 32552 18935 32555
rect 19058 32552 19064 32564
rect 18923 32524 19064 32552
rect 18923 32521 18935 32524
rect 18877 32515 18935 32521
rect 19058 32512 19064 32524
rect 19116 32512 19122 32564
rect 20622 32512 20628 32564
rect 20680 32552 20686 32564
rect 21085 32555 21143 32561
rect 21085 32552 21097 32555
rect 20680 32524 21097 32552
rect 20680 32512 20686 32524
rect 21085 32521 21097 32524
rect 21131 32521 21143 32555
rect 21085 32515 21143 32521
rect 17460 32456 17894 32484
rect 17460 32444 17466 32456
rect 12345 32419 12403 32425
rect 12345 32416 12357 32419
rect 12268 32388 12357 32416
rect 12345 32385 12357 32388
rect 12391 32385 12403 32419
rect 12345 32379 12403 32385
rect 14458 32376 14464 32428
rect 14516 32416 14522 32428
rect 14553 32419 14611 32425
rect 14553 32416 14565 32419
rect 14516 32388 14565 32416
rect 14516 32376 14522 32388
rect 14553 32385 14565 32388
rect 14599 32385 14611 32419
rect 14553 32379 14611 32385
rect 20714 32376 20720 32428
rect 20772 32376 20778 32428
rect 8938 32308 8944 32360
rect 8996 32348 9002 32360
rect 9401 32351 9459 32357
rect 9401 32348 9413 32351
rect 8996 32320 9413 32348
rect 8996 32308 9002 32320
rect 9401 32317 9413 32320
rect 9447 32317 9459 32351
rect 9401 32311 9459 32317
rect 10689 32351 10747 32357
rect 10689 32317 10701 32351
rect 10735 32348 10747 32351
rect 10735 32320 12434 32348
rect 10735 32317 10747 32320
rect 10689 32311 10747 32317
rect 11330 32280 11336 32292
rect 8680 32252 11336 32280
rect 7892 32240 7898 32252
rect 11330 32240 11336 32252
rect 11388 32240 11394 32292
rect 7650 32172 7656 32224
rect 7708 32172 7714 32224
rect 10045 32215 10103 32221
rect 10045 32181 10057 32215
rect 10091 32212 10103 32215
rect 11238 32212 11244 32224
rect 10091 32184 11244 32212
rect 10091 32181 10103 32184
rect 10045 32175 10103 32181
rect 11238 32172 11244 32184
rect 11296 32172 11302 32224
rect 12406 32212 12434 32320
rect 12618 32308 12624 32360
rect 12676 32348 12682 32360
rect 13354 32348 13360 32360
rect 12676 32320 13360 32348
rect 12676 32308 12682 32320
rect 13354 32308 13360 32320
rect 13412 32308 13418 32360
rect 13814 32308 13820 32360
rect 13872 32348 13878 32360
rect 14093 32351 14151 32357
rect 14093 32348 14105 32351
rect 13872 32320 14105 32348
rect 13872 32308 13878 32320
rect 14093 32317 14105 32320
rect 14139 32317 14151 32351
rect 14829 32351 14887 32357
rect 14829 32348 14841 32351
rect 14093 32311 14151 32317
rect 14292 32320 14841 32348
rect 12618 32212 12624 32224
rect 12406 32184 12624 32212
rect 12618 32172 12624 32184
rect 12676 32172 12682 32224
rect 13814 32172 13820 32224
rect 13872 32212 13878 32224
rect 14292 32212 14320 32320
rect 14829 32317 14841 32320
rect 14875 32348 14887 32351
rect 14918 32348 14924 32360
rect 14875 32320 14924 32348
rect 14875 32317 14887 32320
rect 14829 32311 14887 32317
rect 14918 32308 14924 32320
rect 14976 32308 14982 32360
rect 17129 32351 17187 32357
rect 17129 32317 17141 32351
rect 17175 32348 17187 32351
rect 17405 32351 17463 32357
rect 17175 32320 17264 32348
rect 17175 32317 17187 32320
rect 17129 32311 17187 32317
rect 13872 32184 14320 32212
rect 13872 32172 13878 32184
rect 14918 32172 14924 32224
rect 14976 32212 14982 32224
rect 16942 32212 16948 32224
rect 14976 32184 16948 32212
rect 14976 32172 14982 32184
rect 16942 32172 16948 32184
rect 17000 32172 17006 32224
rect 17236 32212 17264 32320
rect 17405 32317 17417 32351
rect 17451 32348 17463 32351
rect 17494 32348 17500 32360
rect 17451 32320 17500 32348
rect 17451 32317 17463 32320
rect 17405 32311 17463 32317
rect 17494 32308 17500 32320
rect 17552 32308 17558 32360
rect 17862 32308 17868 32360
rect 17920 32348 17926 32360
rect 19337 32351 19395 32357
rect 19337 32348 19349 32351
rect 17920 32320 19349 32348
rect 17920 32308 17926 32320
rect 19337 32317 19349 32320
rect 19383 32317 19395 32351
rect 19337 32311 19395 32317
rect 19613 32351 19671 32357
rect 19613 32317 19625 32351
rect 19659 32348 19671 32351
rect 21450 32348 21456 32360
rect 19659 32320 21456 32348
rect 19659 32317 19671 32320
rect 19613 32311 19671 32317
rect 17862 32212 17868 32224
rect 17236 32184 17868 32212
rect 17862 32172 17868 32184
rect 17920 32172 17926 32224
rect 19352 32212 19380 32311
rect 21450 32308 21456 32320
rect 21508 32308 21514 32360
rect 19702 32212 19708 32224
rect 19352 32184 19708 32212
rect 19702 32172 19708 32184
rect 19760 32172 19766 32224
rect 1104 32122 49864 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 32950 32122
rect 33002 32070 33014 32122
rect 33066 32070 33078 32122
rect 33130 32070 33142 32122
rect 33194 32070 33206 32122
rect 33258 32070 42950 32122
rect 43002 32070 43014 32122
rect 43066 32070 43078 32122
rect 43130 32070 43142 32122
rect 43194 32070 43206 32122
rect 43258 32070 49864 32122
rect 1104 32048 49864 32070
rect 6656 31980 9168 32008
rect 1302 31832 1308 31884
rect 1360 31872 1366 31884
rect 6656 31881 6684 31980
rect 2041 31875 2099 31881
rect 2041 31872 2053 31875
rect 1360 31844 2053 31872
rect 1360 31832 1366 31844
rect 2041 31841 2053 31844
rect 2087 31841 2099 31875
rect 2041 31835 2099 31841
rect 6641 31875 6699 31881
rect 6641 31841 6653 31875
rect 6687 31841 6699 31875
rect 6641 31835 6699 31841
rect 6914 31832 6920 31884
rect 6972 31832 6978 31884
rect 9140 31881 9168 31980
rect 10594 31968 10600 32020
rect 10652 32008 10658 32020
rect 10870 32008 10876 32020
rect 10652 31980 10876 32008
rect 10652 31968 10658 31980
rect 10870 31968 10876 31980
rect 10928 31968 10934 32020
rect 12240 32011 12298 32017
rect 12240 31977 12252 32011
rect 12286 32008 12298 32011
rect 13722 32008 13728 32020
rect 12286 31980 13728 32008
rect 12286 31977 12298 31980
rect 12240 31971 12298 31977
rect 13722 31968 13728 31980
rect 13780 31968 13786 32020
rect 14918 31968 14924 32020
rect 14976 31968 14982 32020
rect 16758 32008 16764 32020
rect 16132 31980 16764 32008
rect 11974 31900 11980 31952
rect 12032 31900 12038 31952
rect 9125 31875 9183 31881
rect 9125 31841 9137 31875
rect 9171 31872 9183 31875
rect 10134 31872 10140 31884
rect 9171 31844 10140 31872
rect 9171 31841 9183 31844
rect 9125 31835 9183 31841
rect 10134 31832 10140 31844
rect 10192 31832 10198 31884
rect 11992 31872 12020 31900
rect 12342 31872 12348 31884
rect 11992 31844 12348 31872
rect 12342 31832 12348 31844
rect 12400 31872 12406 31884
rect 13725 31875 13783 31881
rect 13725 31872 13737 31875
rect 12400 31844 13737 31872
rect 12400 31832 12406 31844
rect 13725 31841 13737 31844
rect 13771 31841 13783 31875
rect 13725 31835 13783 31841
rect 15286 31832 15292 31884
rect 15344 31872 15350 31884
rect 15381 31875 15439 31881
rect 15381 31872 15393 31875
rect 15344 31844 15393 31872
rect 15344 31832 15350 31844
rect 15381 31841 15393 31844
rect 15427 31841 15439 31875
rect 15381 31835 15439 31841
rect 15565 31875 15623 31881
rect 15565 31841 15577 31875
rect 15611 31872 15623 31875
rect 16022 31872 16028 31884
rect 15611 31844 16028 31872
rect 15611 31841 15623 31844
rect 15565 31835 15623 31841
rect 16022 31832 16028 31844
rect 16080 31832 16086 31884
rect 16132 31881 16160 31980
rect 16758 31968 16764 31980
rect 16816 31968 16822 32020
rect 17494 31968 17500 32020
rect 17552 32008 17558 32020
rect 17678 32008 17684 32020
rect 17552 31980 17684 32008
rect 17552 31968 17558 31980
rect 17678 31968 17684 31980
rect 17736 32008 17742 32020
rect 17865 32011 17923 32017
rect 17865 32008 17877 32011
rect 17736 31980 17877 32008
rect 17736 31968 17742 31980
rect 17865 31977 17877 31980
rect 17911 31977 17923 32011
rect 17865 31971 17923 31977
rect 16117 31875 16175 31881
rect 16117 31841 16129 31875
rect 16163 31841 16175 31875
rect 16117 31835 16175 31841
rect 16393 31875 16451 31881
rect 16393 31841 16405 31875
rect 16439 31872 16451 31875
rect 17770 31872 17776 31884
rect 16439 31844 17776 31872
rect 16439 31841 16451 31844
rect 16393 31835 16451 31841
rect 17770 31832 17776 31844
rect 17828 31832 17834 31884
rect 1765 31807 1823 31813
rect 1765 31773 1777 31807
rect 1811 31804 1823 31807
rect 5626 31804 5632 31816
rect 1811 31776 5632 31804
rect 1811 31773 1823 31776
rect 1765 31767 1823 31773
rect 5626 31764 5632 31776
rect 5684 31764 5690 31816
rect 11698 31764 11704 31816
rect 11756 31804 11762 31816
rect 11977 31807 12035 31813
rect 11977 31804 11989 31807
rect 11756 31776 11989 31804
rect 11756 31764 11762 31776
rect 11977 31773 11989 31776
rect 12023 31773 12035 31807
rect 11977 31767 12035 31773
rect 14461 31807 14519 31813
rect 14461 31773 14473 31807
rect 14507 31804 14519 31807
rect 14507 31776 15332 31804
rect 14507 31773 14519 31776
rect 14461 31767 14519 31773
rect 9401 31739 9459 31745
rect 7116 31708 7406 31736
rect 7116 31680 7144 31708
rect 9401 31705 9413 31739
rect 9447 31705 9459 31739
rect 9401 31699 9459 31705
rect 7098 31628 7104 31680
rect 7156 31628 7162 31680
rect 7742 31628 7748 31680
rect 7800 31668 7806 31680
rect 8389 31671 8447 31677
rect 8389 31668 8401 31671
rect 7800 31640 8401 31668
rect 7800 31628 7806 31640
rect 8389 31637 8401 31640
rect 8435 31637 8447 31671
rect 9416 31668 9444 31699
rect 10410 31696 10416 31748
rect 10468 31696 10474 31748
rect 12526 31696 12532 31748
rect 12584 31736 12590 31748
rect 12710 31736 12716 31748
rect 12584 31708 12716 31736
rect 12584 31696 12590 31708
rect 12710 31696 12716 31708
rect 12768 31696 12774 31748
rect 15304 31745 15332 31776
rect 15289 31739 15347 31745
rect 15289 31705 15301 31739
rect 15335 31736 15347 31739
rect 15335 31708 15369 31736
rect 15335 31705 15347 31708
rect 15289 31699 15347 31705
rect 15654 31696 15660 31748
rect 15712 31736 15718 31748
rect 15712 31708 16882 31736
rect 15712 31696 15718 31708
rect 10226 31668 10232 31680
rect 9416 31640 10232 31668
rect 8389 31631 8447 31637
rect 10226 31628 10232 31640
rect 10284 31628 10290 31680
rect 1104 31578 49864 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 27950 31578
rect 28002 31526 28014 31578
rect 28066 31526 28078 31578
rect 28130 31526 28142 31578
rect 28194 31526 28206 31578
rect 28258 31526 37950 31578
rect 38002 31526 38014 31578
rect 38066 31526 38078 31578
rect 38130 31526 38142 31578
rect 38194 31526 38206 31578
rect 38258 31526 47950 31578
rect 48002 31526 48014 31578
rect 48066 31526 48078 31578
rect 48130 31526 48142 31578
rect 48194 31526 48206 31578
rect 48258 31526 49864 31578
rect 1104 31504 49864 31526
rect 12710 31424 12716 31476
rect 12768 31464 12774 31476
rect 12768 31436 14228 31464
rect 12768 31424 12774 31436
rect 10410 31356 10416 31408
rect 10468 31356 10474 31408
rect 10686 31356 10692 31408
rect 10744 31396 10750 31408
rect 11149 31399 11207 31405
rect 11149 31396 11161 31399
rect 10744 31368 11161 31396
rect 10744 31356 10750 31368
rect 11149 31365 11161 31368
rect 11195 31365 11207 31399
rect 11149 31359 11207 31365
rect 12526 31356 12532 31408
rect 12584 31356 12590 31408
rect 13538 31356 13544 31408
rect 13596 31396 13602 31408
rect 13725 31399 13783 31405
rect 13725 31396 13737 31399
rect 13596 31368 13737 31396
rect 13596 31356 13602 31368
rect 13725 31365 13737 31368
rect 13771 31365 13783 31399
rect 14200 31396 14228 31436
rect 15102 31424 15108 31476
rect 15160 31464 15166 31476
rect 16301 31467 16359 31473
rect 16301 31464 16313 31467
rect 15160 31436 16313 31464
rect 15160 31424 15166 31436
rect 16301 31433 16313 31436
rect 16347 31433 16359 31467
rect 16301 31427 16359 31433
rect 19426 31424 19432 31476
rect 19484 31424 19490 31476
rect 14918 31396 14924 31408
rect 14200 31368 14924 31396
rect 13725 31359 13783 31365
rect 14918 31356 14924 31368
rect 14976 31396 14982 31408
rect 17862 31396 17868 31408
rect 14976 31368 15318 31396
rect 17696 31368 17868 31396
rect 14976 31356 14982 31368
rect 1765 31331 1823 31337
rect 1765 31297 1777 31331
rect 1811 31328 1823 31331
rect 5534 31328 5540 31340
rect 1811 31300 5540 31328
rect 1811 31297 1823 31300
rect 1765 31291 1823 31297
rect 5534 31288 5540 31300
rect 5592 31288 5598 31340
rect 16758 31288 16764 31340
rect 16816 31328 16822 31340
rect 17696 31337 17724 31368
rect 17862 31356 17868 31368
rect 17920 31356 17926 31408
rect 18414 31356 18420 31408
rect 18472 31356 18478 31408
rect 17681 31331 17739 31337
rect 17681 31328 17693 31331
rect 16816 31300 17693 31328
rect 16816 31288 16822 31300
rect 17681 31297 17693 31300
rect 17727 31297 17739 31331
rect 17681 31291 17739 31297
rect 1302 31220 1308 31272
rect 1360 31260 1366 31272
rect 2041 31263 2099 31269
rect 2041 31260 2053 31263
rect 1360 31232 2053 31260
rect 1360 31220 1366 31232
rect 2041 31229 2053 31232
rect 2087 31229 2099 31263
rect 2041 31223 2099 31229
rect 8386 31220 8392 31272
rect 8444 31260 8450 31272
rect 9125 31263 9183 31269
rect 9125 31260 9137 31263
rect 8444 31232 9137 31260
rect 8444 31220 8450 31232
rect 9125 31229 9137 31232
rect 9171 31229 9183 31263
rect 9125 31223 9183 31229
rect 9401 31263 9459 31269
rect 9401 31229 9413 31263
rect 9447 31260 9459 31263
rect 11330 31260 11336 31272
rect 9447 31232 11336 31260
rect 9447 31229 9459 31232
rect 9401 31223 9459 31229
rect 11330 31220 11336 31232
rect 11388 31220 11394 31272
rect 11698 31220 11704 31272
rect 11756 31220 11762 31272
rect 11977 31263 12035 31269
rect 11977 31229 11989 31263
rect 12023 31260 12035 31263
rect 13538 31260 13544 31272
rect 12023 31232 13544 31260
rect 12023 31229 12035 31232
rect 11977 31223 12035 31229
rect 13538 31220 13544 31232
rect 13596 31220 13602 31272
rect 14550 31220 14556 31272
rect 14608 31220 14614 31272
rect 14826 31220 14832 31272
rect 14884 31260 14890 31272
rect 17494 31260 17500 31272
rect 14884 31232 17500 31260
rect 14884 31220 14890 31232
rect 17494 31220 17500 31232
rect 17552 31220 17558 31272
rect 17957 31263 18015 31269
rect 17957 31229 17969 31263
rect 18003 31260 18015 31263
rect 18322 31260 18328 31272
rect 18003 31232 18328 31260
rect 18003 31229 18015 31232
rect 17957 31223 18015 31229
rect 18322 31220 18328 31232
rect 18380 31260 18386 31272
rect 20622 31260 20628 31272
rect 18380 31232 20628 31260
rect 18380 31220 18386 31232
rect 20622 31220 20628 31232
rect 20680 31220 20686 31272
rect 1104 31034 49864 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 32950 31034
rect 33002 30982 33014 31034
rect 33066 30982 33078 31034
rect 33130 30982 33142 31034
rect 33194 30982 33206 31034
rect 33258 30982 42950 31034
rect 43002 30982 43014 31034
rect 43066 30982 43078 31034
rect 43130 30982 43142 31034
rect 43194 30982 43206 31034
rect 43258 30982 49864 31034
rect 1104 30960 49864 30982
rect 7837 30923 7895 30929
rect 7837 30889 7849 30923
rect 7883 30920 7895 30923
rect 9766 30920 9772 30932
rect 7883 30892 9772 30920
rect 7883 30889 7895 30892
rect 7837 30883 7895 30889
rect 9766 30880 9772 30892
rect 9824 30880 9830 30932
rect 14918 30880 14924 30932
rect 14976 30920 14982 30932
rect 15654 30920 15660 30932
rect 14976 30892 15660 30920
rect 14976 30880 14982 30892
rect 15654 30880 15660 30892
rect 15712 30880 15718 30932
rect 16669 30923 16727 30929
rect 16669 30889 16681 30923
rect 16715 30920 16727 30923
rect 16850 30920 16856 30932
rect 16715 30892 16856 30920
rect 16715 30889 16727 30892
rect 16669 30883 16727 30889
rect 16850 30880 16856 30892
rect 16908 30880 16914 30932
rect 7742 30812 7748 30864
rect 7800 30852 7806 30864
rect 7800 30824 8432 30852
rect 7800 30812 7806 30824
rect 7834 30744 7840 30796
rect 7892 30784 7898 30796
rect 8404 30793 8432 30824
rect 8297 30787 8355 30793
rect 8297 30784 8309 30787
rect 7892 30756 8309 30784
rect 7892 30744 7898 30756
rect 8297 30753 8309 30756
rect 8343 30753 8355 30787
rect 8297 30747 8355 30753
rect 8389 30787 8447 30793
rect 8389 30753 8401 30787
rect 8435 30753 8447 30787
rect 8389 30747 8447 30753
rect 10134 30744 10140 30796
rect 10192 30784 10198 30796
rect 10229 30787 10287 30793
rect 10229 30784 10241 30787
rect 10192 30756 10241 30784
rect 10192 30744 10198 30756
rect 10229 30753 10241 30756
rect 10275 30784 10287 30787
rect 10873 30787 10931 30793
rect 10873 30784 10885 30787
rect 10275 30756 10885 30784
rect 10275 30753 10287 30756
rect 10229 30747 10287 30753
rect 10873 30753 10885 30756
rect 10919 30784 10931 30787
rect 11698 30784 11704 30796
rect 10919 30756 11704 30784
rect 10919 30753 10931 30756
rect 10873 30747 10931 30753
rect 11698 30744 11704 30756
rect 11756 30744 11762 30796
rect 14550 30744 14556 30796
rect 14608 30784 14614 30796
rect 14921 30787 14979 30793
rect 14921 30784 14933 30787
rect 14608 30756 14933 30784
rect 14608 30744 14614 30756
rect 14921 30753 14933 30756
rect 14967 30784 14979 30787
rect 16758 30784 16764 30796
rect 14967 30756 16764 30784
rect 14967 30753 14979 30756
rect 14921 30747 14979 30753
rect 16758 30744 16764 30756
rect 16816 30744 16822 30796
rect 7650 30676 7656 30728
rect 7708 30716 7714 30728
rect 8205 30719 8263 30725
rect 8205 30716 8217 30719
rect 7708 30688 8217 30716
rect 7708 30676 7714 30688
rect 8205 30685 8217 30688
rect 8251 30685 8263 30719
rect 8205 30679 8263 30685
rect 9490 30676 9496 30728
rect 9548 30676 9554 30728
rect 14458 30676 14464 30728
rect 14516 30676 14522 30728
rect 9508 30580 9536 30676
rect 11054 30608 11060 30660
rect 11112 30648 11118 30660
rect 11149 30651 11207 30657
rect 11149 30648 11161 30651
rect 11112 30620 11161 30648
rect 11112 30608 11118 30620
rect 11149 30617 11161 30620
rect 11195 30617 11207 30651
rect 11149 30611 11207 30617
rect 11606 30608 11612 30660
rect 11664 30608 11670 30660
rect 12544 30620 12756 30648
rect 11882 30580 11888 30592
rect 9508 30552 11888 30580
rect 11882 30540 11888 30552
rect 11940 30580 11946 30592
rect 12544 30580 12572 30620
rect 11940 30552 12572 30580
rect 11940 30540 11946 30552
rect 12618 30540 12624 30592
rect 12676 30540 12682 30592
rect 12728 30580 12756 30620
rect 15102 30608 15108 30660
rect 15160 30648 15166 30660
rect 15197 30651 15255 30657
rect 15197 30648 15209 30651
rect 15160 30620 15209 30648
rect 15160 30608 15166 30620
rect 15197 30617 15209 30620
rect 15243 30617 15255 30651
rect 15197 30611 15255 30617
rect 15654 30608 15660 30660
rect 15712 30608 15718 30660
rect 15378 30580 15384 30592
rect 12728 30552 15384 30580
rect 15378 30540 15384 30552
rect 15436 30540 15442 30592
rect 1104 30490 49864 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 27950 30490
rect 28002 30438 28014 30490
rect 28066 30438 28078 30490
rect 28130 30438 28142 30490
rect 28194 30438 28206 30490
rect 28258 30438 37950 30490
rect 38002 30438 38014 30490
rect 38066 30438 38078 30490
rect 38130 30438 38142 30490
rect 38194 30438 38206 30490
rect 38258 30438 47950 30490
rect 48002 30438 48014 30490
rect 48066 30438 48078 30490
rect 48130 30438 48142 30490
rect 48194 30438 48206 30490
rect 48258 30438 49864 30490
rect 1104 30416 49864 30438
rect 10410 30376 10416 30388
rect 9646 30348 10416 30376
rect 9646 30308 9674 30348
rect 10410 30336 10416 30348
rect 10468 30336 10474 30388
rect 11054 30336 11060 30388
rect 11112 30376 11118 30388
rect 11698 30376 11704 30388
rect 11112 30348 11704 30376
rect 11112 30336 11118 30348
rect 11698 30336 11704 30348
rect 11756 30336 11762 30388
rect 9522 30280 9674 30308
rect 10042 30268 10048 30320
rect 10100 30268 10106 30320
rect 10428 30308 10456 30336
rect 11606 30308 11612 30320
rect 10428 30280 11612 30308
rect 11606 30268 11612 30280
rect 11664 30308 11670 30320
rect 12526 30308 12532 30320
rect 11664 30280 12532 30308
rect 11664 30268 11670 30280
rect 12526 30268 12532 30280
rect 12584 30268 12590 30320
rect 1762 30200 1768 30252
rect 1820 30200 1826 30252
rect 9582 30200 9588 30252
rect 9640 30240 9646 30252
rect 11790 30240 11796 30252
rect 9640 30212 11796 30240
rect 9640 30200 9646 30212
rect 11790 30200 11796 30212
rect 11848 30200 11854 30252
rect 14369 30243 14427 30249
rect 14369 30209 14381 30243
rect 14415 30240 14427 30243
rect 15381 30243 15439 30249
rect 15381 30240 15393 30243
rect 14415 30212 15393 30240
rect 14415 30209 14427 30212
rect 14369 30203 14427 30209
rect 15381 30209 15393 30212
rect 15427 30209 15439 30243
rect 15381 30203 15439 30209
rect 1302 30132 1308 30184
rect 1360 30172 1366 30184
rect 2041 30175 2099 30181
rect 2041 30172 2053 30175
rect 1360 30144 2053 30172
rect 1360 30132 1366 30144
rect 2041 30141 2053 30144
rect 2087 30141 2099 30175
rect 2041 30135 2099 30141
rect 8021 30175 8079 30181
rect 8021 30141 8033 30175
rect 8067 30141 8079 30175
rect 8021 30135 8079 30141
rect 8297 30175 8355 30181
rect 8297 30141 8309 30175
rect 8343 30172 8355 30175
rect 9674 30172 9680 30184
rect 8343 30144 9680 30172
rect 8343 30141 8355 30144
rect 8297 30135 8355 30141
rect 8036 30036 8064 30135
rect 9674 30132 9680 30144
rect 9732 30132 9738 30184
rect 12069 30175 12127 30181
rect 12069 30141 12081 30175
rect 12115 30172 12127 30175
rect 12618 30172 12624 30184
rect 12115 30144 12624 30172
rect 12115 30141 12127 30144
rect 12069 30135 12127 30141
rect 12618 30132 12624 30144
rect 12676 30132 12682 30184
rect 13538 30132 13544 30184
rect 13596 30132 13602 30184
rect 13814 30132 13820 30184
rect 13872 30172 13878 30184
rect 14461 30175 14519 30181
rect 14461 30172 14473 30175
rect 13872 30144 14473 30172
rect 13872 30132 13878 30144
rect 14461 30141 14473 30144
rect 14507 30141 14519 30175
rect 14461 30135 14519 30141
rect 14645 30175 14703 30181
rect 14645 30141 14657 30175
rect 14691 30172 14703 30175
rect 17310 30172 17316 30184
rect 14691 30144 17316 30172
rect 14691 30141 14703 30144
rect 14645 30135 14703 30141
rect 17310 30132 17316 30144
rect 17368 30132 17374 30184
rect 14001 30107 14059 30113
rect 14001 30073 14013 30107
rect 14047 30104 14059 30107
rect 14090 30104 14096 30116
rect 14047 30076 14096 30104
rect 14047 30073 14059 30076
rect 14001 30067 14059 30073
rect 14090 30064 14096 30076
rect 14148 30064 14154 30116
rect 8386 30036 8392 30048
rect 8036 30008 8392 30036
rect 8386 29996 8392 30008
rect 8444 29996 8450 30048
rect 9030 29996 9036 30048
rect 9088 30036 9094 30048
rect 14642 30036 14648 30048
rect 9088 30008 14648 30036
rect 9088 29996 9094 30008
rect 14642 29996 14648 30008
rect 14700 29996 14706 30048
rect 1104 29946 49864 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 32950 29946
rect 33002 29894 33014 29946
rect 33066 29894 33078 29946
rect 33130 29894 33142 29946
rect 33194 29894 33206 29946
rect 33258 29894 42950 29946
rect 43002 29894 43014 29946
rect 43066 29894 43078 29946
rect 43130 29894 43142 29946
rect 43194 29894 43206 29946
rect 43258 29894 49864 29946
rect 1104 29872 49864 29894
rect 1762 29792 1768 29844
rect 1820 29832 1826 29844
rect 9030 29832 9036 29844
rect 1820 29804 9036 29832
rect 1820 29792 1826 29804
rect 9030 29792 9036 29804
rect 9088 29792 9094 29844
rect 11146 29832 11152 29844
rect 9232 29804 11152 29832
rect 9232 29696 9260 29804
rect 11146 29792 11152 29804
rect 11204 29792 11210 29844
rect 11330 29792 11336 29844
rect 11388 29832 11394 29844
rect 11425 29835 11483 29841
rect 11425 29832 11437 29835
rect 11388 29804 11437 29832
rect 11388 29792 11394 29804
rect 11425 29801 11437 29804
rect 11471 29801 11483 29835
rect 11425 29795 11483 29801
rect 14277 29835 14335 29841
rect 14277 29801 14289 29835
rect 14323 29832 14335 29835
rect 14366 29832 14372 29844
rect 14323 29804 14372 29832
rect 14323 29801 14335 29804
rect 14277 29795 14335 29801
rect 14366 29792 14372 29804
rect 14424 29792 14430 29844
rect 1780 29668 9260 29696
rect 9677 29699 9735 29705
rect 1780 29637 1808 29668
rect 9677 29665 9689 29699
rect 9723 29696 9735 29699
rect 10042 29696 10048 29708
rect 9723 29668 10048 29696
rect 9723 29665 9735 29668
rect 9677 29659 9735 29665
rect 10042 29656 10048 29668
rect 10100 29656 10106 29708
rect 11790 29656 11796 29708
rect 11848 29696 11854 29708
rect 12621 29699 12679 29705
rect 12621 29696 12633 29699
rect 11848 29668 12633 29696
rect 11848 29656 11854 29668
rect 12621 29665 12633 29668
rect 12667 29665 12679 29699
rect 12621 29659 12679 29665
rect 13262 29656 13268 29708
rect 13320 29696 13326 29708
rect 13722 29696 13728 29708
rect 13320 29668 13728 29696
rect 13320 29656 13326 29668
rect 13722 29656 13728 29668
rect 13780 29656 13786 29708
rect 14921 29699 14979 29705
rect 14921 29665 14933 29699
rect 14967 29696 14979 29699
rect 16114 29696 16120 29708
rect 14967 29668 16120 29696
rect 14967 29665 14979 29668
rect 14921 29659 14979 29665
rect 16114 29656 16120 29668
rect 16172 29656 16178 29708
rect 1765 29631 1823 29637
rect 1765 29597 1777 29631
rect 1811 29597 1823 29631
rect 1765 29591 1823 29597
rect 11882 29588 11888 29640
rect 11940 29588 11946 29640
rect 14458 29588 14464 29640
rect 14516 29628 14522 29640
rect 14645 29631 14703 29637
rect 14645 29628 14657 29631
rect 14516 29600 14657 29628
rect 14516 29588 14522 29600
rect 14645 29597 14657 29600
rect 14691 29597 14703 29631
rect 14645 29591 14703 29597
rect 14734 29588 14740 29640
rect 14792 29588 14798 29640
rect 1302 29520 1308 29572
rect 1360 29560 1366 29572
rect 2501 29563 2559 29569
rect 2501 29560 2513 29563
rect 1360 29532 2513 29560
rect 1360 29520 1366 29532
rect 2501 29529 2513 29532
rect 2547 29529 2559 29563
rect 2501 29523 2559 29529
rect 9953 29563 10011 29569
rect 9953 29529 9965 29563
rect 9999 29529 10011 29563
rect 9953 29523 10011 29529
rect 9968 29492 9996 29523
rect 10042 29520 10048 29572
rect 10100 29560 10106 29572
rect 10410 29560 10416 29572
rect 10100 29532 10416 29560
rect 10100 29520 10106 29532
rect 10410 29520 10416 29532
rect 10468 29520 10474 29572
rect 13722 29520 13728 29572
rect 13780 29560 13786 29572
rect 14752 29560 14780 29588
rect 13780 29532 14780 29560
rect 13780 29520 13786 29532
rect 10594 29492 10600 29504
rect 9968 29464 10600 29492
rect 10594 29452 10600 29464
rect 10652 29452 10658 29504
rect 14734 29452 14740 29504
rect 14792 29452 14798 29504
rect 1104 29402 49864 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 27950 29402
rect 28002 29350 28014 29402
rect 28066 29350 28078 29402
rect 28130 29350 28142 29402
rect 28194 29350 28206 29402
rect 28258 29350 37950 29402
rect 38002 29350 38014 29402
rect 38066 29350 38078 29402
rect 38130 29350 38142 29402
rect 38194 29350 38206 29402
rect 38258 29350 47950 29402
rect 48002 29350 48014 29402
rect 48066 29350 48078 29402
rect 48130 29350 48142 29402
rect 48194 29350 48206 29402
rect 48258 29350 49864 29402
rect 1104 29328 49864 29350
rect 8386 29288 8392 29300
rect 7484 29260 8392 29288
rect 7484 29161 7512 29260
rect 8386 29248 8392 29260
rect 8444 29288 8450 29300
rect 9582 29288 9588 29300
rect 8444 29260 9588 29288
rect 8444 29248 8450 29260
rect 9582 29248 9588 29260
rect 9640 29248 9646 29300
rect 9950 29248 9956 29300
rect 10008 29288 10014 29300
rect 10597 29291 10655 29297
rect 10597 29288 10609 29291
rect 10008 29260 10609 29288
rect 10008 29248 10014 29260
rect 10597 29257 10609 29260
rect 10643 29257 10655 29291
rect 10597 29251 10655 29257
rect 13265 29291 13323 29297
rect 13265 29257 13277 29291
rect 13311 29288 13323 29291
rect 15010 29288 15016 29300
rect 13311 29260 15016 29288
rect 13311 29257 13323 29260
rect 13265 29251 13323 29257
rect 15010 29248 15016 29260
rect 15068 29248 15074 29300
rect 7742 29180 7748 29232
rect 7800 29180 7806 29232
rect 10042 29220 10048 29232
rect 8970 29192 10048 29220
rect 10042 29180 10048 29192
rect 10100 29180 10106 29232
rect 12618 29180 12624 29232
rect 12676 29220 12682 29232
rect 12676 29192 13492 29220
rect 12676 29180 12682 29192
rect 7469 29155 7527 29161
rect 7469 29121 7481 29155
rect 7515 29121 7527 29155
rect 7469 29115 7527 29121
rect 10594 29112 10600 29164
rect 10652 29152 10658 29164
rect 10652 29124 10824 29152
rect 10652 29112 10658 29124
rect 9217 29087 9275 29093
rect 9217 29053 9229 29087
rect 9263 29084 9275 29087
rect 9674 29084 9680 29096
rect 9263 29056 9680 29084
rect 9263 29053 9275 29056
rect 9217 29047 9275 29053
rect 9674 29044 9680 29056
rect 9732 29044 9738 29096
rect 10686 29044 10692 29096
rect 10744 29044 10750 29096
rect 10796 29093 10824 29124
rect 10781 29087 10839 29093
rect 10781 29053 10793 29087
rect 10827 29053 10839 29087
rect 10781 29047 10839 29053
rect 12526 29044 12532 29096
rect 12584 29084 12590 29096
rect 12802 29084 12808 29096
rect 12584 29056 12808 29084
rect 12584 29044 12590 29056
rect 12802 29044 12808 29056
rect 12860 29044 12866 29096
rect 13354 29044 13360 29096
rect 13412 29044 13418 29096
rect 13464 29093 13492 29192
rect 13449 29087 13507 29093
rect 13449 29053 13461 29087
rect 13495 29053 13507 29087
rect 13449 29047 13507 29053
rect 10229 29019 10287 29025
rect 10229 28985 10241 29019
rect 10275 29016 10287 29019
rect 12066 29016 12072 29028
rect 10275 28988 12072 29016
rect 10275 28985 10287 28988
rect 10229 28979 10287 28985
rect 12066 28976 12072 28988
rect 12124 28976 12130 29028
rect 12728 28994 13032 29016
rect 12636 28988 13032 28994
rect 12636 28966 12756 28988
rect 8202 28908 8208 28960
rect 8260 28948 8266 28960
rect 12636 28948 12664 28966
rect 8260 28920 12664 28948
rect 8260 28908 8266 28920
rect 12802 28908 12808 28960
rect 12860 28948 12866 28960
rect 12897 28951 12955 28957
rect 12897 28948 12909 28951
rect 12860 28920 12909 28948
rect 12860 28908 12866 28920
rect 12897 28917 12909 28920
rect 12943 28917 12955 28951
rect 13004 28948 13032 28988
rect 13998 28948 14004 28960
rect 13004 28920 14004 28948
rect 12897 28911 12955 28917
rect 13998 28908 14004 28920
rect 14056 28908 14062 28960
rect 1104 28858 49864 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 32950 28858
rect 33002 28806 33014 28858
rect 33066 28806 33078 28858
rect 33130 28806 33142 28858
rect 33194 28806 33206 28858
rect 33258 28806 42950 28858
rect 43002 28806 43014 28858
rect 43066 28806 43078 28858
rect 43130 28806 43142 28858
rect 43194 28806 43206 28858
rect 43258 28806 49864 28858
rect 1104 28784 49864 28806
rect 7834 28704 7840 28756
rect 7892 28704 7898 28756
rect 9861 28747 9919 28753
rect 9861 28713 9873 28747
rect 9907 28744 9919 28747
rect 10686 28744 10692 28756
rect 9907 28716 10692 28744
rect 9907 28713 9919 28716
rect 9861 28707 9919 28713
rect 10686 28704 10692 28716
rect 10744 28704 10750 28756
rect 11149 28747 11207 28753
rect 11149 28713 11161 28747
rect 11195 28744 11207 28747
rect 13354 28744 13360 28756
rect 11195 28716 13360 28744
rect 11195 28713 11207 28716
rect 11149 28707 11207 28713
rect 13354 28704 13360 28716
rect 13412 28704 13418 28756
rect 13538 28704 13544 28756
rect 13596 28704 13602 28756
rect 7466 28636 7472 28688
rect 7524 28676 7530 28688
rect 7524 28648 8432 28676
rect 7524 28636 7530 28648
rect 1302 28568 1308 28620
rect 1360 28608 1366 28620
rect 2041 28611 2099 28617
rect 2041 28608 2053 28611
rect 1360 28580 2053 28608
rect 1360 28568 1366 28580
rect 2041 28577 2053 28580
rect 2087 28577 2099 28611
rect 2041 28571 2099 28577
rect 7558 28568 7564 28620
rect 7616 28608 7622 28620
rect 8404 28617 8432 28648
rect 11606 28636 11612 28688
rect 11664 28676 11670 28688
rect 12345 28679 12403 28685
rect 11664 28648 12112 28676
rect 11664 28636 11670 28648
rect 8297 28611 8355 28617
rect 8297 28608 8309 28611
rect 7616 28580 8309 28608
rect 7616 28568 7622 28580
rect 8297 28577 8309 28580
rect 8343 28577 8355 28611
rect 8297 28571 8355 28577
rect 8389 28611 8447 28617
rect 8389 28577 8401 28611
rect 8435 28577 8447 28611
rect 8389 28571 8447 28577
rect 10226 28568 10232 28620
rect 10284 28608 10290 28620
rect 10413 28611 10471 28617
rect 10413 28608 10425 28611
rect 10284 28580 10425 28608
rect 10284 28568 10290 28580
rect 10413 28577 10425 28580
rect 10459 28577 10471 28611
rect 11624 28608 11652 28636
rect 10413 28571 10471 28577
rect 11532 28580 11652 28608
rect 1762 28500 1768 28552
rect 1820 28500 1826 28552
rect 7742 28500 7748 28552
rect 7800 28540 7806 28552
rect 8202 28540 8208 28552
rect 7800 28512 8208 28540
rect 7800 28500 7806 28512
rect 8202 28500 8208 28512
rect 8260 28500 8266 28552
rect 10321 28543 10379 28549
rect 10321 28509 10333 28543
rect 10367 28540 10379 28543
rect 11422 28540 11428 28552
rect 10367 28512 11428 28540
rect 10367 28509 10379 28512
rect 10321 28503 10379 28509
rect 11422 28500 11428 28512
rect 11480 28500 11486 28552
rect 11532 28549 11560 28580
rect 11698 28568 11704 28620
rect 11756 28568 11762 28620
rect 11517 28543 11575 28549
rect 11517 28509 11529 28543
rect 11563 28509 11575 28543
rect 11517 28503 11575 28509
rect 11609 28543 11667 28549
rect 11609 28509 11621 28543
rect 11655 28540 11667 28543
rect 11974 28540 11980 28552
rect 11655 28512 11980 28540
rect 11655 28509 11667 28512
rect 11609 28503 11667 28509
rect 11974 28500 11980 28512
rect 12032 28500 12038 28552
rect 12084 28540 12112 28648
rect 12345 28645 12357 28679
rect 12391 28676 12403 28679
rect 13556 28676 13584 28704
rect 12391 28648 13584 28676
rect 12391 28645 12403 28648
rect 12345 28639 12403 28645
rect 12434 28568 12440 28620
rect 12492 28608 12498 28620
rect 12897 28611 12955 28617
rect 12897 28608 12909 28611
rect 12492 28580 12909 28608
rect 12492 28568 12498 28580
rect 12897 28577 12909 28580
rect 12943 28577 12955 28611
rect 12897 28571 12955 28577
rect 15286 28540 15292 28552
rect 12084 28512 15292 28540
rect 15286 28500 15292 28512
rect 15344 28500 15350 28552
rect 10226 28432 10232 28484
rect 10284 28472 10290 28484
rect 14734 28472 14740 28484
rect 10284 28444 14740 28472
rect 10284 28432 10290 28444
rect 14734 28432 14740 28444
rect 14792 28432 14798 28484
rect 12710 28364 12716 28416
rect 12768 28364 12774 28416
rect 12805 28407 12863 28413
rect 12805 28373 12817 28407
rect 12851 28404 12863 28407
rect 19886 28404 19892 28416
rect 12851 28376 19892 28404
rect 12851 28373 12863 28376
rect 12805 28367 12863 28373
rect 19886 28364 19892 28376
rect 19944 28364 19950 28416
rect 1104 28314 49864 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 27950 28314
rect 28002 28262 28014 28314
rect 28066 28262 28078 28314
rect 28130 28262 28142 28314
rect 28194 28262 28206 28314
rect 28258 28262 37950 28314
rect 38002 28262 38014 28314
rect 38066 28262 38078 28314
rect 38130 28262 38142 28314
rect 38194 28262 38206 28314
rect 38258 28262 47950 28314
rect 48002 28262 48014 28314
rect 48066 28262 48078 28314
rect 48130 28262 48142 28314
rect 48194 28262 48206 28314
rect 48258 28262 49864 28314
rect 1104 28240 49864 28262
rect 9766 28160 9772 28212
rect 9824 28160 9830 28212
rect 9858 28160 9864 28212
rect 9916 28160 9922 28212
rect 12802 28160 12808 28212
rect 12860 28200 12866 28212
rect 12989 28203 13047 28209
rect 12989 28200 13001 28203
rect 12860 28172 13001 28200
rect 12860 28160 12866 28172
rect 12989 28169 13001 28172
rect 13035 28169 13047 28203
rect 12989 28163 13047 28169
rect 6886 28104 12434 28132
rect 1765 28067 1823 28073
rect 1765 28033 1777 28067
rect 1811 28064 1823 28067
rect 6886 28064 6914 28104
rect 1811 28036 6914 28064
rect 12406 28064 12434 28104
rect 12618 28092 12624 28144
rect 12676 28132 12682 28144
rect 13081 28135 13139 28141
rect 13081 28132 13093 28135
rect 12676 28104 13093 28132
rect 12676 28092 12682 28104
rect 13081 28101 13093 28104
rect 13127 28101 13139 28135
rect 13081 28095 13139 28101
rect 20990 28064 20996 28076
rect 12406 28036 20996 28064
rect 1811 28033 1823 28036
rect 1765 28027 1823 28033
rect 20990 28024 20996 28036
rect 21048 28024 21054 28076
rect 1302 27956 1308 28008
rect 1360 27996 1366 28008
rect 2041 27999 2099 28005
rect 2041 27996 2053 27999
rect 1360 27968 2053 27996
rect 1360 27956 1366 27968
rect 2041 27965 2053 27968
rect 2087 27965 2099 27999
rect 2041 27959 2099 27965
rect 9953 27999 10011 28005
rect 9953 27965 9965 27999
rect 9999 27965 10011 27999
rect 9953 27959 10011 27965
rect 13265 27999 13323 28005
rect 13265 27965 13277 27999
rect 13311 27996 13323 27999
rect 13630 27996 13636 28008
rect 13311 27968 13636 27996
rect 13311 27965 13323 27968
rect 13265 27959 13323 27965
rect 9674 27888 9680 27940
rect 9732 27928 9738 27940
rect 9968 27928 9996 27959
rect 13630 27956 13636 27968
rect 13688 27956 13694 28008
rect 9732 27900 9996 27928
rect 9732 27888 9738 27900
rect 9398 27820 9404 27872
rect 9456 27820 9462 27872
rect 12621 27863 12679 27869
rect 12621 27829 12633 27863
rect 12667 27860 12679 27863
rect 15102 27860 15108 27872
rect 12667 27832 15108 27860
rect 12667 27829 12679 27832
rect 12621 27823 12679 27829
rect 15102 27820 15108 27832
rect 15160 27820 15166 27872
rect 1104 27770 49864 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 32950 27770
rect 33002 27718 33014 27770
rect 33066 27718 33078 27770
rect 33130 27718 33142 27770
rect 33194 27718 33206 27770
rect 33258 27718 42950 27770
rect 43002 27718 43014 27770
rect 43066 27718 43078 27770
rect 43130 27718 43142 27770
rect 43194 27718 43206 27770
rect 43258 27718 49864 27770
rect 1104 27696 49864 27718
rect 11514 27548 11520 27600
rect 11572 27588 11578 27600
rect 11701 27591 11759 27597
rect 11701 27588 11713 27591
rect 11572 27560 11713 27588
rect 11572 27548 11578 27560
rect 11701 27557 11713 27560
rect 11747 27557 11759 27591
rect 11701 27551 11759 27557
rect 12342 27480 12348 27532
rect 12400 27480 12406 27532
rect 13173 27455 13231 27461
rect 13173 27421 13185 27455
rect 13219 27452 13231 27455
rect 14182 27452 14188 27464
rect 13219 27424 14188 27452
rect 13219 27421 13231 27424
rect 13173 27415 13231 27421
rect 14182 27412 14188 27424
rect 14240 27412 14246 27464
rect 12069 27387 12127 27393
rect 12069 27384 12081 27387
rect 6886 27356 12081 27384
rect 1670 27276 1676 27328
rect 1728 27316 1734 27328
rect 6886 27316 6914 27356
rect 12069 27353 12081 27356
rect 12115 27353 12127 27387
rect 12069 27347 12127 27353
rect 12161 27387 12219 27393
rect 12161 27353 12173 27387
rect 12207 27384 12219 27387
rect 18690 27384 18696 27396
rect 12207 27356 18696 27384
rect 12207 27353 12219 27356
rect 12161 27347 12219 27353
rect 18690 27344 18696 27356
rect 18748 27344 18754 27396
rect 1728 27288 6914 27316
rect 12989 27319 13047 27325
rect 1728 27276 1734 27288
rect 12989 27285 13001 27319
rect 13035 27316 13047 27319
rect 17126 27316 17132 27328
rect 13035 27288 17132 27316
rect 13035 27285 13047 27288
rect 12989 27279 13047 27285
rect 17126 27276 17132 27288
rect 17184 27276 17190 27328
rect 1104 27226 49864 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 27950 27226
rect 28002 27174 28014 27226
rect 28066 27174 28078 27226
rect 28130 27174 28142 27226
rect 28194 27174 28206 27226
rect 28258 27174 37950 27226
rect 38002 27174 38014 27226
rect 38066 27174 38078 27226
rect 38130 27174 38142 27226
rect 38194 27174 38206 27226
rect 38258 27174 47950 27226
rect 48002 27174 48014 27226
rect 48066 27174 48078 27226
rect 48130 27174 48142 27226
rect 48194 27174 48206 27226
rect 48258 27174 49864 27226
rect 1104 27152 49864 27174
rect 12066 27072 12072 27124
rect 12124 27072 12130 27124
rect 1857 27047 1915 27053
rect 1857 27013 1869 27047
rect 1903 27044 1915 27047
rect 6454 27044 6460 27056
rect 1903 27016 6460 27044
rect 1903 27013 1915 27016
rect 1857 27007 1915 27013
rect 6454 27004 6460 27016
rect 6512 27004 6518 27056
rect 9306 27004 9312 27056
rect 9364 27044 9370 27056
rect 12161 27047 12219 27053
rect 12161 27044 12173 27047
rect 9364 27016 12173 27044
rect 9364 27004 9370 27016
rect 12161 27013 12173 27016
rect 12207 27013 12219 27047
rect 12161 27007 12219 27013
rect 934 26936 940 26988
rect 992 26976 998 26988
rect 1673 26979 1731 26985
rect 1673 26976 1685 26979
rect 992 26948 1685 26976
rect 992 26936 998 26948
rect 1673 26945 1685 26948
rect 1719 26945 1731 26979
rect 1673 26939 1731 26945
rect 11330 26936 11336 26988
rect 11388 26976 11394 26988
rect 11388 26948 12296 26976
rect 11388 26936 11394 26948
rect 12268 26917 12296 26948
rect 12253 26911 12311 26917
rect 12253 26877 12265 26911
rect 12299 26877 12311 26911
rect 12253 26871 12311 26877
rect 11701 26775 11759 26781
rect 11701 26741 11713 26775
rect 11747 26772 11759 26775
rect 16206 26772 16212 26784
rect 11747 26744 16212 26772
rect 11747 26741 11759 26744
rect 11701 26735 11759 26741
rect 16206 26732 16212 26744
rect 16264 26732 16270 26784
rect 1104 26682 49864 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 32950 26682
rect 33002 26630 33014 26682
rect 33066 26630 33078 26682
rect 33130 26630 33142 26682
rect 33194 26630 33206 26682
rect 33258 26630 42950 26682
rect 43002 26630 43014 26682
rect 43066 26630 43078 26682
rect 43130 26630 43142 26682
rect 43194 26630 43206 26682
rect 43258 26630 49864 26682
rect 1104 26608 49864 26630
rect 1854 26392 1860 26444
rect 1912 26392 1918 26444
rect 1578 26324 1584 26376
rect 1636 26324 1642 26376
rect 1104 26138 49864 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 27950 26138
rect 28002 26086 28014 26138
rect 28066 26086 28078 26138
rect 28130 26086 28142 26138
rect 28194 26086 28206 26138
rect 28258 26086 37950 26138
rect 38002 26086 38014 26138
rect 38066 26086 38078 26138
rect 38130 26086 38142 26138
rect 38194 26086 38206 26138
rect 38258 26086 47950 26138
rect 48002 26086 48014 26138
rect 48066 26086 48078 26138
rect 48130 26086 48142 26138
rect 48194 26086 48206 26138
rect 48258 26086 49864 26138
rect 1104 26064 49864 26086
rect 1104 25594 49864 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 32950 25594
rect 33002 25542 33014 25594
rect 33066 25542 33078 25594
rect 33130 25542 33142 25594
rect 33194 25542 33206 25594
rect 33258 25542 42950 25594
rect 43002 25542 43014 25594
rect 43066 25542 43078 25594
rect 43130 25542 43142 25594
rect 43194 25542 43206 25594
rect 43258 25542 49864 25594
rect 1104 25520 49864 25542
rect 10229 25483 10287 25489
rect 10229 25449 10241 25483
rect 10275 25480 10287 25483
rect 12526 25480 12532 25492
rect 10275 25452 12532 25480
rect 10275 25449 10287 25452
rect 10229 25443 10287 25449
rect 12526 25440 12532 25452
rect 12584 25440 12590 25492
rect 1857 25347 1915 25353
rect 1857 25313 1869 25347
rect 1903 25344 1915 25347
rect 4982 25344 4988 25356
rect 1903 25316 4988 25344
rect 1903 25313 1915 25316
rect 1857 25307 1915 25313
rect 4982 25304 4988 25316
rect 5040 25304 5046 25356
rect 10870 25304 10876 25356
rect 10928 25304 10934 25356
rect 934 25236 940 25288
rect 992 25276 998 25288
rect 1581 25279 1639 25285
rect 1581 25276 1593 25279
rect 992 25248 1593 25276
rect 992 25236 998 25248
rect 1581 25245 1593 25248
rect 1627 25245 1639 25279
rect 1581 25239 1639 25245
rect 10597 25279 10655 25285
rect 10597 25245 10609 25279
rect 10643 25276 10655 25279
rect 11609 25279 11667 25285
rect 11609 25276 11621 25279
rect 10643 25248 11621 25276
rect 10643 25245 10655 25248
rect 10597 25239 10655 25245
rect 11609 25245 11621 25248
rect 11655 25245 11667 25279
rect 11609 25239 11667 25245
rect 10318 25100 10324 25152
rect 10376 25140 10382 25152
rect 10689 25143 10747 25149
rect 10689 25140 10701 25143
rect 10376 25112 10701 25140
rect 10376 25100 10382 25112
rect 10689 25109 10701 25112
rect 10735 25109 10747 25143
rect 10689 25103 10747 25109
rect 1104 25050 49864 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 27950 25050
rect 28002 24998 28014 25050
rect 28066 24998 28078 25050
rect 28130 24998 28142 25050
rect 28194 24998 28206 25050
rect 28258 24998 37950 25050
rect 38002 24998 38014 25050
rect 38066 24998 38078 25050
rect 38130 24998 38142 25050
rect 38194 24998 38206 25050
rect 38258 24998 47950 25050
rect 48002 24998 48014 25050
rect 48066 24998 48078 25050
rect 48130 24998 48142 25050
rect 48194 24998 48206 25050
rect 48258 24998 49864 25050
rect 1104 24976 49864 24998
rect 1578 24896 1584 24948
rect 1636 24936 1642 24948
rect 10318 24936 10324 24948
rect 1636 24908 10324 24936
rect 1636 24896 1642 24908
rect 10318 24896 10324 24908
rect 10376 24896 10382 24948
rect 934 24760 940 24812
rect 992 24800 998 24812
rect 1673 24803 1731 24809
rect 1673 24800 1685 24803
rect 992 24772 1685 24800
rect 992 24760 998 24772
rect 1673 24769 1685 24772
rect 1719 24769 1731 24803
rect 1673 24763 1731 24769
rect 1857 24803 1915 24809
rect 1857 24769 1869 24803
rect 1903 24800 1915 24803
rect 4890 24800 4896 24812
rect 1903 24772 4896 24800
rect 1903 24769 1915 24772
rect 1857 24763 1915 24769
rect 4890 24760 4896 24772
rect 4948 24760 4954 24812
rect 33686 24760 33692 24812
rect 33744 24760 33750 24812
rect 24118 24692 24124 24744
rect 24176 24732 24182 24744
rect 24670 24732 24676 24744
rect 24176 24704 24676 24732
rect 24176 24692 24182 24704
rect 24670 24692 24676 24704
rect 24728 24732 24734 24744
rect 32309 24735 32367 24741
rect 32309 24732 32321 24735
rect 24728 24704 32321 24732
rect 24728 24692 24734 24704
rect 32309 24701 32321 24704
rect 32355 24701 32367 24735
rect 32585 24735 32643 24741
rect 32585 24732 32597 24735
rect 32309 24695 32367 24701
rect 32416 24704 32597 24732
rect 26418 24624 26424 24676
rect 26476 24664 26482 24676
rect 32416 24664 32444 24704
rect 32585 24701 32597 24704
rect 32631 24701 32643 24735
rect 32585 24695 32643 24701
rect 34330 24692 34336 24744
rect 34388 24732 34394 24744
rect 47854 24732 47860 24744
rect 34388 24704 47860 24732
rect 34388 24692 34394 24704
rect 47854 24692 47860 24704
rect 47912 24692 47918 24744
rect 26476 24636 32444 24664
rect 26476 24624 26482 24636
rect 10778 24556 10784 24608
rect 10836 24596 10842 24608
rect 10965 24599 11023 24605
rect 10965 24596 10977 24599
rect 10836 24568 10977 24596
rect 10836 24556 10842 24568
rect 10965 24565 10977 24568
rect 11011 24565 11023 24599
rect 10965 24559 11023 24565
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 10413 24395 10471 24401
rect 10413 24361 10425 24395
rect 10459 24392 10471 24395
rect 13906 24392 13912 24404
rect 10459 24364 13912 24392
rect 10459 24361 10471 24364
rect 10413 24355 10471 24361
rect 13906 24352 13912 24364
rect 13964 24352 13970 24404
rect 10965 24259 11023 24265
rect 10965 24225 10977 24259
rect 11011 24256 11023 24259
rect 14826 24256 14832 24268
rect 11011 24228 14832 24256
rect 11011 24225 11023 24228
rect 10965 24219 11023 24225
rect 14826 24216 14832 24228
rect 14884 24216 14890 24268
rect 10778 24148 10784 24200
rect 10836 24148 10842 24200
rect 12434 24148 12440 24200
rect 12492 24148 12498 24200
rect 12802 24148 12808 24200
rect 12860 24188 12866 24200
rect 13814 24188 13820 24200
rect 12860 24160 13820 24188
rect 12860 24148 12866 24160
rect 13814 24148 13820 24160
rect 13872 24148 13878 24200
rect 10870 24012 10876 24064
rect 10928 24012 10934 24064
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 12069 23851 12127 23857
rect 12069 23817 12081 23851
rect 12115 23848 12127 23851
rect 18782 23848 18788 23860
rect 12115 23820 18788 23848
rect 12115 23817 12127 23820
rect 12069 23811 12127 23817
rect 18782 23808 18788 23820
rect 18840 23808 18846 23860
rect 1857 23715 1915 23721
rect 1857 23681 1869 23715
rect 1903 23712 1915 23715
rect 3510 23712 3516 23724
rect 1903 23684 3516 23712
rect 1903 23681 1915 23684
rect 1857 23675 1915 23681
rect 3510 23672 3516 23684
rect 3568 23672 3574 23724
rect 12437 23715 12495 23721
rect 12437 23681 12449 23715
rect 12483 23712 12495 23715
rect 13449 23715 13507 23721
rect 13449 23712 13461 23715
rect 12483 23684 13461 23712
rect 12483 23681 12495 23684
rect 12437 23675 12495 23681
rect 13449 23681 13461 23684
rect 13495 23681 13507 23715
rect 13449 23675 13507 23681
rect 934 23604 940 23656
rect 992 23644 998 23656
rect 1581 23647 1639 23653
rect 1581 23644 1593 23647
rect 992 23616 1593 23644
rect 992 23604 998 23616
rect 1581 23613 1593 23616
rect 1627 23613 1639 23647
rect 1581 23607 1639 23613
rect 12526 23604 12532 23656
rect 12584 23604 12590 23656
rect 12713 23647 12771 23653
rect 12713 23613 12725 23647
rect 12759 23644 12771 23647
rect 17402 23644 17408 23656
rect 12759 23616 17408 23644
rect 12759 23613 12771 23616
rect 12713 23607 12771 23613
rect 17402 23604 17408 23616
rect 17460 23604 17466 23656
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 11885 23307 11943 23313
rect 11885 23273 11897 23307
rect 11931 23304 11943 23307
rect 17586 23304 17592 23316
rect 11931 23276 17592 23304
rect 11931 23273 11943 23276
rect 11885 23267 11943 23273
rect 17586 23264 17592 23276
rect 17644 23264 17650 23316
rect 1857 23171 1915 23177
rect 1857 23137 1869 23171
rect 1903 23168 1915 23171
rect 5902 23168 5908 23180
rect 1903 23140 5908 23168
rect 1903 23137 1915 23140
rect 1857 23131 1915 23137
rect 5902 23128 5908 23140
rect 5960 23128 5966 23180
rect 12529 23171 12587 23177
rect 12529 23137 12541 23171
rect 12575 23168 12587 23171
rect 18322 23168 18328 23180
rect 12575 23140 18328 23168
rect 12575 23137 12587 23140
rect 12529 23131 12587 23137
rect 18322 23128 18328 23140
rect 18380 23128 18386 23180
rect 934 23060 940 23112
rect 992 23100 998 23112
rect 1581 23103 1639 23109
rect 1581 23100 1593 23103
rect 992 23072 1593 23100
rect 992 23060 998 23072
rect 1581 23069 1593 23072
rect 1627 23069 1639 23103
rect 1581 23063 1639 23069
rect 12253 23103 12311 23109
rect 12253 23069 12265 23103
rect 12299 23100 12311 23103
rect 12299 23072 12434 23100
rect 12299 23069 12311 23072
rect 12253 23063 12311 23069
rect 12406 23044 12434 23072
rect 12406 23004 12440 23044
rect 12434 22992 12440 23004
rect 12492 22992 12498 23044
rect 12342 22924 12348 22976
rect 12400 22924 12406 22976
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 1857 22083 1915 22089
rect 1857 22049 1869 22083
rect 1903 22080 1915 22083
rect 3418 22080 3424 22092
rect 1903 22052 3424 22080
rect 1903 22049 1915 22052
rect 1857 22043 1915 22049
rect 3418 22040 3424 22052
rect 3476 22040 3482 22092
rect 934 21972 940 22024
rect 992 22012 998 22024
rect 1581 22015 1639 22021
rect 1581 22012 1593 22015
rect 992 21984 1593 22012
rect 992 21972 998 21984
rect 1581 21981 1593 21984
rect 1627 21981 1639 22015
rect 1581 21975 1639 21981
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 1857 21539 1915 21545
rect 1857 21505 1869 21539
rect 1903 21536 1915 21539
rect 4798 21536 4804 21548
rect 1903 21508 4804 21536
rect 1903 21505 1915 21508
rect 1857 21499 1915 21505
rect 4798 21496 4804 21508
rect 4856 21496 4862 21548
rect 934 21428 940 21480
rect 992 21468 998 21480
rect 1581 21471 1639 21477
rect 1581 21468 1593 21471
rect 992 21440 1593 21468
rect 992 21428 998 21440
rect 1581 21437 1593 21440
rect 1627 21437 1639 21471
rect 1581 21431 1639 21437
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 14277 21063 14335 21069
rect 14277 21029 14289 21063
rect 14323 21060 14335 21063
rect 19150 21060 19156 21072
rect 14323 21032 19156 21060
rect 14323 21029 14335 21032
rect 14277 21023 14335 21029
rect 19150 21020 19156 21032
rect 19208 21020 19214 21072
rect 9398 20884 9404 20936
rect 9456 20924 9462 20936
rect 14461 20927 14519 20933
rect 14461 20924 14473 20927
rect 9456 20896 14473 20924
rect 9456 20884 9462 20896
rect 14461 20893 14473 20896
rect 14507 20893 14519 20927
rect 14461 20887 14519 20893
rect 15102 20884 15108 20936
rect 15160 20924 15166 20936
rect 15841 20927 15899 20933
rect 15841 20924 15853 20927
rect 15160 20896 15853 20924
rect 15160 20884 15166 20896
rect 15841 20893 15853 20896
rect 15887 20893 15899 20927
rect 15841 20887 15899 20893
rect 15657 20791 15715 20797
rect 15657 20757 15669 20791
rect 15703 20788 15715 20791
rect 18598 20788 18604 20800
rect 15703 20760 18604 20788
rect 15703 20757 15715 20760
rect 15657 20751 15715 20757
rect 18598 20748 18604 20760
rect 18656 20748 18662 20800
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 1857 20451 1915 20457
rect 1857 20417 1869 20451
rect 1903 20448 1915 20451
rect 7098 20448 7104 20460
rect 1903 20420 7104 20448
rect 1903 20417 1915 20420
rect 1857 20411 1915 20417
rect 7098 20408 7104 20420
rect 7156 20408 7162 20460
rect 16206 20408 16212 20460
rect 16264 20408 16270 20460
rect 25866 20408 25872 20460
rect 25924 20448 25930 20460
rect 30101 20451 30159 20457
rect 30101 20448 30113 20451
rect 25924 20420 30113 20448
rect 25924 20408 25930 20420
rect 30101 20417 30113 20420
rect 30147 20417 30159 20451
rect 30101 20411 30159 20417
rect 934 20340 940 20392
rect 992 20380 998 20392
rect 1581 20383 1639 20389
rect 1581 20380 1593 20383
rect 992 20352 1593 20380
rect 992 20340 998 20352
rect 1581 20349 1593 20352
rect 1627 20349 1639 20383
rect 1581 20343 1639 20349
rect 30561 20315 30619 20321
rect 30561 20312 30573 20315
rect 26206 20284 30573 20312
rect 16025 20247 16083 20253
rect 16025 20213 16037 20247
rect 16071 20244 16083 20247
rect 18690 20244 18696 20256
rect 16071 20216 18696 20244
rect 16071 20213 16083 20216
rect 16025 20207 16083 20213
rect 18690 20204 18696 20216
rect 18748 20204 18754 20256
rect 23566 20204 23572 20256
rect 23624 20244 23630 20256
rect 26206 20244 26234 20284
rect 30561 20281 30573 20284
rect 30607 20281 30619 20315
rect 30561 20275 30619 20281
rect 23624 20216 26234 20244
rect 30377 20247 30435 20253
rect 23624 20204 23630 20216
rect 30377 20213 30389 20247
rect 30423 20244 30435 20247
rect 34330 20244 34336 20256
rect 30423 20216 34336 20244
rect 30423 20213 30435 20216
rect 30377 20207 30435 20213
rect 34330 20204 34336 20216
rect 34388 20204 34394 20256
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 1854 19932 1860 19984
rect 1912 19932 1918 19984
rect 934 19728 940 19780
rect 992 19768 998 19780
rect 1673 19771 1731 19777
rect 1673 19768 1685 19771
rect 992 19740 1685 19768
rect 992 19728 998 19740
rect 1673 19737 1685 19740
rect 1719 19737 1731 19771
rect 1673 19731 1731 19737
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18952 1639 18955
rect 8386 18952 8392 18964
rect 1627 18924 8392 18952
rect 1627 18921 1639 18924
rect 1581 18915 1639 18921
rect 8386 18912 8392 18924
rect 8444 18912 8450 18964
rect 934 18708 940 18760
rect 992 18748 998 18760
rect 1765 18751 1823 18757
rect 1765 18748 1777 18751
rect 992 18720 1777 18748
rect 992 18708 998 18720
rect 1765 18717 1777 18720
rect 1811 18717 1823 18751
rect 1765 18711 1823 18717
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 1581 18411 1639 18417
rect 1581 18377 1593 18411
rect 1627 18408 1639 18411
rect 8662 18408 8668 18420
rect 1627 18380 8668 18408
rect 1627 18377 1639 18380
rect 1581 18371 1639 18377
rect 8662 18368 8668 18380
rect 8720 18368 8726 18420
rect 1762 18232 1768 18284
rect 1820 18232 1826 18284
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 25406 17688 25412 17740
rect 25464 17688 25470 17740
rect 26142 17688 26148 17740
rect 26200 17728 26206 17740
rect 27709 17731 27767 17737
rect 27709 17728 27721 17731
rect 26200 17700 27721 17728
rect 26200 17688 26206 17700
rect 27709 17697 27721 17700
rect 27755 17697 27767 17731
rect 27709 17691 27767 17697
rect 24946 17620 24952 17672
rect 25004 17620 25010 17672
rect 27246 17620 27252 17672
rect 27304 17620 27310 17672
rect 25130 17552 25136 17604
rect 25188 17552 25194 17604
rect 27433 17595 27491 17601
rect 27433 17592 27445 17595
rect 26206 17564 27445 17592
rect 24486 17484 24492 17536
rect 24544 17524 24550 17536
rect 26206 17524 26234 17564
rect 27433 17561 27445 17564
rect 27479 17561 27491 17595
rect 27433 17555 27491 17561
rect 24544 17496 26234 17524
rect 24544 17484 24550 17496
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 26418 17280 26424 17332
rect 26476 17280 26482 17332
rect 20714 17212 20720 17264
rect 20772 17252 20778 17264
rect 20772 17224 25438 17252
rect 20772 17212 20778 17224
rect 30742 17212 30748 17264
rect 30800 17212 30806 17264
rect 934 17144 940 17196
rect 992 17184 998 17196
rect 1673 17187 1731 17193
rect 1673 17184 1685 17187
rect 992 17156 1685 17184
rect 992 17144 998 17156
rect 1673 17153 1685 17156
rect 1719 17153 1731 17187
rect 1673 17147 1731 17153
rect 17126 17144 17132 17196
rect 17184 17144 17190 17196
rect 17313 17187 17371 17193
rect 17313 17153 17325 17187
rect 17359 17184 17371 17187
rect 23566 17184 23572 17196
rect 17359 17156 23572 17184
rect 17359 17153 17371 17156
rect 17313 17147 17371 17153
rect 1854 17076 1860 17128
rect 1912 17076 1918 17128
rect 15838 17076 15844 17128
rect 15896 17116 15902 17128
rect 17328 17116 17356 17147
rect 23566 17144 23572 17156
rect 23624 17144 23630 17196
rect 24670 17144 24676 17196
rect 24728 17144 24734 17196
rect 24949 17119 25007 17125
rect 24949 17116 24961 17119
rect 15896 17088 17356 17116
rect 24688 17088 24961 17116
rect 15896 17076 15902 17088
rect 24688 17060 24716 17088
rect 24949 17085 24961 17088
rect 24995 17085 25007 17119
rect 24949 17079 25007 17085
rect 28902 17076 28908 17128
rect 28960 17076 28966 17128
rect 29086 17076 29092 17128
rect 29144 17076 29150 17128
rect 24670 17008 24676 17060
rect 24728 17008 24734 17060
rect 17770 16940 17776 16992
rect 17828 16940 17834 16992
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 1857 16711 1915 16717
rect 1857 16677 1869 16711
rect 1903 16708 1915 16711
rect 1946 16708 1952 16720
rect 1903 16680 1952 16708
rect 1903 16677 1915 16680
rect 1857 16671 1915 16677
rect 1946 16668 1952 16680
rect 2004 16668 2010 16720
rect 31018 16600 31024 16652
rect 31076 16600 31082 16652
rect 23566 16532 23572 16584
rect 23624 16581 23630 16584
rect 23624 16575 23662 16581
rect 23650 16541 23662 16575
rect 23624 16535 23662 16541
rect 23707 16575 23765 16581
rect 23707 16541 23719 16575
rect 23753 16572 23765 16575
rect 25130 16572 25136 16584
rect 23753 16544 25136 16572
rect 23753 16541 23765 16544
rect 23707 16535 23765 16541
rect 23624 16532 23630 16535
rect 25130 16532 25136 16544
rect 25188 16532 25194 16584
rect 32858 16532 32864 16584
rect 32916 16532 32922 16584
rect 934 16464 940 16516
rect 992 16504 998 16516
rect 1673 16507 1731 16513
rect 1673 16504 1685 16507
rect 992 16476 1685 16504
rect 992 16464 998 16476
rect 1673 16473 1685 16476
rect 1719 16473 1731 16507
rect 1673 16467 1731 16473
rect 31202 16464 31208 16516
rect 31260 16464 31266 16516
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 26145 15691 26203 15697
rect 26145 15657 26157 15691
rect 26191 15688 26203 15691
rect 26418 15688 26424 15700
rect 26191 15660 26424 15688
rect 26191 15657 26203 15660
rect 26145 15651 26203 15657
rect 26418 15648 26424 15660
rect 26476 15648 26482 15700
rect 1857 15623 1915 15629
rect 1857 15589 1869 15623
rect 1903 15620 1915 15623
rect 7650 15620 7656 15632
rect 1903 15592 7656 15620
rect 1903 15589 1915 15592
rect 1857 15583 1915 15589
rect 7650 15580 7656 15592
rect 7708 15580 7714 15632
rect 25866 15444 25872 15496
rect 25924 15444 25930 15496
rect 934 15376 940 15428
rect 992 15416 998 15428
rect 1673 15419 1731 15425
rect 1673 15416 1685 15419
rect 992 15388 1685 15416
rect 992 15376 998 15388
rect 1673 15385 1685 15388
rect 1719 15385 1731 15419
rect 1673 15379 1731 15385
rect 25958 15308 25964 15360
rect 26016 15348 26022 15360
rect 26329 15351 26387 15357
rect 26329 15348 26341 15351
rect 26016 15320 26341 15348
rect 26016 15308 26022 15320
rect 26329 15317 26341 15320
rect 26375 15317 26387 15351
rect 26329 15311 26387 15317
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 24486 15153 24492 15156
rect 24443 15147 24492 15153
rect 24443 15113 24455 15147
rect 24489 15113 24492 15147
rect 24443 15107 24492 15113
rect 24486 15104 24492 15107
rect 24544 15104 24550 15156
rect 1857 15011 1915 15017
rect 1857 14977 1869 15011
rect 1903 15008 1915 15011
rect 6914 15008 6920 15020
rect 1903 14980 6920 15008
rect 1903 14977 1915 14980
rect 1857 14971 1915 14977
rect 6914 14968 6920 14980
rect 6972 14968 6978 15020
rect 17862 14968 17868 15020
rect 17920 15008 17926 15020
rect 24340 15011 24398 15017
rect 24340 15008 24352 15011
rect 17920 14980 24352 15008
rect 17920 14968 17926 14980
rect 24340 14977 24352 14980
rect 24386 15008 24398 15011
rect 25958 15008 25964 15020
rect 24386 14980 25964 15008
rect 24386 14977 24398 14980
rect 24340 14971 24398 14977
rect 25958 14968 25964 14980
rect 26016 14968 26022 15020
rect 934 14900 940 14952
rect 992 14940 998 14952
rect 1581 14943 1639 14949
rect 1581 14940 1593 14943
rect 992 14912 1593 14940
rect 992 14900 998 14912
rect 1581 14909 1593 14912
rect 1627 14909 1639 14943
rect 1581 14903 1639 14909
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 25038 14356 25044 14408
rect 25096 14396 25102 14408
rect 25260 14399 25318 14405
rect 25260 14396 25272 14399
rect 25096 14368 25272 14396
rect 25096 14356 25102 14368
rect 25260 14365 25272 14368
rect 25306 14365 25318 14399
rect 25260 14359 25318 14365
rect 25363 14263 25421 14269
rect 25363 14229 25375 14263
rect 25409 14260 25421 14263
rect 29086 14260 29092 14272
rect 25409 14232 29092 14260
rect 25409 14229 25421 14232
rect 25363 14223 25421 14229
rect 29086 14220 29092 14232
rect 29144 14220 29150 14272
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 1670 14056 1676 14068
rect 1627 14028 1676 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 1670 14016 1676 14028
rect 1728 14016 1734 14068
rect 19245 14059 19303 14065
rect 19245 14025 19257 14059
rect 19291 14056 19303 14059
rect 20898 14056 20904 14068
rect 19291 14028 20904 14056
rect 19291 14025 19303 14028
rect 19245 14019 19303 14025
rect 20898 14016 20904 14028
rect 20956 14016 20962 14068
rect 21453 14059 21511 14065
rect 21453 14025 21465 14059
rect 21499 14056 21511 14059
rect 24670 14056 24676 14068
rect 21499 14028 24676 14056
rect 21499 14025 21511 14028
rect 21453 14019 21511 14025
rect 24670 14016 24676 14028
rect 24728 14016 24734 14068
rect 27295 14059 27353 14065
rect 27295 14025 27307 14059
rect 27341 14056 27353 14059
rect 31202 14056 31208 14068
rect 27341 14028 31208 14056
rect 27341 14025 27353 14028
rect 27295 14019 27353 14025
rect 31202 14016 31208 14028
rect 31260 14016 31266 14068
rect 20714 13948 20720 14000
rect 20772 13948 20778 14000
rect 934 13880 940 13932
rect 992 13920 998 13932
rect 1765 13923 1823 13929
rect 1765 13920 1777 13923
rect 992 13892 1777 13920
rect 992 13880 998 13892
rect 1765 13889 1777 13892
rect 1811 13889 1823 13923
rect 1765 13883 1823 13889
rect 18598 13880 18604 13932
rect 18656 13880 18662 13932
rect 19702 13880 19708 13932
rect 19760 13880 19766 13932
rect 26694 13880 26700 13932
rect 26752 13920 26758 13932
rect 27192 13923 27250 13929
rect 27192 13920 27204 13923
rect 26752 13892 27204 13920
rect 26752 13880 26758 13892
rect 27192 13889 27204 13892
rect 27238 13889 27250 13923
rect 27192 13883 27250 13889
rect 17218 13812 17224 13864
rect 17276 13852 17282 13864
rect 17862 13852 17868 13864
rect 17276 13824 17868 13852
rect 17276 13812 17282 13824
rect 17862 13812 17868 13824
rect 17920 13852 17926 13864
rect 18785 13855 18843 13861
rect 18785 13852 18797 13855
rect 17920 13824 18797 13852
rect 17920 13812 17926 13824
rect 18785 13821 18797 13824
rect 18831 13821 18843 13855
rect 18785 13815 18843 13821
rect 19968 13719 20026 13725
rect 19968 13685 19980 13719
rect 20014 13716 20026 13719
rect 20622 13716 20628 13728
rect 20014 13688 20628 13716
rect 20014 13685 20026 13688
rect 19968 13679 20026 13685
rect 20622 13676 20628 13688
rect 20680 13676 20686 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 24670 13472 24676 13524
rect 24728 13472 24734 13524
rect 934 13268 940 13320
rect 992 13308 998 13320
rect 1765 13311 1823 13317
rect 1765 13308 1777 13311
rect 992 13280 1777 13308
rect 992 13268 998 13280
rect 1765 13277 1777 13280
rect 1811 13277 1823 13311
rect 1765 13271 1823 13277
rect 23382 13268 23388 13320
rect 23440 13308 23446 13320
rect 24581 13311 24639 13317
rect 24581 13308 24593 13311
rect 23440 13280 24593 13308
rect 23440 13268 23446 13280
rect 24581 13277 24593 13280
rect 24627 13308 24639 13311
rect 25501 13311 25559 13317
rect 25501 13308 25513 13311
rect 24627 13280 25513 13308
rect 24627 13277 24639 13280
rect 24581 13271 24639 13277
rect 25501 13277 25513 13280
rect 25547 13308 25559 13311
rect 25866 13308 25872 13320
rect 25547 13280 25872 13308
rect 25547 13277 25559 13280
rect 25501 13271 25559 13277
rect 25866 13268 25872 13280
rect 25924 13308 25930 13320
rect 25924 13280 26234 13308
rect 25924 13268 25930 13280
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 12710 13172 12716 13184
rect 1627 13144 12716 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 19334 13132 19340 13184
rect 19392 13172 19398 13184
rect 25038 13172 25044 13184
rect 19392 13144 25044 13172
rect 19392 13132 19398 13144
rect 25038 13132 25044 13144
rect 25096 13132 25102 13184
rect 26206 13172 26234 13280
rect 45554 13172 45560 13184
rect 26206 13144 45560 13172
rect 45554 13132 45560 13144
rect 45612 13132 45618 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 18690 12860 18696 12912
rect 18748 12900 18754 12912
rect 18748 12872 20852 12900
rect 18748 12860 18754 12872
rect 19150 12792 19156 12844
rect 19208 12792 19214 12844
rect 20824 12841 20852 12872
rect 20809 12835 20867 12841
rect 20809 12801 20821 12835
rect 20855 12801 20867 12835
rect 20809 12795 20867 12801
rect 19334 12724 19340 12776
rect 19392 12724 19398 12776
rect 20993 12767 21051 12773
rect 20993 12733 21005 12767
rect 21039 12764 21051 12767
rect 21358 12764 21364 12776
rect 21039 12736 21364 12764
rect 21039 12733 21051 12736
rect 20993 12727 21051 12733
rect 21358 12724 21364 12736
rect 21416 12724 21422 12776
rect 19797 12699 19855 12705
rect 19797 12665 19809 12699
rect 19843 12696 19855 12699
rect 22646 12696 22652 12708
rect 19843 12668 22652 12696
rect 19843 12665 19855 12668
rect 19797 12659 19855 12665
rect 22646 12656 22652 12668
rect 22704 12656 22710 12708
rect 21453 12631 21511 12637
rect 21453 12597 21465 12631
rect 21499 12628 21511 12631
rect 24118 12628 24124 12640
rect 21499 12600 24124 12628
rect 21499 12597 21511 12600
rect 21453 12591 21511 12597
rect 24118 12588 24124 12600
rect 24176 12588 24182 12640
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 21358 12384 21364 12436
rect 21416 12424 21422 12436
rect 26694 12424 26700 12436
rect 21416 12396 26700 12424
rect 21416 12384 21422 12396
rect 26694 12384 26700 12396
rect 26752 12384 26758 12436
rect 934 12112 940 12164
rect 992 12152 998 12164
rect 1673 12155 1731 12161
rect 1673 12152 1685 12155
rect 992 12124 1685 12152
rect 992 12112 998 12124
rect 1673 12121 1685 12124
rect 1719 12121 1731 12155
rect 1673 12115 1731 12121
rect 1765 12087 1823 12093
rect 1765 12053 1777 12087
rect 1811 12084 1823 12087
rect 11974 12084 11980 12096
rect 1811 12056 11980 12084
rect 1811 12053 1823 12056
rect 1765 12047 1823 12053
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 1673 11747 1731 11753
rect 1673 11744 1685 11747
rect 992 11716 1685 11744
rect 992 11704 998 11716
rect 1673 11713 1685 11716
rect 1719 11713 1731 11747
rect 1673 11707 1731 11713
rect 1765 11543 1823 11549
rect 1765 11509 1777 11543
rect 1811 11540 1823 11543
rect 10962 11540 10968 11552
rect 1811 11512 10968 11540
rect 1811 11509 1823 11512
rect 1765 11503 1823 11509
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 20622 11296 20628 11348
rect 20680 11336 20686 11348
rect 22097 11339 22155 11345
rect 22097 11336 22109 11339
rect 20680 11308 22109 11336
rect 20680 11296 20686 11308
rect 22097 11305 22109 11308
rect 22143 11305 22155 11339
rect 22097 11299 22155 11305
rect 21358 11160 21364 11212
rect 21416 11200 21422 11212
rect 22465 11203 22523 11209
rect 22465 11200 22477 11203
rect 21416 11172 22477 11200
rect 21416 11160 21422 11172
rect 22465 11169 22477 11172
rect 22511 11169 22523 11203
rect 22465 11163 22523 11169
rect 21545 11135 21603 11141
rect 21545 11101 21557 11135
rect 21591 11132 21603 11135
rect 22005 11135 22063 11141
rect 22005 11132 22017 11135
rect 21591 11104 22017 11132
rect 21591 11101 21603 11104
rect 21545 11095 21603 11101
rect 22005 11101 22017 11104
rect 22051 11132 22063 11135
rect 23382 11132 23388 11144
rect 22051 11104 23388 11132
rect 22051 11101 22063 11104
rect 22005 11095 22063 11101
rect 23382 11092 23388 11104
rect 23440 11092 23446 11144
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 934 10616 940 10668
rect 992 10656 998 10668
rect 1673 10659 1731 10665
rect 1673 10656 1685 10659
rect 992 10628 1685 10656
rect 992 10616 998 10628
rect 1673 10625 1685 10628
rect 1719 10625 1731 10659
rect 1673 10619 1731 10625
rect 1765 10455 1823 10461
rect 1765 10421 1777 10455
rect 1811 10452 1823 10455
rect 12802 10452 12808 10464
rect 1811 10424 12808 10452
rect 1811 10421 1823 10424
rect 1765 10415 1823 10421
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 934 9936 940 9988
rect 992 9976 998 9988
rect 1673 9979 1731 9985
rect 1673 9976 1685 9979
rect 992 9948 1685 9976
rect 992 9936 998 9948
rect 1673 9945 1685 9948
rect 1719 9945 1731 9979
rect 1673 9939 1731 9945
rect 1765 9911 1823 9917
rect 1765 9877 1777 9911
rect 1811 9908 1823 9911
rect 10686 9908 10692 9920
rect 1811 9880 10692 9908
rect 1811 9877 1823 9880
rect 1765 9871 1823 9877
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 1578 9120 1584 9172
rect 1636 9120 1642 9172
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1765 8959 1823 8965
rect 1765 8956 1777 8959
rect 992 8928 1777 8956
rect 992 8916 998 8928
rect 1765 8925 1777 8928
rect 1811 8925 1823 8959
rect 1765 8919 1823 8925
rect 17770 8916 17776 8968
rect 17828 8956 17834 8968
rect 18325 8959 18383 8965
rect 18325 8956 18337 8959
rect 17828 8928 18337 8956
rect 17828 8916 17834 8928
rect 18325 8925 18337 8928
rect 18371 8925 18383 8959
rect 18325 8919 18383 8925
rect 18509 8891 18567 8897
rect 18509 8857 18521 8891
rect 18555 8888 18567 8891
rect 19426 8888 19432 8900
rect 18555 8860 19432 8888
rect 18555 8857 18567 8860
rect 18509 8851 18567 8857
rect 19426 8848 19432 8860
rect 19484 8848 19490 8900
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 1762 8440 1768 8492
rect 1820 8440 1826 8492
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 10870 8344 10876 8356
rect 1627 8316 10876 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 10870 8304 10876 8316
rect 10928 8304 10934 8356
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 13357 8075 13415 8081
rect 13357 8072 13369 8075
rect 6972 8044 13369 8072
rect 6972 8032 6978 8044
rect 13357 8041 13369 8044
rect 13403 8041 13415 8075
rect 13357 8035 13415 8041
rect 9582 7896 9588 7948
rect 9640 7936 9646 7948
rect 10413 7939 10471 7945
rect 10413 7936 10425 7939
rect 9640 7908 10425 7936
rect 9640 7896 9646 7908
rect 10413 7905 10425 7908
rect 10459 7905 10471 7939
rect 20714 7936 20720 7948
rect 10413 7899 10471 7905
rect 11808 7908 20720 7936
rect 11808 7854 11836 7908
rect 20714 7896 20720 7908
rect 20772 7896 20778 7948
rect 13265 7871 13323 7877
rect 13265 7837 13277 7871
rect 13311 7868 13323 7871
rect 15838 7868 15844 7880
rect 13311 7840 15844 7868
rect 13311 7837 13323 7840
rect 13265 7831 13323 7837
rect 15838 7828 15844 7840
rect 15896 7828 15902 7880
rect 10686 7760 10692 7812
rect 10744 7760 10750 7812
rect 20622 7800 20628 7812
rect 12176 7772 20628 7800
rect 12176 7741 12204 7772
rect 20622 7760 20628 7772
rect 20680 7760 20686 7812
rect 12161 7735 12219 7741
rect 12161 7701 12173 7735
rect 12207 7701 12219 7735
rect 12161 7695 12219 7701
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 934 7352 940 7404
rect 992 7392 998 7404
rect 1673 7395 1731 7401
rect 1673 7392 1685 7395
rect 992 7364 1685 7392
rect 992 7352 998 7364
rect 1673 7361 1685 7364
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 1765 7191 1823 7197
rect 1765 7157 1777 7191
rect 1811 7188 1823 7191
rect 10226 7188 10232 7200
rect 1811 7160 10232 7188
rect 1811 7157 1823 7160
rect 1765 7151 1823 7157
rect 10226 7148 10232 7160
rect 10284 7148 10290 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 1857 6851 1915 6857
rect 1857 6817 1869 6851
rect 1903 6848 1915 6851
rect 7742 6848 7748 6860
rect 1903 6820 7748 6848
rect 1903 6817 1915 6820
rect 1857 6811 1915 6817
rect 7742 6808 7748 6820
rect 7800 6808 7806 6860
rect 15013 6783 15071 6789
rect 15013 6749 15025 6783
rect 15059 6780 15071 6783
rect 17218 6780 17224 6792
rect 15059 6752 17224 6780
rect 15059 6749 15071 6752
rect 15013 6743 15071 6749
rect 17218 6740 17224 6752
rect 17276 6740 17282 6792
rect 20898 6740 20904 6792
rect 20956 6740 20962 6792
rect 22646 6740 22652 6792
rect 22704 6740 22710 6792
rect 934 6672 940 6724
rect 992 6712 998 6724
rect 1673 6715 1731 6721
rect 1673 6712 1685 6715
rect 992 6684 1685 6712
rect 992 6672 998 6684
rect 1673 6681 1685 6684
rect 1719 6681 1731 6715
rect 1673 6675 1731 6681
rect 15197 6715 15255 6721
rect 15197 6681 15209 6715
rect 15243 6712 15255 6715
rect 15286 6712 15292 6724
rect 15243 6684 15292 6712
rect 15243 6681 15255 6684
rect 15197 6675 15255 6681
rect 15286 6672 15292 6684
rect 15344 6672 15350 6724
rect 21085 6715 21143 6721
rect 21085 6681 21097 6715
rect 21131 6712 21143 6715
rect 22186 6712 22192 6724
rect 21131 6684 22192 6712
rect 21131 6681 21143 6684
rect 21085 6675 21143 6681
rect 22186 6672 22192 6684
rect 22244 6672 22250 6724
rect 22833 6715 22891 6721
rect 22833 6681 22845 6715
rect 22879 6712 22891 6715
rect 23474 6712 23480 6724
rect 22879 6684 23480 6712
rect 22879 6681 22891 6684
rect 22833 6675 22891 6681
rect 23474 6672 23480 6684
rect 23532 6672 23538 6724
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 16945 6375 17003 6381
rect 16945 6341 16957 6375
rect 16991 6372 17003 6375
rect 19334 6372 19340 6384
rect 16991 6344 19340 6372
rect 16991 6341 17003 6344
rect 16945 6335 17003 6341
rect 19334 6332 19340 6344
rect 19392 6332 19398 6384
rect 24118 6332 24124 6384
rect 24176 6372 24182 6384
rect 25133 6375 25191 6381
rect 25133 6372 25145 6375
rect 24176 6344 25145 6372
rect 24176 6332 24182 6344
rect 25133 6341 25145 6344
rect 25179 6341 25191 6375
rect 25133 6335 25191 6341
rect 25317 6171 25375 6177
rect 25317 6137 25329 6171
rect 25363 6168 25375 6171
rect 28810 6168 28816 6180
rect 25363 6140 28816 6168
rect 25363 6137 25375 6140
rect 25317 6131 25375 6137
rect 28810 6128 28816 6140
rect 28868 6128 28874 6180
rect 15194 6060 15200 6112
rect 15252 6100 15258 6112
rect 17037 6103 17095 6109
rect 17037 6100 17049 6103
rect 15252 6072 17049 6100
rect 15252 6060 15258 6072
rect 17037 6069 17049 6072
rect 17083 6069 17095 6103
rect 17037 6063 17095 6069
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 19521 5695 19579 5701
rect 19521 5661 19533 5695
rect 19567 5692 19579 5695
rect 21358 5692 21364 5704
rect 19567 5664 21364 5692
rect 19567 5661 19579 5664
rect 19521 5655 19579 5661
rect 21358 5652 21364 5664
rect 21416 5652 21422 5704
rect 934 5584 940 5636
rect 992 5624 998 5636
rect 1673 5627 1731 5633
rect 1673 5624 1685 5627
rect 992 5596 1685 5624
rect 992 5584 998 5596
rect 1673 5593 1685 5596
rect 1719 5593 1731 5627
rect 1673 5587 1731 5593
rect 1765 5559 1823 5565
rect 1765 5525 1777 5559
rect 1811 5556 1823 5559
rect 11514 5556 11520 5568
rect 1811 5528 11520 5556
rect 1811 5525 1823 5528
rect 1765 5519 1823 5525
rect 11514 5516 11520 5528
rect 11572 5516 11578 5568
rect 18322 5516 18328 5568
rect 18380 5556 18386 5568
rect 19613 5559 19671 5565
rect 19613 5556 19625 5559
rect 18380 5528 19625 5556
rect 18380 5516 18386 5528
rect 19613 5525 19625 5528
rect 19659 5525 19671 5559
rect 19613 5519 19671 5525
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 1857 5287 1915 5293
rect 1857 5253 1869 5287
rect 1903 5284 1915 5287
rect 9214 5284 9220 5296
rect 1903 5256 9220 5284
rect 1903 5253 1915 5256
rect 1857 5247 1915 5253
rect 9214 5244 9220 5256
rect 9272 5244 9278 5296
rect 934 5176 940 5228
rect 992 5216 998 5228
rect 1673 5219 1731 5225
rect 1673 5216 1685 5219
rect 992 5188 1685 5216
rect 992 5176 998 5188
rect 1673 5185 1685 5188
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 934 4020 940 4072
rect 992 4060 998 4072
rect 1581 4063 1639 4069
rect 1581 4060 1593 4063
rect 992 4032 1593 4060
rect 992 4020 998 4032
rect 1581 4029 1593 4032
rect 1627 4029 1639 4063
rect 1581 4023 1639 4029
rect 1857 4063 1915 4069
rect 1857 4029 1869 4063
rect 1903 4060 1915 4063
rect 12342 4060 12348 4072
rect 1903 4032 12348 4060
rect 1903 4029 1915 4032
rect 1857 4023 1915 4029
rect 12342 4020 12348 4032
rect 12400 4020 12406 4072
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 934 3476 940 3528
rect 992 3516 998 3528
rect 1581 3519 1639 3525
rect 1581 3516 1593 3519
rect 992 3488 1593 3516
rect 992 3476 998 3488
rect 1581 3485 1593 3488
rect 1627 3485 1639 3519
rect 1581 3479 1639 3485
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 12526 3516 12532 3528
rect 1903 3488 12532 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 12526 3476 12532 3488
rect 12584 3476 12590 3528
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 28810 3000 28816 3052
rect 28868 3000 28874 3052
rect 46661 3043 46719 3049
rect 46661 3009 46673 3043
rect 46707 3040 46719 3043
rect 48590 3040 48596 3052
rect 46707 3012 48596 3040
rect 46707 3009 46719 3012
rect 46661 3003 46719 3009
rect 48590 3000 48596 3012
rect 48648 3000 48654 3052
rect 28718 2932 28724 2984
rect 28776 2972 28782 2984
rect 29273 2975 29331 2981
rect 29273 2972 29285 2975
rect 28776 2944 29285 2972
rect 28776 2932 28782 2944
rect 29273 2941 29285 2944
rect 29319 2941 29331 2975
rect 29273 2935 29331 2941
rect 19518 2796 19524 2848
rect 19576 2836 19582 2848
rect 46845 2839 46903 2845
rect 46845 2836 46857 2839
rect 19576 2808 46857 2836
rect 19576 2796 19582 2808
rect 46845 2805 46857 2808
rect 46891 2805 46903 2839
rect 46845 2799 46903 2805
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 31018 2592 31024 2644
rect 31076 2632 31082 2644
rect 31076 2604 42932 2632
rect 31076 2592 31082 2604
rect 24946 2524 24952 2576
rect 25004 2564 25010 2576
rect 25004 2536 26234 2564
rect 25004 2524 25010 2536
rect 5534 2456 5540 2508
rect 5592 2496 5598 2508
rect 7009 2499 7067 2505
rect 7009 2496 7021 2499
rect 5592 2468 7021 2496
rect 5592 2456 5598 2468
rect 7009 2465 7021 2468
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 8846 2456 8852 2508
rect 8904 2496 8910 2508
rect 9677 2499 9735 2505
rect 9677 2496 9689 2499
rect 8904 2468 9689 2496
rect 8904 2456 8910 2468
rect 9677 2465 9689 2468
rect 9723 2465 9735 2499
rect 9677 2459 9735 2465
rect 12158 2456 12164 2508
rect 12216 2496 12222 2508
rect 12713 2499 12771 2505
rect 12713 2496 12725 2499
rect 12216 2468 12725 2496
rect 12216 2456 12222 2468
rect 12713 2465 12725 2468
rect 12759 2465 12771 2499
rect 15194 2496 15200 2508
rect 12713 2459 12771 2465
rect 14384 2468 15200 2496
rect 2222 2388 2228 2440
rect 2280 2428 2286 2440
rect 2501 2431 2559 2437
rect 2501 2428 2513 2431
rect 2280 2400 2513 2428
rect 2280 2388 2286 2400
rect 2501 2397 2513 2400
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 6914 2428 6920 2440
rect 6779 2400 6920 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 6914 2388 6920 2400
rect 6972 2388 6978 2440
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2397 9367 2431
rect 9309 2391 9367 2397
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2428 12403 2431
rect 14384 2428 14412 2468
rect 15194 2456 15200 2468
rect 15252 2456 15258 2508
rect 15470 2456 15476 2508
rect 15528 2456 15534 2508
rect 18782 2456 18788 2508
rect 18840 2496 18846 2508
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 18840 2468 19901 2496
rect 18840 2456 18846 2468
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 22094 2456 22100 2508
rect 22152 2496 22158 2508
rect 22649 2499 22707 2505
rect 22649 2496 22661 2499
rect 22152 2468 22661 2496
rect 22152 2456 22158 2468
rect 22649 2465 22661 2468
rect 22695 2465 22707 2499
rect 22649 2459 22707 2465
rect 25406 2456 25412 2508
rect 25464 2496 25470 2508
rect 25685 2499 25743 2505
rect 25685 2496 25697 2499
rect 25464 2468 25697 2496
rect 25464 2456 25470 2468
rect 25685 2465 25697 2468
rect 25731 2465 25743 2499
rect 26206 2496 26234 2536
rect 28902 2524 28908 2576
rect 28960 2564 28966 2576
rect 28960 2536 35894 2564
rect 28960 2524 28966 2536
rect 32585 2499 32643 2505
rect 32585 2496 32597 2499
rect 26206 2468 32597 2496
rect 25685 2459 25743 2465
rect 32585 2465 32597 2468
rect 32631 2465 32643 2499
rect 35866 2496 35894 2536
rect 42904 2505 42932 2604
rect 45554 2592 45560 2644
rect 45612 2592 45618 2644
rect 38933 2499 38991 2505
rect 38933 2496 38945 2499
rect 35866 2468 38945 2496
rect 32585 2459 32643 2465
rect 38933 2465 38945 2468
rect 38979 2465 38991 2499
rect 38933 2459 38991 2465
rect 42889 2499 42947 2505
rect 42889 2465 42901 2499
rect 42935 2465 42947 2499
rect 42889 2459 42947 2465
rect 12391 2400 14412 2428
rect 15105 2431 15163 2437
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 15105 2397 15117 2431
rect 15151 2428 15163 2431
rect 18322 2428 18328 2440
rect 15151 2400 18328 2428
rect 15151 2397 15163 2400
rect 15105 2391 15163 2397
rect 9324 2360 9352 2391
rect 18322 2388 18328 2400
rect 18380 2388 18386 2440
rect 19426 2388 19432 2440
rect 19484 2388 19490 2440
rect 22186 2388 22192 2440
rect 22244 2388 22250 2440
rect 23474 2388 23480 2440
rect 23532 2428 23538 2440
rect 25225 2431 25283 2437
rect 25225 2428 25237 2431
rect 23532 2400 25237 2428
rect 23532 2388 23538 2400
rect 25225 2397 25237 2400
rect 25271 2397 25283 2431
rect 25225 2391 25283 2397
rect 32030 2388 32036 2440
rect 32088 2428 32094 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 32088 2400 32321 2428
rect 32088 2388 32094 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 35342 2388 35348 2440
rect 35400 2428 35406 2440
rect 35437 2431 35495 2437
rect 35437 2428 35449 2431
rect 35400 2400 35449 2428
rect 35400 2388 35406 2400
rect 35437 2397 35449 2400
rect 35483 2397 35495 2431
rect 35437 2391 35495 2397
rect 35713 2431 35771 2437
rect 35713 2397 35725 2431
rect 35759 2397 35771 2431
rect 35713 2391 35771 2397
rect 15286 2360 15292 2372
rect 9324 2332 15292 2360
rect 15286 2320 15292 2332
rect 15344 2320 15350 2372
rect 27246 2320 27252 2372
rect 27304 2360 27310 2372
rect 35728 2360 35756 2391
rect 38654 2388 38660 2440
rect 38712 2388 38718 2440
rect 41966 2388 41972 2440
rect 42024 2428 42030 2440
rect 42613 2431 42671 2437
rect 42613 2428 42625 2431
rect 42024 2400 42625 2428
rect 42024 2388 42030 2400
rect 42613 2397 42625 2400
rect 42659 2397 42671 2431
rect 42613 2391 42671 2397
rect 27304 2332 35756 2360
rect 27304 2320 27310 2332
rect 45278 2320 45284 2372
rect 45336 2360 45342 2372
rect 45465 2363 45523 2369
rect 45465 2360 45477 2363
rect 45336 2332 45477 2360
rect 45336 2320 45342 2332
rect 45465 2329 45477 2332
rect 45511 2329 45523 2363
rect 45465 2323 45523 2329
rect 2317 2295 2375 2301
rect 2317 2261 2329 2295
rect 2363 2292 2375 2295
rect 10686 2292 10692 2304
rect 2363 2264 10692 2292
rect 2363 2261 2375 2264
rect 2317 2255 2375 2261
rect 10686 2252 10692 2264
rect 10744 2252 10750 2304
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
<< via1 >>
rect 10416 54680 10468 54732
rect 28908 54680 28960 54732
rect 12716 54612 12768 54664
rect 27712 54612 27764 54664
rect 11612 54544 11664 54596
rect 32772 54544 32824 54596
rect 18696 54476 18748 54528
rect 22560 54476 22612 54528
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 27950 54374 28002 54426
rect 28014 54374 28066 54426
rect 28078 54374 28130 54426
rect 28142 54374 28194 54426
rect 28206 54374 28258 54426
rect 37950 54374 38002 54426
rect 38014 54374 38066 54426
rect 38078 54374 38130 54426
rect 38142 54374 38194 54426
rect 38206 54374 38258 54426
rect 47950 54374 48002 54426
rect 48014 54374 48066 54426
rect 48078 54374 48130 54426
rect 48142 54374 48194 54426
rect 48206 54374 48258 54426
rect 19984 54272 20036 54324
rect 22468 54272 22520 54324
rect 22560 54315 22612 54324
rect 22560 54281 22569 54315
rect 22569 54281 22603 54315
rect 22603 54281 22612 54315
rect 22560 54272 22612 54281
rect 22652 54272 22704 54324
rect 23572 54272 23624 54324
rect 27712 54272 27764 54324
rect 28908 54315 28960 54324
rect 28908 54281 28917 54315
rect 28917 54281 28951 54315
rect 28951 54281 28960 54315
rect 28908 54272 28960 54281
rect 32772 54315 32824 54324
rect 32772 54281 32781 54315
rect 32781 54281 32815 54315
rect 32815 54281 32824 54315
rect 32772 54272 32824 54281
rect 3516 54204 3568 54256
rect 8668 54204 8720 54256
rect 10600 54204 10652 54256
rect 13820 54204 13872 54256
rect 15752 54204 15804 54256
rect 18972 54204 19024 54256
rect 20536 54204 20588 54256
rect 2320 54136 2372 54188
rect 4896 54136 4948 54188
rect 7748 54136 7800 54188
rect 10876 54136 10928 54188
rect 12532 54179 12584 54188
rect 12532 54145 12541 54179
rect 12541 54145 12575 54179
rect 12575 54145 12584 54179
rect 12532 54136 12584 54145
rect 12624 54136 12676 54188
rect 17868 54136 17920 54188
rect 19708 54136 19760 54188
rect 5448 54111 5500 54120
rect 5448 54077 5457 54111
rect 5457 54077 5491 54111
rect 5491 54077 5500 54111
rect 5448 54068 5500 54077
rect 10600 54068 10652 54120
rect 20352 54136 20404 54188
rect 22836 54136 22888 54188
rect 23480 54136 23532 54188
rect 24124 54136 24176 54188
rect 24860 54136 24912 54188
rect 25412 54136 25464 54188
rect 26240 54136 26292 54188
rect 26700 54136 26752 54188
rect 27620 54136 27672 54188
rect 28632 54204 28684 54256
rect 29276 54204 29328 54256
rect 30564 54204 30616 54256
rect 20260 54068 20312 54120
rect 16488 54000 16540 54052
rect 22560 54068 22612 54120
rect 22652 54068 22704 54120
rect 28908 54068 28960 54120
rect 30380 54136 30432 54188
rect 32496 54204 32548 54256
rect 33140 54204 33192 54256
rect 33784 54204 33836 54256
rect 34428 54204 34480 54256
rect 37648 54204 37700 54256
rect 38936 54204 38988 54256
rect 42156 54204 42208 54256
rect 35072 54136 35124 54188
rect 35900 54136 35952 54188
rect 39580 54136 39632 54188
rect 44732 54136 44784 54188
rect 45560 54136 45612 54188
rect 46020 54136 46072 54188
rect 47308 54136 47360 54188
rect 47860 54136 47912 54188
rect 18512 53932 18564 53984
rect 22468 53932 22520 53984
rect 27160 53975 27212 53984
rect 27160 53941 27169 53975
rect 27169 53941 27203 53975
rect 27203 53941 27212 53975
rect 27160 53932 27212 53941
rect 29828 53932 29880 53984
rect 30472 53975 30524 53984
rect 30472 53941 30481 53975
rect 30481 53941 30515 53975
rect 30515 53941 30524 53975
rect 30472 53932 30524 53941
rect 31116 53975 31168 53984
rect 31116 53941 31125 53975
rect 31125 53941 31159 53975
rect 31159 53941 31168 53975
rect 31116 53932 31168 53941
rect 33784 54000 33836 54052
rect 38844 54068 38896 54120
rect 40316 54111 40368 54120
rect 40316 54077 40325 54111
rect 40325 54077 40359 54111
rect 40359 54077 40368 54111
rect 40316 54068 40368 54077
rect 34244 53975 34296 53984
rect 34244 53941 34253 53975
rect 34253 53941 34287 53975
rect 34287 53941 34296 53975
rect 34244 53932 34296 53941
rect 35072 53975 35124 53984
rect 35072 53941 35081 53975
rect 35081 53941 35115 53975
rect 35115 53941 35124 53975
rect 35072 53932 35124 53941
rect 37832 53932 37884 53984
rect 43904 53975 43956 53984
rect 43904 53941 43913 53975
rect 43913 53941 43947 53975
rect 43947 53941 43956 53975
rect 43904 53932 43956 53941
rect 45284 53932 45336 53984
rect 46112 53975 46164 53984
rect 46112 53941 46121 53975
rect 46121 53941 46155 53975
rect 46155 53941 46164 53975
rect 46112 53932 46164 53941
rect 46848 53975 46900 53984
rect 46848 53941 46857 53975
rect 46857 53941 46891 53975
rect 46891 53941 46900 53975
rect 46848 53932 46900 53941
rect 47768 53932 47820 53984
rect 48688 53975 48740 53984
rect 48688 53941 48697 53975
rect 48697 53941 48731 53975
rect 48731 53941 48740 53975
rect 48688 53932 48740 53941
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 32950 53830 33002 53882
rect 33014 53830 33066 53882
rect 33078 53830 33130 53882
rect 33142 53830 33194 53882
rect 33206 53830 33258 53882
rect 42950 53830 43002 53882
rect 43014 53830 43066 53882
rect 43078 53830 43130 53882
rect 43142 53830 43194 53882
rect 43206 53830 43258 53882
rect 30380 53728 30432 53780
rect 23480 53660 23532 53712
rect 33508 53660 33560 53712
rect 2872 53635 2924 53644
rect 2872 53601 2881 53635
rect 2881 53601 2915 53635
rect 2915 53601 2924 53635
rect 2872 53592 2924 53601
rect 6092 53635 6144 53644
rect 6092 53601 6101 53635
rect 6101 53601 6135 53635
rect 6135 53601 6144 53635
rect 6092 53592 6144 53601
rect 7840 53635 7892 53644
rect 7840 53601 7849 53635
rect 7849 53601 7883 53635
rect 7883 53601 7892 53635
rect 7840 53592 7892 53601
rect 11244 53635 11296 53644
rect 11244 53601 11253 53635
rect 11253 53601 11287 53635
rect 11287 53601 11296 53635
rect 11244 53592 11296 53601
rect 13360 53635 13412 53644
rect 13360 53601 13369 53635
rect 13369 53601 13403 53635
rect 13403 53601 13412 53635
rect 13360 53592 13412 53601
rect 16396 53635 16448 53644
rect 16396 53601 16405 53635
rect 16405 53601 16439 53635
rect 16439 53601 16448 53635
rect 16396 53592 16448 53601
rect 18328 53635 18380 53644
rect 18328 53601 18337 53635
rect 18337 53601 18371 53635
rect 18371 53601 18380 53635
rect 18328 53592 18380 53601
rect 20904 53592 20956 53644
rect 4712 53524 4764 53576
rect 5540 53524 5592 53576
rect 7380 53567 7432 53576
rect 7380 53533 7389 53567
rect 7389 53533 7423 53567
rect 7423 53533 7432 53567
rect 7380 53524 7432 53533
rect 11704 53524 11756 53576
rect 12348 53567 12400 53576
rect 12348 53533 12357 53567
rect 12357 53533 12391 53567
rect 12391 53533 12400 53567
rect 12348 53524 12400 53533
rect 13820 53524 13872 53576
rect 20812 53524 20864 53576
rect 20996 53567 21048 53576
rect 20996 53533 21005 53567
rect 21005 53533 21039 53567
rect 21039 53533 21048 53567
rect 20996 53524 21048 53533
rect 22192 53524 22244 53576
rect 27804 53524 27856 53576
rect 31208 53524 31260 53576
rect 31852 53524 31904 53576
rect 36360 53524 36412 53576
rect 37004 53524 37056 53576
rect 38292 53524 38344 53576
rect 40224 53524 40276 53576
rect 44088 53524 44140 53576
rect 46664 53524 46716 53576
rect 49240 53592 49292 53644
rect 48596 53524 48648 53576
rect 24860 53456 24912 53508
rect 18420 53388 18472 53440
rect 25044 53388 25096 53440
rect 38660 53499 38712 53508
rect 38660 53465 38669 53499
rect 38669 53465 38703 53499
rect 38703 53465 38712 53499
rect 38660 53456 38712 53465
rect 40040 53388 40092 53440
rect 44364 53431 44416 53440
rect 44364 53397 44373 53431
rect 44373 53397 44407 53431
rect 44407 53397 44416 53431
rect 44364 53388 44416 53397
rect 46940 53431 46992 53440
rect 46940 53397 46949 53431
rect 46949 53397 46983 53431
rect 46983 53397 46992 53431
rect 46940 53388 46992 53397
rect 47032 53388 47084 53440
rect 48872 53431 48924 53440
rect 48872 53397 48881 53431
rect 48881 53397 48915 53431
rect 48915 53397 48924 53431
rect 48872 53388 48924 53397
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 27950 53286 28002 53338
rect 28014 53286 28066 53338
rect 28078 53286 28130 53338
rect 28142 53286 28194 53338
rect 28206 53286 28258 53338
rect 37950 53286 38002 53338
rect 38014 53286 38066 53338
rect 38078 53286 38130 53338
rect 38142 53286 38194 53338
rect 38206 53286 38258 53338
rect 47950 53286 48002 53338
rect 48014 53286 48066 53338
rect 48078 53286 48130 53338
rect 48142 53286 48194 53338
rect 48206 53286 48258 53338
rect 14372 53116 14424 53168
rect 25044 53116 25096 53168
rect 2688 53048 2740 53100
rect 5816 53048 5868 53100
rect 9036 53048 9088 53100
rect 9956 53091 10008 53100
rect 9956 53057 9965 53091
rect 9965 53057 9999 53091
rect 9999 53057 10008 53091
rect 9956 53048 10008 53057
rect 12164 53048 12216 53100
rect 15568 53048 15620 53100
rect 17776 53091 17828 53100
rect 17776 53057 17785 53091
rect 17785 53057 17819 53091
rect 17819 53057 17828 53091
rect 17776 53048 17828 53057
rect 19892 53091 19944 53100
rect 19892 53057 19901 53091
rect 19901 53057 19935 53091
rect 19935 53057 19944 53091
rect 19892 53048 19944 53057
rect 21548 53048 21600 53100
rect 49056 53091 49108 53100
rect 49056 53057 49065 53091
rect 49065 53057 49099 53091
rect 49099 53057 49108 53091
rect 49056 53048 49108 53057
rect 2228 52980 2280 53032
rect 4804 52980 4856 53032
rect 7564 52980 7616 53032
rect 10048 52980 10100 53032
rect 12440 52980 12492 53032
rect 17684 52980 17736 53032
rect 19616 52980 19668 53032
rect 15108 52912 15160 52964
rect 21272 52844 21324 52896
rect 48780 52844 48832 52896
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 32950 52742 33002 52794
rect 33014 52742 33066 52794
rect 33078 52742 33130 52794
rect 33142 52742 33194 52794
rect 33206 52742 33258 52794
rect 42950 52742 43002 52794
rect 43014 52742 43066 52794
rect 43078 52742 43130 52794
rect 43142 52742 43194 52794
rect 43206 52742 43258 52794
rect 2780 52640 2832 52692
rect 14648 52640 14700 52692
rect 20996 52683 21048 52692
rect 20996 52649 21005 52683
rect 21005 52649 21039 52683
rect 21039 52649 21048 52683
rect 20996 52640 21048 52649
rect 1584 52504 1636 52556
rect 8484 52572 8536 52624
rect 49148 52572 49200 52624
rect 4160 52504 4212 52556
rect 6736 52504 6788 52556
rect 9312 52504 9364 52556
rect 11888 52504 11940 52556
rect 14464 52504 14516 52556
rect 17040 52504 17092 52556
rect 4252 52479 4304 52488
rect 4252 52445 4261 52479
rect 4261 52445 4295 52479
rect 4295 52445 4304 52479
rect 4252 52436 4304 52445
rect 9220 52436 9272 52488
rect 9680 52436 9732 52488
rect 11796 52436 11848 52488
rect 14556 52479 14608 52488
rect 14556 52445 14565 52479
rect 14565 52445 14599 52479
rect 14599 52445 14608 52479
rect 14556 52436 14608 52445
rect 16856 52436 16908 52488
rect 21180 52479 21232 52488
rect 21180 52445 21189 52479
rect 21189 52445 21223 52479
rect 21223 52445 21232 52479
rect 21180 52436 21232 52445
rect 49056 52479 49108 52488
rect 49056 52445 49065 52479
rect 49065 52445 49099 52479
rect 49099 52445 49108 52479
rect 49056 52436 49108 52445
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 27950 52198 28002 52250
rect 28014 52198 28066 52250
rect 28078 52198 28130 52250
rect 28142 52198 28194 52250
rect 28206 52198 28258 52250
rect 37950 52198 38002 52250
rect 38014 52198 38066 52250
rect 38078 52198 38130 52250
rect 38142 52198 38194 52250
rect 38206 52198 38258 52250
rect 47950 52198 48002 52250
rect 48014 52198 48066 52250
rect 48078 52198 48130 52250
rect 48142 52198 48194 52250
rect 48206 52198 48258 52250
rect 5816 52096 5868 52148
rect 9680 52139 9732 52148
rect 9680 52105 9689 52139
rect 9689 52105 9723 52139
rect 9723 52105 9732 52139
rect 9680 52096 9732 52105
rect 9956 52096 10008 52148
rect 15568 52139 15620 52148
rect 15568 52105 15577 52139
rect 15577 52105 15611 52139
rect 15611 52105 15620 52139
rect 15568 52096 15620 52105
rect 17776 52096 17828 52148
rect 17868 52096 17920 52148
rect 4896 52028 4948 52080
rect 8392 51960 8444 52012
rect 9864 52003 9916 52012
rect 9864 51969 9873 52003
rect 9873 51969 9907 52003
rect 9907 51969 9916 52003
rect 9864 51960 9916 51969
rect 10508 52003 10560 52012
rect 10508 51969 10517 52003
rect 10517 51969 10551 52003
rect 10551 51969 10560 52003
rect 10508 51960 10560 51969
rect 14464 51960 14516 52012
rect 17684 51960 17736 52012
rect 18972 51960 19024 52012
rect 10692 51892 10744 51944
rect 16304 51756 16356 51808
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 32950 51654 33002 51706
rect 33014 51654 33066 51706
rect 33078 51654 33130 51706
rect 33142 51654 33194 51706
rect 33206 51654 33258 51706
rect 42950 51654 43002 51706
rect 43014 51654 43066 51706
rect 43078 51654 43130 51706
rect 43142 51654 43194 51706
rect 43206 51654 43258 51706
rect 7380 51552 7432 51604
rect 9220 51595 9272 51604
rect 9220 51561 9229 51595
rect 9229 51561 9263 51595
rect 9263 51561 9272 51595
rect 9220 51552 9272 51561
rect 10876 51595 10928 51604
rect 10876 51561 10885 51595
rect 10885 51561 10919 51595
rect 10919 51561 10928 51595
rect 10876 51552 10928 51561
rect 14556 51552 14608 51604
rect 14648 51552 14700 51604
rect 18604 51552 18656 51604
rect 5540 51484 5592 51536
rect 17316 51484 17368 51536
rect 1308 51416 1360 51468
rect 3332 51416 3384 51468
rect 5172 51348 5224 51400
rect 7840 51391 7892 51400
rect 7840 51357 7849 51391
rect 7849 51357 7883 51391
rect 7883 51357 7892 51391
rect 7840 51348 7892 51357
rect 10968 51348 11020 51400
rect 11060 51391 11112 51400
rect 11060 51357 11069 51391
rect 11069 51357 11103 51391
rect 11103 51357 11112 51391
rect 11060 51348 11112 51357
rect 10784 51280 10836 51332
rect 13360 51416 13412 51468
rect 16120 51416 16172 51468
rect 19984 51459 20036 51468
rect 19984 51425 19993 51459
rect 19993 51425 20027 51459
rect 20027 51425 20036 51459
rect 19984 51416 20036 51425
rect 14188 51348 14240 51400
rect 15844 51391 15896 51400
rect 15844 51357 15853 51391
rect 15853 51357 15887 51391
rect 15887 51357 15896 51391
rect 15844 51348 15896 51357
rect 18512 51391 18564 51400
rect 18512 51357 18521 51391
rect 18521 51357 18555 51391
rect 18555 51357 18564 51391
rect 18512 51348 18564 51357
rect 15660 51280 15712 51332
rect 16028 51280 16080 51332
rect 17408 51280 17460 51332
rect 17500 51212 17552 51264
rect 18604 51212 18656 51264
rect 19524 51255 19576 51264
rect 19524 51221 19533 51255
rect 19533 51221 19567 51255
rect 19567 51221 19576 51255
rect 19524 51212 19576 51221
rect 19616 51212 19668 51264
rect 20444 51212 20496 51264
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 27950 51110 28002 51162
rect 28014 51110 28066 51162
rect 28078 51110 28130 51162
rect 28142 51110 28194 51162
rect 28206 51110 28258 51162
rect 37950 51110 38002 51162
rect 38014 51110 38066 51162
rect 38078 51110 38130 51162
rect 38142 51110 38194 51162
rect 38206 51110 38258 51162
rect 47950 51110 48002 51162
rect 48014 51110 48066 51162
rect 48078 51110 48130 51162
rect 48142 51110 48194 51162
rect 48206 51110 48258 51162
rect 7748 51008 7800 51060
rect 9036 51051 9088 51060
rect 9036 51017 9045 51051
rect 9045 51017 9079 51051
rect 9079 51017 9088 51051
rect 9036 51008 9088 51017
rect 12348 51008 12400 51060
rect 12532 51008 12584 51060
rect 14372 50940 14424 50992
rect 3332 50872 3384 50924
rect 7656 50872 7708 50924
rect 9220 50915 9272 50924
rect 9220 50881 9229 50915
rect 9229 50881 9263 50915
rect 9263 50881 9272 50915
rect 9220 50872 9272 50881
rect 12348 50915 12400 50924
rect 12348 50881 12357 50915
rect 12357 50881 12391 50915
rect 12391 50881 12400 50915
rect 12348 50872 12400 50881
rect 12808 50872 12860 50924
rect 1308 50804 1360 50856
rect 14096 50804 14148 50856
rect 15844 51008 15896 51060
rect 15292 50940 15344 50992
rect 17408 51008 17460 51060
rect 17316 50983 17368 50992
rect 17316 50949 17325 50983
rect 17325 50949 17359 50983
rect 17359 50949 17368 50983
rect 17316 50940 17368 50949
rect 20812 51008 20864 51060
rect 23480 51051 23532 51060
rect 23480 51017 23489 51051
rect 23489 51017 23523 51051
rect 23523 51017 23532 51051
rect 23480 51008 23532 51017
rect 33416 51008 33468 51060
rect 22652 50940 22704 50992
rect 43904 50940 43956 50992
rect 17040 50915 17092 50924
rect 17040 50881 17049 50915
rect 17049 50881 17083 50915
rect 17083 50881 17092 50915
rect 17040 50872 17092 50881
rect 18420 50872 18472 50924
rect 19432 50872 19484 50924
rect 20168 50915 20220 50924
rect 20168 50881 20177 50915
rect 20177 50881 20211 50915
rect 20211 50881 20220 50915
rect 20168 50872 20220 50881
rect 21456 50872 21508 50924
rect 21548 50872 21600 50924
rect 26148 50872 26200 50924
rect 16120 50804 16172 50856
rect 17776 50804 17828 50856
rect 20444 50804 20496 50856
rect 20168 50736 20220 50788
rect 23296 50804 23348 50856
rect 37556 50847 37608 50856
rect 37556 50813 37565 50847
rect 37565 50813 37599 50847
rect 37599 50813 37608 50847
rect 37556 50804 37608 50813
rect 47032 50804 47084 50856
rect 13636 50711 13688 50720
rect 13636 50677 13645 50711
rect 13645 50677 13679 50711
rect 13679 50677 13688 50711
rect 13636 50668 13688 50677
rect 15844 50668 15896 50720
rect 16028 50668 16080 50720
rect 17408 50668 17460 50720
rect 19524 50668 19576 50720
rect 22468 50668 22520 50720
rect 24768 50736 24820 50788
rect 24952 50668 25004 50720
rect 27620 50668 27672 50720
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 32950 50566 33002 50618
rect 33014 50566 33066 50618
rect 33078 50566 33130 50618
rect 33142 50566 33194 50618
rect 33206 50566 33258 50618
rect 42950 50566 43002 50618
rect 43014 50566 43066 50618
rect 43078 50566 43130 50618
rect 43142 50566 43194 50618
rect 43206 50566 43258 50618
rect 11704 50507 11756 50516
rect 11704 50473 11713 50507
rect 11713 50473 11747 50507
rect 11747 50473 11756 50507
rect 11704 50464 11756 50473
rect 1584 50396 1636 50448
rect 13636 50396 13688 50448
rect 16120 50507 16172 50516
rect 16120 50473 16129 50507
rect 16129 50473 16163 50507
rect 16163 50473 16172 50507
rect 16120 50464 16172 50473
rect 17592 50464 17644 50516
rect 19616 50464 19668 50516
rect 20076 50464 20128 50516
rect 21548 50464 21600 50516
rect 21732 50464 21784 50516
rect 16856 50396 16908 50448
rect 16212 50328 16264 50380
rect 17408 50371 17460 50380
rect 17408 50337 17417 50371
rect 17417 50337 17451 50371
rect 17451 50337 17460 50371
rect 17408 50328 17460 50337
rect 18604 50328 18656 50380
rect 20076 50328 20128 50380
rect 11888 50303 11940 50312
rect 11888 50269 11897 50303
rect 11897 50269 11931 50303
rect 11931 50269 11940 50303
rect 11888 50260 11940 50269
rect 14096 50260 14148 50312
rect 17040 50260 17092 50312
rect 18972 50260 19024 50312
rect 21548 50328 21600 50380
rect 20904 50303 20956 50312
rect 20904 50269 20913 50303
rect 20913 50269 20947 50303
rect 20947 50269 20956 50303
rect 20904 50260 20956 50269
rect 22652 50328 22704 50380
rect 23388 50260 23440 50312
rect 13636 50192 13688 50244
rect 15200 50192 15252 50244
rect 18420 50192 18472 50244
rect 20076 50235 20128 50244
rect 20076 50201 20085 50235
rect 20085 50201 20119 50235
rect 20119 50201 20128 50235
rect 20076 50192 20128 50201
rect 20260 50192 20312 50244
rect 21456 50192 21508 50244
rect 15568 50124 15620 50176
rect 17776 50124 17828 50176
rect 19616 50124 19668 50176
rect 23572 50192 23624 50244
rect 24860 50260 24912 50312
rect 49056 50303 49108 50312
rect 49056 50269 49065 50303
rect 49065 50269 49099 50303
rect 49099 50269 49108 50303
rect 49056 50260 49108 50269
rect 31208 50192 31260 50244
rect 22652 50167 22704 50176
rect 22652 50133 22661 50167
rect 22661 50133 22695 50167
rect 22695 50133 22704 50167
rect 22652 50124 22704 50133
rect 23664 50167 23716 50176
rect 23664 50133 23673 50167
rect 23673 50133 23707 50167
rect 23707 50133 23716 50167
rect 23664 50124 23716 50133
rect 49240 50167 49292 50176
rect 49240 50133 49249 50167
rect 49249 50133 49283 50167
rect 49283 50133 49292 50167
rect 49240 50124 49292 50133
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 27950 50022 28002 50074
rect 28014 50022 28066 50074
rect 28078 50022 28130 50074
rect 28142 50022 28194 50074
rect 28206 50022 28258 50074
rect 37950 50022 38002 50074
rect 38014 50022 38066 50074
rect 38078 50022 38130 50074
rect 38142 50022 38194 50074
rect 38206 50022 38258 50074
rect 47950 50022 48002 50074
rect 48014 50022 48066 50074
rect 48078 50022 48130 50074
rect 48142 50022 48194 50074
rect 48206 50022 48258 50074
rect 13728 49920 13780 49972
rect 16580 49920 16632 49972
rect 18696 49920 18748 49972
rect 12164 49895 12216 49904
rect 12164 49861 12173 49895
rect 12173 49861 12207 49895
rect 12207 49861 12216 49895
rect 12164 49852 12216 49861
rect 12716 49895 12768 49904
rect 12716 49861 12725 49895
rect 12725 49861 12759 49895
rect 12759 49861 12768 49895
rect 12716 49852 12768 49861
rect 13820 49852 13872 49904
rect 14832 49852 14884 49904
rect 17040 49852 17092 49904
rect 20996 49920 21048 49972
rect 22744 49920 22796 49972
rect 31116 49920 31168 49972
rect 31208 49920 31260 49972
rect 33416 49920 33468 49972
rect 33692 49920 33744 49972
rect 4620 49784 4672 49836
rect 11980 49827 12032 49836
rect 11980 49793 11989 49827
rect 11989 49793 12023 49827
rect 12023 49793 12032 49827
rect 11980 49784 12032 49793
rect 1308 49716 1360 49768
rect 5356 49716 5408 49768
rect 15660 49784 15712 49836
rect 17592 49784 17644 49836
rect 18328 49827 18380 49836
rect 18328 49793 18337 49827
rect 18337 49793 18371 49827
rect 18371 49793 18380 49827
rect 21548 49852 21600 49904
rect 18328 49784 18380 49793
rect 14096 49759 14148 49768
rect 14096 49725 14105 49759
rect 14105 49725 14139 49759
rect 14139 49725 14148 49759
rect 14096 49716 14148 49725
rect 16028 49716 16080 49768
rect 21456 49759 21508 49768
rect 21456 49725 21465 49759
rect 21465 49725 21499 49759
rect 21499 49725 21508 49759
rect 21456 49716 21508 49725
rect 15660 49648 15712 49700
rect 20996 49648 21048 49700
rect 24860 49784 24912 49836
rect 21824 49716 21876 49768
rect 37556 49716 37608 49768
rect 16396 49580 16448 49632
rect 21088 49580 21140 49632
rect 21456 49580 21508 49632
rect 21548 49580 21600 49632
rect 27160 49580 27212 49632
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 32950 49478 33002 49530
rect 33014 49478 33066 49530
rect 33078 49478 33130 49530
rect 33142 49478 33194 49530
rect 33206 49478 33258 49530
rect 42950 49478 43002 49530
rect 43014 49478 43066 49530
rect 43078 49478 43130 49530
rect 43142 49478 43194 49530
rect 43206 49478 43258 49530
rect 9956 49376 10008 49428
rect 11796 49351 11848 49360
rect 11796 49317 11805 49351
rect 11805 49317 11839 49351
rect 11839 49317 11848 49351
rect 11796 49308 11848 49317
rect 12624 49308 12676 49360
rect 1308 49240 1360 49292
rect 3608 49240 3660 49292
rect 15844 49376 15896 49428
rect 16488 49376 16540 49428
rect 13820 49308 13872 49360
rect 3424 49172 3476 49224
rect 13360 49215 13412 49224
rect 13360 49181 13369 49215
rect 13369 49181 13403 49215
rect 13403 49181 13412 49215
rect 13360 49172 13412 49181
rect 14924 49240 14976 49292
rect 15016 49240 15068 49292
rect 16488 49283 16540 49292
rect 16488 49249 16497 49283
rect 16497 49249 16531 49283
rect 16531 49249 16540 49283
rect 16488 49240 16540 49249
rect 14648 49172 14700 49224
rect 18512 49376 18564 49428
rect 21548 49376 21600 49428
rect 21640 49376 21692 49428
rect 18604 49308 18656 49360
rect 19340 49308 19392 49360
rect 19708 49351 19760 49360
rect 19708 49317 19717 49351
rect 19717 49317 19751 49351
rect 19751 49317 19760 49351
rect 19708 49308 19760 49317
rect 17040 49240 17092 49292
rect 17776 49240 17828 49292
rect 18880 49283 18932 49292
rect 18880 49249 18889 49283
rect 18889 49249 18923 49283
rect 18923 49249 18932 49283
rect 18880 49240 18932 49249
rect 19064 49172 19116 49224
rect 21456 49240 21508 49292
rect 22560 49240 22612 49292
rect 26056 49283 26108 49292
rect 26056 49249 26065 49283
rect 26065 49249 26099 49283
rect 26099 49249 26108 49283
rect 26056 49240 26108 49249
rect 23388 49172 23440 49224
rect 30472 49172 30524 49224
rect 9772 49104 9824 49156
rect 12716 49104 12768 49156
rect 13544 49036 13596 49088
rect 14924 49036 14976 49088
rect 16120 49036 16172 49088
rect 18420 49104 18472 49156
rect 18696 49104 18748 49156
rect 17500 49036 17552 49088
rect 17776 49036 17828 49088
rect 23204 49104 23256 49156
rect 22192 49036 22244 49088
rect 22560 49036 22612 49088
rect 24768 49147 24820 49156
rect 24768 49113 24777 49147
rect 24777 49113 24811 49147
rect 24811 49113 24820 49147
rect 24768 49104 24820 49113
rect 25504 49079 25556 49088
rect 25504 49045 25513 49079
rect 25513 49045 25547 49079
rect 25547 49045 25556 49079
rect 25504 49036 25556 49045
rect 25872 49079 25924 49088
rect 25872 49045 25881 49079
rect 25881 49045 25915 49079
rect 25915 49045 25924 49079
rect 25872 49036 25924 49045
rect 33784 49036 33836 49088
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 27950 48934 28002 48986
rect 28014 48934 28066 48986
rect 28078 48934 28130 48986
rect 28142 48934 28194 48986
rect 28206 48934 28258 48986
rect 37950 48934 38002 48986
rect 38014 48934 38066 48986
rect 38078 48934 38130 48986
rect 38142 48934 38194 48986
rect 38206 48934 38258 48986
rect 47950 48934 48002 48986
rect 48014 48934 48066 48986
rect 48078 48934 48130 48986
rect 48142 48934 48194 48986
rect 48206 48934 48258 48986
rect 9220 48832 9272 48884
rect 11244 48696 11296 48748
rect 14096 48832 14148 48884
rect 16304 48832 16356 48884
rect 14740 48764 14792 48816
rect 18604 48764 18656 48816
rect 19892 48832 19944 48884
rect 21088 48832 21140 48884
rect 23296 48832 23348 48884
rect 28908 48832 28960 48884
rect 16120 48696 16172 48748
rect 15016 48628 15068 48680
rect 16212 48671 16264 48680
rect 16212 48637 16221 48671
rect 16221 48637 16255 48671
rect 16255 48637 16264 48671
rect 16212 48628 16264 48637
rect 18512 48696 18564 48748
rect 21272 48764 21324 48816
rect 21456 48764 21508 48816
rect 16672 48560 16724 48612
rect 13360 48492 13412 48544
rect 14648 48492 14700 48544
rect 15200 48492 15252 48544
rect 17316 48535 17368 48544
rect 17316 48501 17325 48535
rect 17325 48501 17359 48535
rect 17359 48501 17368 48535
rect 17316 48492 17368 48501
rect 17500 48560 17552 48612
rect 19156 48628 19208 48680
rect 21916 48696 21968 48748
rect 23388 48696 23440 48748
rect 24860 48696 24912 48748
rect 30748 48696 30800 48748
rect 20260 48628 20312 48680
rect 21456 48628 21508 48680
rect 22376 48628 22428 48680
rect 23664 48628 23716 48680
rect 24768 48628 24820 48680
rect 20720 48492 20772 48544
rect 20996 48535 21048 48544
rect 20996 48501 21005 48535
rect 21005 48501 21039 48535
rect 21039 48501 21048 48535
rect 20996 48492 21048 48501
rect 22468 48492 22520 48544
rect 24952 48492 25004 48544
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 32950 48390 33002 48442
rect 33014 48390 33066 48442
rect 33078 48390 33130 48442
rect 33142 48390 33194 48442
rect 33206 48390 33258 48442
rect 42950 48390 43002 48442
rect 43014 48390 43066 48442
rect 43078 48390 43130 48442
rect 43142 48390 43194 48442
rect 43206 48390 43258 48442
rect 12716 48288 12768 48340
rect 13268 48288 13320 48340
rect 16396 48331 16448 48340
rect 16396 48297 16405 48331
rect 16405 48297 16439 48331
rect 16439 48297 16448 48331
rect 16396 48288 16448 48297
rect 19432 48288 19484 48340
rect 25504 48288 25556 48340
rect 1308 48152 1360 48204
rect 13636 48195 13688 48204
rect 13636 48161 13645 48195
rect 13645 48161 13679 48195
rect 13679 48161 13688 48195
rect 13636 48152 13688 48161
rect 14096 48152 14148 48204
rect 17040 48152 17092 48204
rect 17408 48195 17460 48204
rect 17408 48161 17417 48195
rect 17417 48161 17451 48195
rect 17451 48161 17460 48195
rect 17408 48152 17460 48161
rect 18880 48152 18932 48204
rect 20536 48152 20588 48204
rect 3884 48084 3936 48136
rect 12532 48127 12584 48136
rect 12532 48093 12541 48127
rect 12541 48093 12575 48127
rect 12575 48093 12584 48127
rect 12532 48084 12584 48093
rect 13360 48127 13412 48136
rect 13360 48093 13369 48127
rect 13369 48093 13403 48127
rect 13403 48093 13412 48127
rect 13360 48084 13412 48093
rect 13820 48084 13872 48136
rect 20996 48084 21048 48136
rect 21272 48127 21324 48136
rect 21272 48093 21281 48127
rect 21281 48093 21315 48127
rect 21315 48093 21324 48127
rect 21272 48084 21324 48093
rect 21916 48152 21968 48204
rect 24860 48220 24912 48272
rect 26056 48220 26108 48272
rect 22560 48195 22612 48204
rect 22560 48161 22569 48195
rect 22569 48161 22603 48195
rect 22603 48161 22612 48195
rect 22560 48152 22612 48161
rect 14924 48059 14976 48068
rect 14924 48025 14933 48059
rect 14933 48025 14967 48059
rect 14967 48025 14976 48059
rect 14924 48016 14976 48025
rect 16212 48016 16264 48068
rect 17868 48016 17920 48068
rect 12624 47948 12676 48000
rect 16764 47948 16816 48000
rect 18972 47948 19024 48000
rect 21732 48016 21784 48068
rect 21180 47948 21232 48000
rect 22284 48127 22336 48136
rect 22284 48093 22293 48127
rect 22293 48093 22327 48127
rect 22327 48093 22336 48127
rect 22284 48084 22336 48093
rect 23572 48016 23624 48068
rect 25872 48084 25924 48136
rect 32864 48084 32916 48136
rect 25780 47991 25832 48000
rect 25780 47957 25789 47991
rect 25789 47957 25823 47991
rect 25823 47957 25832 47991
rect 25780 47948 25832 47957
rect 48964 48059 49016 48068
rect 48964 48025 48973 48059
rect 48973 48025 49007 48059
rect 49007 48025 49016 48059
rect 48964 48016 49016 48025
rect 40040 47948 40092 48000
rect 49056 47991 49108 48000
rect 49056 47957 49065 47991
rect 49065 47957 49099 47991
rect 49099 47957 49108 47991
rect 49056 47948 49108 47957
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 27950 47846 28002 47898
rect 28014 47846 28066 47898
rect 28078 47846 28130 47898
rect 28142 47846 28194 47898
rect 28206 47846 28258 47898
rect 37950 47846 38002 47898
rect 38014 47846 38066 47898
rect 38078 47846 38130 47898
rect 38142 47846 38194 47898
rect 38206 47846 38258 47898
rect 47950 47846 48002 47898
rect 48014 47846 48066 47898
rect 48078 47846 48130 47898
rect 48142 47846 48194 47898
rect 48206 47846 48258 47898
rect 9864 47744 9916 47796
rect 10508 47744 10560 47796
rect 10692 47744 10744 47796
rect 12532 47744 12584 47796
rect 19524 47744 19576 47796
rect 4160 47608 4212 47660
rect 9864 47651 9916 47660
rect 9864 47617 9873 47651
rect 9873 47617 9907 47651
rect 9907 47617 9916 47651
rect 9864 47608 9916 47617
rect 11612 47676 11664 47728
rect 13728 47676 13780 47728
rect 1308 47540 1360 47592
rect 14740 47608 14792 47660
rect 12532 47540 12584 47592
rect 8392 47472 8444 47524
rect 13636 47583 13688 47592
rect 13636 47549 13645 47583
rect 13645 47549 13679 47583
rect 13679 47549 13688 47583
rect 13636 47540 13688 47549
rect 14004 47540 14056 47592
rect 16212 47676 16264 47728
rect 17408 47676 17460 47728
rect 17960 47676 18012 47728
rect 22284 47744 22336 47796
rect 15016 47540 15068 47592
rect 20996 47608 21048 47660
rect 30380 47744 30432 47796
rect 48964 47744 49016 47796
rect 49148 47744 49200 47796
rect 23572 47676 23624 47728
rect 26148 47651 26200 47660
rect 26148 47617 26157 47651
rect 26157 47617 26191 47651
rect 26191 47617 26200 47651
rect 26148 47608 26200 47617
rect 17132 47540 17184 47592
rect 18972 47540 19024 47592
rect 20628 47540 20680 47592
rect 20720 47540 20772 47592
rect 17316 47472 17368 47524
rect 24032 47540 24084 47592
rect 24768 47583 24820 47592
rect 24768 47549 24777 47583
rect 24777 47549 24811 47583
rect 24811 47549 24820 47583
rect 24768 47540 24820 47549
rect 14280 47404 14332 47456
rect 14740 47404 14792 47456
rect 17408 47404 17460 47456
rect 19248 47404 19300 47456
rect 24308 47472 24360 47524
rect 21456 47447 21508 47456
rect 21456 47413 21465 47447
rect 21465 47413 21499 47447
rect 21499 47413 21508 47447
rect 21456 47404 21508 47413
rect 22468 47404 22520 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 32950 47302 33002 47354
rect 33014 47302 33066 47354
rect 33078 47302 33130 47354
rect 33142 47302 33194 47354
rect 33206 47302 33258 47354
rect 42950 47302 43002 47354
rect 43014 47302 43066 47354
rect 43078 47302 43130 47354
rect 43142 47302 43194 47354
rect 43206 47302 43258 47354
rect 10784 47200 10836 47252
rect 8760 47132 8812 47184
rect 13544 47200 13596 47252
rect 12716 47132 12768 47184
rect 13912 47132 13964 47184
rect 13636 47107 13688 47116
rect 13636 47073 13645 47107
rect 13645 47073 13679 47107
rect 13679 47073 13688 47107
rect 16304 47200 16356 47252
rect 19064 47200 19116 47252
rect 21640 47200 21692 47252
rect 24032 47243 24084 47252
rect 24032 47209 24041 47243
rect 24041 47209 24075 47243
rect 24075 47209 24084 47243
rect 24032 47200 24084 47209
rect 16028 47175 16080 47184
rect 16028 47141 16037 47175
rect 16037 47141 16071 47175
rect 16071 47141 16080 47175
rect 16028 47132 16080 47141
rect 16396 47132 16448 47184
rect 13636 47064 13688 47073
rect 14280 47107 14332 47116
rect 14280 47073 14289 47107
rect 14289 47073 14323 47107
rect 14323 47073 14332 47107
rect 14280 47064 14332 47073
rect 14556 47064 14608 47116
rect 17408 47107 17460 47116
rect 17408 47073 17417 47107
rect 17417 47073 17451 47107
rect 17451 47073 17460 47107
rect 17408 47064 17460 47073
rect 24860 47064 24912 47116
rect 12440 46996 12492 47048
rect 12532 46996 12584 47048
rect 12900 46928 12952 46980
rect 14004 46996 14056 47048
rect 16028 46996 16080 47048
rect 19616 47039 19668 47048
rect 19616 47005 19625 47039
rect 19625 47005 19659 47039
rect 19659 47005 19668 47039
rect 19616 46996 19668 47005
rect 22284 47039 22336 47048
rect 22284 47005 22293 47039
rect 22293 47005 22327 47039
rect 22327 47005 22336 47039
rect 22284 46996 22336 47005
rect 13360 46903 13412 46912
rect 13360 46869 13369 46903
rect 13369 46869 13403 46903
rect 13403 46869 13412 46903
rect 13360 46860 13412 46869
rect 13912 46928 13964 46980
rect 14648 46928 14700 46980
rect 16212 46928 16264 46980
rect 17868 46928 17920 46980
rect 19248 46928 19300 46980
rect 20904 46928 20956 46980
rect 23572 46928 23624 46980
rect 13544 46860 13596 46912
rect 18328 46860 18380 46912
rect 18788 46860 18840 46912
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 27950 46758 28002 46810
rect 28014 46758 28066 46810
rect 28078 46758 28130 46810
rect 28142 46758 28194 46810
rect 28206 46758 28258 46810
rect 37950 46758 38002 46810
rect 38014 46758 38066 46810
rect 38078 46758 38130 46810
rect 38142 46758 38194 46810
rect 38206 46758 38258 46810
rect 47950 46758 48002 46810
rect 48014 46758 48066 46810
rect 48078 46758 48130 46810
rect 48142 46758 48194 46810
rect 48206 46758 48258 46810
rect 2320 46656 2372 46708
rect 5172 46699 5224 46708
rect 5172 46665 5181 46699
rect 5181 46665 5215 46699
rect 5215 46665 5224 46699
rect 5172 46656 5224 46665
rect 10968 46699 11020 46708
rect 10968 46665 10977 46699
rect 10977 46665 11011 46699
rect 11011 46665 11020 46699
rect 10968 46656 11020 46665
rect 16304 46699 16356 46708
rect 16304 46665 16313 46699
rect 16313 46665 16347 46699
rect 16347 46665 16356 46699
rect 16304 46656 16356 46665
rect 16580 46588 16632 46640
rect 1308 46452 1360 46504
rect 4528 46520 4580 46572
rect 9588 46520 9640 46572
rect 12532 46520 12584 46572
rect 12900 46563 12952 46572
rect 12900 46529 12909 46563
rect 12909 46529 12943 46563
rect 12943 46529 12952 46563
rect 12900 46520 12952 46529
rect 14464 46520 14516 46572
rect 16212 46520 16264 46572
rect 17132 46520 17184 46572
rect 19708 46656 19760 46708
rect 20812 46656 20864 46708
rect 21824 46656 21876 46708
rect 23572 46656 23624 46708
rect 17868 46588 17920 46640
rect 20720 46588 20772 46640
rect 24308 46656 24360 46708
rect 25412 46520 25464 46572
rect 4436 46452 4488 46504
rect 14004 46495 14056 46504
rect 14004 46461 14013 46495
rect 14013 46461 14047 46495
rect 14047 46461 14056 46495
rect 14004 46452 14056 46461
rect 14556 46495 14608 46504
rect 14556 46461 14565 46495
rect 14565 46461 14599 46495
rect 14599 46461 14608 46495
rect 14556 46452 14608 46461
rect 17408 46452 17460 46504
rect 19064 46452 19116 46504
rect 19708 46495 19760 46504
rect 19708 46461 19717 46495
rect 19717 46461 19751 46495
rect 19751 46461 19760 46495
rect 19708 46452 19760 46461
rect 19984 46495 20036 46504
rect 19984 46461 19993 46495
rect 19993 46461 20027 46495
rect 20027 46461 20036 46495
rect 19984 46452 20036 46461
rect 22284 46452 22336 46504
rect 22652 46495 22704 46504
rect 22652 46461 22661 46495
rect 22661 46461 22695 46495
rect 22695 46461 22704 46495
rect 22652 46452 22704 46461
rect 33508 46520 33560 46572
rect 11336 46384 11388 46436
rect 24032 46384 24084 46436
rect 17040 46359 17092 46368
rect 17040 46325 17049 46359
rect 17049 46325 17083 46359
rect 17083 46325 17092 46359
rect 17040 46316 17092 46325
rect 18420 46316 18472 46368
rect 19248 46359 19300 46368
rect 19248 46325 19257 46359
rect 19257 46325 19291 46359
rect 19291 46325 19300 46359
rect 19248 46316 19300 46325
rect 25136 46359 25188 46368
rect 25136 46325 25145 46359
rect 25145 46325 25179 46359
rect 25179 46325 25188 46359
rect 25136 46316 25188 46325
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 32950 46214 33002 46266
rect 33014 46214 33066 46266
rect 33078 46214 33130 46266
rect 33142 46214 33194 46266
rect 33206 46214 33258 46266
rect 42950 46214 43002 46266
rect 43014 46214 43066 46266
rect 43078 46214 43130 46266
rect 43142 46214 43194 46266
rect 43206 46214 43258 46266
rect 3332 46112 3384 46164
rect 7840 46112 7892 46164
rect 11060 46112 11112 46164
rect 13360 46112 13412 46164
rect 14004 46112 14056 46164
rect 14924 46112 14976 46164
rect 17408 46112 17460 46164
rect 21640 46112 21692 46164
rect 1308 45976 1360 46028
rect 16120 45976 16172 46028
rect 17132 46019 17184 46028
rect 17132 45985 17141 46019
rect 17141 45985 17175 46019
rect 17175 45985 17184 46019
rect 17132 45976 17184 45985
rect 19524 45976 19576 46028
rect 19708 45976 19760 46028
rect 20352 45976 20404 46028
rect 24768 45976 24820 46028
rect 3700 45908 3752 45960
rect 7748 45908 7800 45960
rect 11428 45951 11480 45960
rect 11428 45917 11437 45951
rect 11437 45917 11471 45951
rect 11471 45917 11480 45951
rect 11428 45908 11480 45917
rect 14556 45951 14608 45960
rect 14556 45917 14565 45951
rect 14565 45917 14599 45951
rect 14599 45917 14608 45951
rect 14556 45908 14608 45917
rect 19340 45908 19392 45960
rect 22284 45951 22336 45960
rect 22284 45917 22293 45951
rect 22293 45917 22327 45951
rect 22327 45917 22336 45951
rect 22284 45908 22336 45917
rect 47860 45908 47912 45960
rect 49148 45951 49200 45960
rect 49148 45917 49157 45951
rect 49157 45917 49191 45951
rect 49191 45917 49200 45951
rect 49148 45908 49200 45917
rect 5448 45840 5500 45892
rect 16212 45840 16264 45892
rect 17868 45840 17920 45892
rect 20812 45840 20864 45892
rect 23572 45840 23624 45892
rect 15108 45772 15160 45824
rect 19984 45772 20036 45824
rect 22652 45772 22704 45824
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 27950 45670 28002 45722
rect 28014 45670 28066 45722
rect 28078 45670 28130 45722
rect 28142 45670 28194 45722
rect 28206 45670 28258 45722
rect 37950 45670 38002 45722
rect 38014 45670 38066 45722
rect 38078 45670 38130 45722
rect 38142 45670 38194 45722
rect 38206 45670 38258 45722
rect 47950 45670 48002 45722
rect 48014 45670 48066 45722
rect 48078 45670 48130 45722
rect 48142 45670 48194 45722
rect 48206 45670 48258 45722
rect 2688 45543 2740 45552
rect 2688 45509 2697 45543
rect 2697 45509 2731 45543
rect 2731 45509 2740 45543
rect 2688 45500 2740 45509
rect 3884 45543 3936 45552
rect 3884 45509 3893 45543
rect 3893 45509 3927 45543
rect 3927 45509 3936 45543
rect 3884 45500 3936 45509
rect 4620 45543 4672 45552
rect 4620 45509 4629 45543
rect 4629 45509 4663 45543
rect 4663 45509 4672 45543
rect 4620 45500 4672 45509
rect 2504 45475 2556 45484
rect 2504 45441 2513 45475
rect 2513 45441 2547 45475
rect 2547 45441 2556 45475
rect 2504 45432 2556 45441
rect 5724 45432 5776 45484
rect 6828 45432 6880 45484
rect 9128 45432 9180 45484
rect 12624 45500 12676 45552
rect 16028 45500 16080 45552
rect 19432 45568 19484 45620
rect 23756 45568 23808 45620
rect 25412 45568 25464 45620
rect 16672 45500 16724 45552
rect 18788 45500 18840 45552
rect 23572 45500 23624 45552
rect 6184 45364 6236 45416
rect 14648 45432 14700 45484
rect 16488 45432 16540 45484
rect 17408 45475 17460 45484
rect 17408 45441 17417 45475
rect 17417 45441 17451 45475
rect 17451 45441 17460 45475
rect 17408 45432 17460 45441
rect 7656 45296 7708 45348
rect 15200 45364 15252 45416
rect 15936 45364 15988 45416
rect 16120 45407 16172 45416
rect 16120 45373 16129 45407
rect 16129 45373 16163 45407
rect 16163 45373 16172 45407
rect 16120 45364 16172 45373
rect 18328 45364 18380 45416
rect 10876 45296 10928 45348
rect 14188 45296 14240 45348
rect 7012 45228 7064 45280
rect 12808 45228 12860 45280
rect 14464 45296 14516 45348
rect 19156 45296 19208 45348
rect 20352 45364 20404 45416
rect 22284 45364 22336 45416
rect 22836 45407 22888 45416
rect 22836 45373 22845 45407
rect 22845 45373 22879 45407
rect 22879 45373 22888 45407
rect 22836 45364 22888 45373
rect 24308 45364 24360 45416
rect 15016 45228 15068 45280
rect 19248 45228 19300 45280
rect 21456 45296 21508 45348
rect 20812 45228 20864 45280
rect 23572 45228 23624 45280
rect 24584 45271 24636 45280
rect 24584 45237 24593 45271
rect 24593 45237 24627 45271
rect 24627 45237 24636 45271
rect 24584 45228 24636 45237
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 32950 45126 33002 45178
rect 33014 45126 33066 45178
rect 33078 45126 33130 45178
rect 33142 45126 33194 45178
rect 33206 45126 33258 45178
rect 42950 45126 43002 45178
rect 43014 45126 43066 45178
rect 43078 45126 43130 45178
rect 43142 45126 43194 45178
rect 43206 45126 43258 45178
rect 3424 45024 3476 45076
rect 4712 45024 4764 45076
rect 5448 45024 5500 45076
rect 11888 45024 11940 45076
rect 12440 45024 12492 45076
rect 13636 45024 13688 45076
rect 14372 45024 14424 45076
rect 1308 44888 1360 44940
rect 4344 44820 4396 44872
rect 5816 44820 5868 44872
rect 12716 44956 12768 45008
rect 13084 44999 13136 45008
rect 13084 44965 13093 44999
rect 13093 44965 13127 44999
rect 13127 44965 13136 44999
rect 13084 44956 13136 44965
rect 9956 44863 10008 44872
rect 9956 44829 9965 44863
rect 9965 44829 9999 44863
rect 9999 44829 10008 44863
rect 9956 44820 10008 44829
rect 14740 44888 14792 44940
rect 4988 44752 5040 44804
rect 5632 44752 5684 44804
rect 5540 44684 5592 44736
rect 6368 44684 6420 44736
rect 12440 44820 12492 44872
rect 12532 44863 12584 44872
rect 12532 44829 12541 44863
rect 12541 44829 12575 44863
rect 12575 44829 12584 44863
rect 12532 44820 12584 44829
rect 12348 44752 12400 44804
rect 14464 44863 14516 44872
rect 14464 44829 14473 44863
rect 14473 44829 14507 44863
rect 14507 44829 14516 44863
rect 14464 44820 14516 44829
rect 16764 45024 16816 45076
rect 16856 44956 16908 45008
rect 16396 44931 16448 44940
rect 16396 44897 16405 44931
rect 16405 44897 16439 44931
rect 16439 44897 16448 44931
rect 16396 44888 16448 44897
rect 17132 44956 17184 45008
rect 13452 44684 13504 44736
rect 15384 44752 15436 44804
rect 18420 44888 18472 44940
rect 22744 45024 22796 45076
rect 19248 44888 19300 44940
rect 19708 44888 19760 44940
rect 22652 44888 22704 44940
rect 27620 44888 27672 44940
rect 17040 44820 17092 44872
rect 17776 44820 17828 44872
rect 19340 44820 19392 44872
rect 20812 44820 20864 44872
rect 24952 44820 25004 44872
rect 15292 44684 15344 44736
rect 16120 44727 16172 44736
rect 16120 44693 16129 44727
rect 16129 44693 16163 44727
rect 16163 44693 16172 44727
rect 16120 44684 16172 44693
rect 19616 44752 19668 44804
rect 19708 44795 19760 44804
rect 19708 44761 19717 44795
rect 19717 44761 19751 44795
rect 19751 44761 19760 44795
rect 19708 44752 19760 44761
rect 23664 44752 23716 44804
rect 46848 44820 46900 44872
rect 19524 44684 19576 44736
rect 20076 44684 20128 44736
rect 21640 44727 21692 44736
rect 21640 44693 21649 44727
rect 21649 44693 21683 44727
rect 21683 44693 21692 44727
rect 21640 44684 21692 44693
rect 22008 44727 22060 44736
rect 22008 44693 22017 44727
rect 22017 44693 22051 44727
rect 22051 44693 22060 44727
rect 22008 44684 22060 44693
rect 26792 44727 26844 44736
rect 26792 44693 26801 44727
rect 26801 44693 26835 44727
rect 26835 44693 26844 44727
rect 26792 44684 26844 44693
rect 27252 44727 27304 44736
rect 27252 44693 27261 44727
rect 27261 44693 27295 44727
rect 27295 44693 27304 44727
rect 27252 44684 27304 44693
rect 44364 44752 44416 44804
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 27950 44582 28002 44634
rect 28014 44582 28066 44634
rect 28078 44582 28130 44634
rect 28142 44582 28194 44634
rect 28206 44582 28258 44634
rect 37950 44582 38002 44634
rect 38014 44582 38066 44634
rect 38078 44582 38130 44634
rect 38142 44582 38194 44634
rect 38206 44582 38258 44634
rect 47950 44582 48002 44634
rect 48014 44582 48066 44634
rect 48078 44582 48130 44634
rect 48142 44582 48194 44634
rect 48206 44582 48258 44634
rect 4160 44480 4212 44532
rect 6828 44480 6880 44532
rect 11980 44480 12032 44532
rect 13912 44480 13964 44532
rect 17132 44480 17184 44532
rect 18696 44480 18748 44532
rect 4252 44412 4304 44464
rect 5540 44412 5592 44464
rect 9956 44412 10008 44464
rect 10416 44412 10468 44464
rect 2044 44319 2096 44328
rect 2044 44285 2053 44319
rect 2053 44285 2087 44319
rect 2087 44285 2096 44319
rect 2044 44276 2096 44285
rect 3516 44344 3568 44396
rect 8760 44387 8812 44396
rect 8760 44353 8769 44387
rect 8769 44353 8803 44387
rect 8803 44353 8812 44387
rect 8760 44344 8812 44353
rect 10232 44344 10284 44396
rect 13084 44412 13136 44464
rect 19892 44412 19944 44464
rect 12808 44344 12860 44396
rect 16120 44344 16172 44396
rect 4160 44276 4212 44328
rect 17776 44344 17828 44396
rect 19156 44387 19208 44396
rect 19156 44353 19165 44387
rect 19165 44353 19199 44387
rect 19199 44353 19208 44387
rect 19156 44344 19208 44353
rect 23296 44480 23348 44532
rect 20444 44412 20496 44464
rect 23572 44412 23624 44464
rect 23848 44412 23900 44464
rect 20904 44344 20956 44396
rect 22008 44344 22060 44396
rect 22836 44344 22888 44396
rect 18420 44276 18472 44328
rect 19984 44276 20036 44328
rect 13820 44208 13872 44260
rect 19708 44208 19760 44260
rect 20536 44208 20588 44260
rect 27620 44276 27672 44328
rect 9404 44183 9456 44192
rect 9404 44149 9413 44183
rect 9413 44149 9447 44183
rect 9447 44149 9456 44183
rect 9404 44140 9456 44149
rect 10784 44140 10836 44192
rect 12348 44183 12400 44192
rect 12348 44149 12357 44183
rect 12357 44149 12391 44183
rect 12391 44149 12400 44183
rect 12348 44140 12400 44149
rect 21364 44140 21416 44192
rect 25228 44140 25280 44192
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 32950 44038 33002 44090
rect 33014 44038 33066 44090
rect 33078 44038 33130 44090
rect 33142 44038 33194 44090
rect 33206 44038 33258 44090
rect 42950 44038 43002 44090
rect 43014 44038 43066 44090
rect 43078 44038 43130 44090
rect 43142 44038 43194 44090
rect 43206 44038 43258 44090
rect 4436 43936 4488 43988
rect 5816 43936 5868 43988
rect 11244 43979 11296 43988
rect 11244 43945 11253 43979
rect 11253 43945 11287 43979
rect 11287 43945 11296 43979
rect 11244 43936 11296 43945
rect 9680 43868 9732 43920
rect 17684 43979 17736 43988
rect 17684 43945 17693 43979
rect 17693 43945 17727 43979
rect 17727 43945 17736 43979
rect 17684 43936 17736 43945
rect 19156 43936 19208 43988
rect 20904 43979 20956 43988
rect 20904 43945 20913 43979
rect 20913 43945 20947 43979
rect 20947 43945 20956 43979
rect 20904 43936 20956 43945
rect 24032 43979 24084 43988
rect 24032 43945 24041 43979
rect 24041 43945 24075 43979
rect 24075 43945 24084 43979
rect 24032 43936 24084 43945
rect 24952 43936 25004 43988
rect 7288 43800 7340 43852
rect 11796 43843 11848 43852
rect 11796 43809 11805 43843
rect 11805 43809 11839 43843
rect 11839 43809 11848 43843
rect 11796 43800 11848 43809
rect 7012 43732 7064 43784
rect 7656 43732 7708 43784
rect 11336 43732 11388 43784
rect 12532 43732 12584 43784
rect 13820 43800 13872 43852
rect 14004 43800 14056 43852
rect 21640 43868 21692 43920
rect 24860 43868 24912 43920
rect 20076 43843 20128 43852
rect 20076 43809 20085 43843
rect 20085 43809 20119 43843
rect 20119 43809 20128 43843
rect 20076 43800 20128 43809
rect 23572 43800 23624 43852
rect 24584 43800 24636 43852
rect 25228 43843 25280 43852
rect 25228 43809 25237 43843
rect 25237 43809 25271 43843
rect 25271 43809 25280 43843
rect 25228 43800 25280 43809
rect 13912 43732 13964 43784
rect 15016 43732 15068 43784
rect 15200 43732 15252 43784
rect 15476 43775 15528 43784
rect 15476 43741 15485 43775
rect 15485 43741 15519 43775
rect 15519 43741 15528 43775
rect 15476 43732 15528 43741
rect 17224 43732 17276 43784
rect 19892 43775 19944 43784
rect 19892 43741 19901 43775
rect 19901 43741 19935 43775
rect 19935 43741 19944 43775
rect 19892 43732 19944 43741
rect 21824 43775 21876 43784
rect 21824 43741 21833 43775
rect 21833 43741 21867 43775
rect 21867 43741 21876 43775
rect 21824 43732 21876 43741
rect 22284 43775 22336 43784
rect 22284 43741 22293 43775
rect 22293 43741 22327 43775
rect 22327 43741 22336 43775
rect 22284 43732 22336 43741
rect 26792 43732 26844 43784
rect 27620 43800 27672 43852
rect 13360 43664 13412 43716
rect 15752 43707 15804 43716
rect 15752 43673 15761 43707
rect 15761 43673 15795 43707
rect 15795 43673 15804 43707
rect 15752 43664 15804 43673
rect 16028 43664 16080 43716
rect 16212 43664 16264 43716
rect 23848 43664 23900 43716
rect 7472 43596 7524 43648
rect 13268 43596 13320 43648
rect 16672 43596 16724 43648
rect 16764 43596 16816 43648
rect 17316 43596 17368 43648
rect 24584 43639 24636 43648
rect 24584 43605 24593 43639
rect 24593 43605 24627 43639
rect 24627 43605 24636 43639
rect 24584 43596 24636 43605
rect 25780 43596 25832 43648
rect 48596 43664 48648 43716
rect 49240 43596 49292 43648
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 27950 43494 28002 43546
rect 28014 43494 28066 43546
rect 28078 43494 28130 43546
rect 28142 43494 28194 43546
rect 28206 43494 28258 43546
rect 37950 43494 38002 43546
rect 38014 43494 38066 43546
rect 38078 43494 38130 43546
rect 38142 43494 38194 43546
rect 38206 43494 38258 43546
rect 47950 43494 48002 43546
rect 48014 43494 48066 43546
rect 48078 43494 48130 43546
rect 48142 43494 48194 43546
rect 48206 43494 48258 43546
rect 9772 43435 9824 43444
rect 9772 43401 9781 43435
rect 9781 43401 9815 43435
rect 9815 43401 9824 43435
rect 9772 43392 9824 43401
rect 9864 43392 9916 43444
rect 10784 43435 10836 43444
rect 10784 43401 10793 43435
rect 10793 43401 10827 43435
rect 10827 43401 10836 43435
rect 10784 43392 10836 43401
rect 11428 43392 11480 43444
rect 12348 43392 12400 43444
rect 12532 43324 12584 43376
rect 5356 43256 5408 43308
rect 9220 43256 9272 43308
rect 10048 43256 10100 43308
rect 1308 43188 1360 43240
rect 5080 43188 5132 43240
rect 10968 43231 11020 43240
rect 10968 43197 10977 43231
rect 10977 43197 11011 43231
rect 11011 43197 11020 43231
rect 10968 43188 11020 43197
rect 12164 43231 12216 43240
rect 12164 43197 12173 43231
rect 12173 43197 12207 43231
rect 12207 43197 12216 43231
rect 12164 43188 12216 43197
rect 12256 43231 12308 43240
rect 12256 43197 12265 43231
rect 12265 43197 12299 43231
rect 12299 43197 12308 43231
rect 12256 43188 12308 43197
rect 13544 43392 13596 43444
rect 17684 43392 17736 43444
rect 17868 43392 17920 43444
rect 17316 43324 17368 43376
rect 14004 43256 14056 43308
rect 14924 43256 14976 43308
rect 15844 43256 15896 43308
rect 17040 43299 17092 43308
rect 17040 43265 17049 43299
rect 17049 43265 17083 43299
rect 17083 43265 17092 43299
rect 17040 43256 17092 43265
rect 17592 43256 17644 43308
rect 9772 43120 9824 43172
rect 11520 43120 11572 43172
rect 9220 43095 9272 43104
rect 9220 43061 9229 43095
rect 9229 43061 9263 43095
rect 9263 43061 9272 43095
rect 9220 43052 9272 43061
rect 9588 43052 9640 43104
rect 15476 43188 15528 43240
rect 18328 43324 18380 43376
rect 19708 43392 19760 43444
rect 21272 43392 21324 43444
rect 21824 43392 21876 43444
rect 22468 43435 22520 43444
rect 22468 43401 22477 43435
rect 22477 43401 22511 43435
rect 22511 43401 22520 43435
rect 22468 43392 22520 43401
rect 24584 43324 24636 43376
rect 20812 43256 20864 43308
rect 17316 43120 17368 43172
rect 21364 43231 21416 43240
rect 21364 43197 21373 43231
rect 21373 43197 21407 43231
rect 21407 43197 21416 43231
rect 21364 43188 21416 43197
rect 23572 43188 23624 43240
rect 15568 43052 15620 43104
rect 16672 43052 16724 43104
rect 17868 43052 17920 43104
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 32950 42950 33002 43002
rect 33014 42950 33066 43002
rect 33078 42950 33130 43002
rect 33142 42950 33194 43002
rect 33206 42950 33258 43002
rect 42950 42950 43002 43002
rect 43014 42950 43066 43002
rect 43078 42950 43130 43002
rect 43142 42950 43194 43002
rect 43206 42950 43258 43002
rect 8944 42848 8996 42900
rect 11796 42848 11848 42900
rect 14188 42848 14240 42900
rect 16764 42848 16816 42900
rect 20260 42848 20312 42900
rect 24032 42848 24084 42900
rect 1308 42712 1360 42764
rect 3700 42712 3752 42764
rect 1584 42687 1636 42696
rect 1584 42653 1593 42687
rect 1593 42653 1627 42687
rect 1627 42653 1636 42687
rect 1584 42644 1636 42653
rect 5632 42644 5684 42696
rect 6000 42644 6052 42696
rect 9312 42687 9364 42696
rect 9312 42653 9321 42687
rect 9321 42653 9355 42687
rect 9355 42653 9364 42687
rect 9312 42644 9364 42653
rect 15200 42712 15252 42764
rect 17316 42712 17368 42764
rect 19984 42755 20036 42764
rect 19984 42721 19993 42755
rect 19993 42721 20027 42755
rect 20027 42721 20036 42755
rect 19984 42712 20036 42721
rect 21456 42712 21508 42764
rect 21732 42712 21784 42764
rect 7564 42576 7616 42628
rect 7012 42508 7064 42560
rect 8484 42551 8536 42560
rect 8484 42517 8493 42551
rect 8493 42517 8527 42551
rect 8527 42517 8536 42551
rect 8484 42508 8536 42517
rect 8760 42576 8812 42628
rect 15476 42644 15528 42696
rect 18328 42644 18380 42696
rect 18512 42644 18564 42696
rect 22928 42712 22980 42764
rect 48780 42712 48832 42764
rect 25136 42644 25188 42696
rect 10324 42576 10376 42628
rect 11336 42576 11388 42628
rect 12716 42576 12768 42628
rect 13820 42576 13872 42628
rect 16028 42576 16080 42628
rect 18696 42619 18748 42628
rect 18696 42585 18705 42619
rect 18705 42585 18739 42619
rect 18739 42585 18748 42619
rect 18696 42576 18748 42585
rect 22468 42576 22520 42628
rect 23848 42576 23900 42628
rect 13636 42508 13688 42560
rect 13912 42508 13964 42560
rect 18512 42508 18564 42560
rect 18788 42551 18840 42560
rect 18788 42517 18797 42551
rect 18797 42517 18831 42551
rect 18831 42517 18840 42551
rect 18788 42508 18840 42517
rect 18972 42508 19024 42560
rect 19800 42551 19852 42560
rect 19800 42517 19809 42551
rect 19809 42517 19843 42551
rect 19843 42517 19852 42551
rect 19800 42508 19852 42517
rect 21732 42508 21784 42560
rect 21916 42508 21968 42560
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 27950 42406 28002 42458
rect 28014 42406 28066 42458
rect 28078 42406 28130 42458
rect 28142 42406 28194 42458
rect 28206 42406 28258 42458
rect 37950 42406 38002 42458
rect 38014 42406 38066 42458
rect 38078 42406 38130 42458
rect 38142 42406 38194 42458
rect 38206 42406 38258 42458
rect 47950 42406 48002 42458
rect 48014 42406 48066 42458
rect 48078 42406 48130 42458
rect 48142 42406 48194 42458
rect 48206 42406 48258 42458
rect 4160 42304 4212 42356
rect 9312 42304 9364 42356
rect 12440 42304 12492 42356
rect 15200 42304 15252 42356
rect 15752 42304 15804 42356
rect 18328 42304 18380 42356
rect 18512 42304 18564 42356
rect 21088 42347 21140 42356
rect 21088 42313 21097 42347
rect 21097 42313 21131 42347
rect 21131 42313 21140 42347
rect 21088 42304 21140 42313
rect 21364 42304 21416 42356
rect 21824 42304 21876 42356
rect 15108 42236 15160 42288
rect 16396 42236 16448 42288
rect 19708 42236 19760 42288
rect 20076 42236 20128 42288
rect 21916 42236 21968 42288
rect 8760 42211 8812 42220
rect 8760 42177 8769 42211
rect 8769 42177 8803 42211
rect 8803 42177 8812 42211
rect 8760 42168 8812 42177
rect 11060 42168 11112 42220
rect 11152 42211 11204 42220
rect 11152 42177 11161 42211
rect 11161 42177 11195 42211
rect 11195 42177 11204 42211
rect 11152 42168 11204 42177
rect 12164 42168 12216 42220
rect 15936 42168 15988 42220
rect 16764 42168 16816 42220
rect 17500 42168 17552 42220
rect 19800 42168 19852 42220
rect 9036 42143 9088 42152
rect 9036 42109 9045 42143
rect 9045 42109 9079 42143
rect 9079 42109 9088 42143
rect 9036 42100 9088 42109
rect 10416 42100 10468 42152
rect 13544 42143 13596 42152
rect 13544 42109 13553 42143
rect 13553 42109 13587 42143
rect 13587 42109 13596 42143
rect 13544 42100 13596 42109
rect 7104 42032 7156 42084
rect 8484 41964 8536 42016
rect 8668 41964 8720 42016
rect 10508 42075 10560 42084
rect 10508 42041 10517 42075
rect 10517 42041 10551 42075
rect 10551 42041 10560 42075
rect 10508 42032 10560 42041
rect 11612 42032 11664 42084
rect 11980 41964 12032 42016
rect 14556 42143 14608 42152
rect 14556 42109 14565 42143
rect 14565 42109 14599 42143
rect 14599 42109 14608 42143
rect 14556 42100 14608 42109
rect 14832 42143 14884 42152
rect 14832 42109 14841 42143
rect 14841 42109 14875 42143
rect 14875 42109 14884 42143
rect 14832 42100 14884 42109
rect 17224 42100 17276 42152
rect 16028 42032 16080 42084
rect 17868 42100 17920 42152
rect 18144 42100 18196 42152
rect 18512 42100 18564 42152
rect 18696 42100 18748 42152
rect 20168 42168 20220 42220
rect 20352 42168 20404 42220
rect 17684 42032 17736 42084
rect 20260 42100 20312 42152
rect 21364 42168 21416 42220
rect 22928 42236 22980 42288
rect 22284 42168 22336 42220
rect 23756 42168 23808 42220
rect 20904 42032 20956 42084
rect 21456 42100 21508 42152
rect 22652 42143 22704 42152
rect 22652 42109 22661 42143
rect 22661 42109 22695 42143
rect 22695 42109 22704 42143
rect 22652 42100 22704 42109
rect 25228 42100 25280 42152
rect 13728 41964 13780 42016
rect 14280 41964 14332 42016
rect 15568 41964 15620 42016
rect 17960 41964 18012 42016
rect 19248 41964 19300 42016
rect 19708 41964 19760 42016
rect 22376 42032 22428 42084
rect 24676 42032 24728 42084
rect 48964 42032 49016 42084
rect 21088 41964 21140 42016
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 32950 41862 33002 41914
rect 33014 41862 33066 41914
rect 33078 41862 33130 41914
rect 33142 41862 33194 41914
rect 33206 41862 33258 41914
rect 42950 41862 43002 41914
rect 43014 41862 43066 41914
rect 43078 41862 43130 41914
rect 43142 41862 43194 41914
rect 43206 41862 43258 41914
rect 4344 41760 4396 41812
rect 1768 41692 1820 41744
rect 1308 41624 1360 41676
rect 9404 41624 9456 41676
rect 10876 41760 10928 41812
rect 11152 41760 11204 41812
rect 7012 41556 7064 41608
rect 8300 41556 8352 41608
rect 10416 41667 10468 41676
rect 10416 41633 10425 41667
rect 10425 41633 10459 41667
rect 10459 41633 10468 41667
rect 10416 41624 10468 41633
rect 11980 41692 12032 41744
rect 12624 41760 12676 41812
rect 11888 41624 11940 41676
rect 9772 41599 9824 41608
rect 9772 41565 9781 41599
rect 9781 41565 9815 41599
rect 9815 41565 9824 41599
rect 9772 41556 9824 41565
rect 12716 41556 12768 41608
rect 10600 41488 10652 41540
rect 17960 41760 18012 41812
rect 20812 41760 20864 41812
rect 20996 41803 21048 41812
rect 20996 41769 21005 41803
rect 21005 41769 21039 41803
rect 21039 41769 21048 41803
rect 20996 41760 21048 41769
rect 22376 41760 22428 41812
rect 24952 41760 25004 41812
rect 14280 41735 14332 41744
rect 14280 41701 14289 41735
rect 14289 41701 14323 41735
rect 14323 41701 14332 41735
rect 14280 41692 14332 41701
rect 14096 41624 14148 41676
rect 15384 41692 15436 41744
rect 17224 41735 17276 41744
rect 17224 41701 17233 41735
rect 17233 41701 17267 41735
rect 17267 41701 17276 41735
rect 17224 41692 17276 41701
rect 17500 41692 17552 41744
rect 18144 41692 18196 41744
rect 14740 41667 14792 41676
rect 14740 41633 14749 41667
rect 14749 41633 14783 41667
rect 14783 41633 14792 41667
rect 14740 41624 14792 41633
rect 15752 41667 15804 41676
rect 15752 41633 15761 41667
rect 15761 41633 15795 41667
rect 15795 41633 15804 41667
rect 15752 41624 15804 41633
rect 18236 41624 18288 41676
rect 22652 41692 22704 41744
rect 14556 41556 14608 41608
rect 18328 41556 18380 41608
rect 5540 41420 5592 41472
rect 12256 41420 12308 41472
rect 22100 41624 22152 41676
rect 20720 41599 20772 41608
rect 20720 41565 20729 41599
rect 20729 41565 20763 41599
rect 20763 41565 20772 41599
rect 20720 41556 20772 41565
rect 20996 41556 21048 41608
rect 24860 41692 24912 41744
rect 23572 41624 23624 41676
rect 23848 41667 23900 41676
rect 23848 41633 23857 41667
rect 23857 41633 23891 41667
rect 23891 41633 23900 41667
rect 23848 41624 23900 41633
rect 15936 41420 15988 41472
rect 16120 41420 16172 41472
rect 23664 41599 23716 41608
rect 23664 41565 23673 41599
rect 23673 41565 23707 41599
rect 23707 41565 23716 41599
rect 23664 41556 23716 41565
rect 22192 41488 22244 41540
rect 24492 41488 24544 41540
rect 17500 41420 17552 41472
rect 20352 41420 20404 41472
rect 20904 41420 20956 41472
rect 21272 41420 21324 41472
rect 21364 41463 21416 41472
rect 21364 41429 21373 41463
rect 21373 41429 21407 41463
rect 21407 41429 21416 41463
rect 21364 41420 21416 41429
rect 21640 41420 21692 41472
rect 23756 41463 23808 41472
rect 23756 41429 23765 41463
rect 23765 41429 23799 41463
rect 23799 41429 23808 41463
rect 23756 41420 23808 41429
rect 27252 41420 27304 41472
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 27950 41318 28002 41370
rect 28014 41318 28066 41370
rect 28078 41318 28130 41370
rect 28142 41318 28194 41370
rect 28206 41318 28258 41370
rect 37950 41318 38002 41370
rect 38014 41318 38066 41370
rect 38078 41318 38130 41370
rect 38142 41318 38194 41370
rect 38206 41318 38258 41370
rect 47950 41318 48002 41370
rect 48014 41318 48066 41370
rect 48078 41318 48130 41370
rect 48142 41318 48194 41370
rect 48206 41318 48258 41370
rect 10324 41216 10376 41268
rect 11520 41216 11572 41268
rect 12072 41216 12124 41268
rect 9220 41148 9272 41200
rect 11336 41148 11388 41200
rect 7840 41080 7892 41132
rect 8484 41080 8536 41132
rect 11704 41080 11756 41132
rect 14556 41216 14608 41268
rect 15752 41216 15804 41268
rect 16488 41216 16540 41268
rect 19248 41259 19300 41268
rect 19248 41225 19257 41259
rect 19257 41225 19291 41259
rect 19291 41225 19300 41259
rect 19248 41216 19300 41225
rect 24400 41216 24452 41268
rect 24492 41259 24544 41268
rect 24492 41225 24501 41259
rect 24501 41225 24535 41259
rect 24535 41225 24544 41259
rect 24492 41216 24544 41225
rect 24860 41259 24912 41268
rect 24860 41225 24869 41259
rect 24869 41225 24903 41259
rect 24903 41225 24912 41259
rect 24860 41216 24912 41225
rect 24952 41259 25004 41268
rect 24952 41225 24961 41259
rect 24961 41225 24995 41259
rect 24995 41225 25004 41259
rect 24952 41216 25004 41225
rect 12716 41148 12768 41200
rect 15936 41080 15988 41132
rect 16488 41080 16540 41132
rect 1308 41012 1360 41064
rect 8576 41012 8628 41064
rect 12256 41012 12308 41064
rect 6920 40987 6972 40996
rect 6920 40953 6929 40987
rect 6929 40953 6963 40987
rect 6963 40953 6972 40987
rect 6920 40944 6972 40953
rect 11336 40944 11388 40996
rect 13636 41012 13688 41064
rect 14096 41055 14148 41064
rect 14096 41021 14105 41055
rect 14105 41021 14139 41055
rect 14139 41021 14148 41055
rect 14096 41012 14148 41021
rect 14188 41012 14240 41064
rect 16304 41012 16356 41064
rect 8208 40876 8260 40928
rect 10692 40876 10744 40928
rect 10876 40876 10928 40928
rect 11888 40919 11940 40928
rect 11888 40885 11897 40919
rect 11897 40885 11931 40919
rect 11931 40885 11940 40919
rect 11888 40876 11940 40885
rect 13636 40876 13688 40928
rect 19524 41148 19576 41200
rect 22192 41148 22244 41200
rect 23204 41148 23256 41200
rect 46112 41216 46164 41268
rect 17868 41012 17920 41064
rect 17500 40876 17552 40928
rect 23388 41080 23440 41132
rect 18788 41012 18840 41064
rect 19616 41012 19668 41064
rect 23940 41080 23992 41132
rect 19524 40944 19576 40996
rect 23848 41012 23900 41064
rect 23480 40944 23532 40996
rect 22652 40876 22704 40928
rect 23204 40876 23256 40928
rect 47768 41080 47820 41132
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 32950 40774 33002 40826
rect 33014 40774 33066 40826
rect 33078 40774 33130 40826
rect 33142 40774 33194 40826
rect 33206 40774 33258 40826
rect 42950 40774 43002 40826
rect 43014 40774 43066 40826
rect 43078 40774 43130 40826
rect 43142 40774 43194 40826
rect 43206 40774 43258 40826
rect 7748 40672 7800 40724
rect 9128 40715 9180 40724
rect 9128 40681 9137 40715
rect 9137 40681 9171 40715
rect 9171 40681 9180 40715
rect 9128 40672 9180 40681
rect 10692 40672 10744 40724
rect 11980 40715 12032 40724
rect 11980 40681 11989 40715
rect 11989 40681 12023 40715
rect 12023 40681 12032 40715
rect 11980 40672 12032 40681
rect 12532 40672 12584 40724
rect 9036 40536 9088 40588
rect 9312 40536 9364 40588
rect 8300 40468 8352 40520
rect 8484 40468 8536 40520
rect 8760 40400 8812 40452
rect 12716 40468 12768 40520
rect 12992 40536 13044 40588
rect 14556 40536 14608 40588
rect 10416 40400 10468 40452
rect 7748 40332 7800 40384
rect 8392 40332 8444 40384
rect 11244 40400 11296 40452
rect 13268 40400 13320 40452
rect 14096 40400 14148 40452
rect 15936 40400 15988 40452
rect 14188 40332 14240 40384
rect 16120 40332 16172 40384
rect 19984 40672 20036 40724
rect 20628 40672 20680 40724
rect 23664 40672 23716 40724
rect 24400 40672 24452 40724
rect 49056 40672 49108 40724
rect 19064 40604 19116 40656
rect 19708 40536 19760 40588
rect 21824 40579 21876 40588
rect 21824 40545 21833 40579
rect 21833 40545 21867 40579
rect 21867 40545 21876 40579
rect 21824 40536 21876 40545
rect 24768 40536 24820 40588
rect 19156 40468 19208 40520
rect 21548 40511 21600 40520
rect 21548 40477 21557 40511
rect 21557 40477 21591 40511
rect 21591 40477 21600 40511
rect 21548 40468 21600 40477
rect 23756 40468 23808 40520
rect 18880 40443 18932 40452
rect 18880 40409 18889 40443
rect 18889 40409 18923 40443
rect 18923 40409 18932 40443
rect 18880 40400 18932 40409
rect 18788 40332 18840 40384
rect 19800 40375 19852 40384
rect 19800 40341 19809 40375
rect 19809 40341 19843 40375
rect 19843 40341 19852 40375
rect 19800 40332 19852 40341
rect 20352 40375 20404 40384
rect 20352 40341 20361 40375
rect 20361 40341 20395 40375
rect 20395 40341 20404 40375
rect 20352 40332 20404 40341
rect 20904 40400 20956 40452
rect 21272 40400 21324 40452
rect 22284 40400 22336 40452
rect 23480 40400 23532 40452
rect 23664 40400 23716 40452
rect 20628 40332 20680 40384
rect 22836 40332 22888 40384
rect 23296 40375 23348 40384
rect 23296 40341 23305 40375
rect 23305 40341 23339 40375
rect 23339 40341 23348 40375
rect 23296 40332 23348 40341
rect 24584 40375 24636 40384
rect 24584 40341 24593 40375
rect 24593 40341 24627 40375
rect 24627 40341 24636 40375
rect 24584 40332 24636 40341
rect 45284 40400 45336 40452
rect 46940 40332 46992 40384
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 27950 40230 28002 40282
rect 28014 40230 28066 40282
rect 28078 40230 28130 40282
rect 28142 40230 28194 40282
rect 28206 40230 28258 40282
rect 37950 40230 38002 40282
rect 38014 40230 38066 40282
rect 38078 40230 38130 40282
rect 38142 40230 38194 40282
rect 38206 40230 38258 40282
rect 47950 40230 48002 40282
rect 48014 40230 48066 40282
rect 48078 40230 48130 40282
rect 48142 40230 48194 40282
rect 48206 40230 48258 40282
rect 8852 40128 8904 40180
rect 4344 40060 4396 40112
rect 8300 40060 8352 40112
rect 10140 40060 10192 40112
rect 11244 40128 11296 40180
rect 12072 40060 12124 40112
rect 12348 40128 12400 40180
rect 17408 40128 17460 40180
rect 17040 40060 17092 40112
rect 20720 40128 20772 40180
rect 18328 40060 18380 40112
rect 18512 40060 18564 40112
rect 8484 40035 8536 40044
rect 8484 40001 8493 40035
rect 8493 40001 8527 40035
rect 8527 40001 8536 40035
rect 8484 39992 8536 40001
rect 11704 40035 11756 40044
rect 11704 40001 11713 40035
rect 11713 40001 11747 40035
rect 11747 40001 11756 40035
rect 11704 39992 11756 40001
rect 2044 39967 2096 39976
rect 2044 39933 2053 39967
rect 2053 39933 2087 39967
rect 2087 39933 2096 39967
rect 2044 39924 2096 39933
rect 8392 39924 8444 39976
rect 10876 39924 10928 39976
rect 11520 39924 11572 39976
rect 11980 39967 12032 39976
rect 11980 39933 11989 39967
rect 11989 39933 12023 39967
rect 12023 39933 12032 39967
rect 11980 39924 12032 39933
rect 12440 39924 12492 39976
rect 13820 39992 13872 40044
rect 13912 39992 13964 40044
rect 13268 39924 13320 39976
rect 13636 39924 13688 39976
rect 19064 40060 19116 40112
rect 19156 40060 19208 40112
rect 3976 39856 4028 39908
rect 4068 39788 4120 39840
rect 11704 39788 11756 39840
rect 18328 39967 18380 39976
rect 18328 39933 18337 39967
rect 18337 39933 18371 39967
rect 18371 39933 18380 39967
rect 18328 39924 18380 39933
rect 18880 39924 18932 39976
rect 19984 40103 20036 40112
rect 19984 40069 19993 40103
rect 19993 40069 20027 40103
rect 20027 40069 20036 40103
rect 19984 40060 20036 40069
rect 19708 40035 19760 40044
rect 19708 40001 19717 40035
rect 19717 40001 19751 40035
rect 19751 40001 19760 40035
rect 19708 39992 19760 40001
rect 21272 40060 21324 40112
rect 21456 40060 21508 40112
rect 24768 40060 24820 40112
rect 23480 39992 23532 40044
rect 24676 40035 24728 40044
rect 24676 40001 24685 40035
rect 24685 40001 24719 40035
rect 24719 40001 24728 40035
rect 24676 39992 24728 40001
rect 21548 39924 21600 39976
rect 23848 39924 23900 39976
rect 15108 39831 15160 39840
rect 15108 39797 15117 39831
rect 15117 39797 15151 39831
rect 15151 39797 15160 39831
rect 15108 39788 15160 39797
rect 21456 39831 21508 39840
rect 21456 39797 21465 39831
rect 21465 39797 21499 39831
rect 21499 39797 21508 39831
rect 21456 39788 21508 39797
rect 21916 39788 21968 39840
rect 23572 39788 23624 39840
rect 23848 39831 23900 39840
rect 23848 39797 23857 39831
rect 23857 39797 23891 39831
rect 23891 39797 23900 39831
rect 23848 39788 23900 39797
rect 24308 39831 24360 39840
rect 24308 39797 24317 39831
rect 24317 39797 24351 39831
rect 24351 39797 24360 39831
rect 24308 39788 24360 39797
rect 38660 39788 38712 39840
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 32950 39686 33002 39738
rect 33014 39686 33066 39738
rect 33078 39686 33130 39738
rect 33142 39686 33194 39738
rect 33206 39686 33258 39738
rect 42950 39686 43002 39738
rect 43014 39686 43066 39738
rect 43078 39686 43130 39738
rect 43142 39686 43194 39738
rect 43206 39686 43258 39738
rect 7564 39584 7616 39636
rect 8208 39584 8260 39636
rect 9036 39584 9088 39636
rect 10784 39584 10836 39636
rect 12256 39584 12308 39636
rect 13360 39584 13412 39636
rect 14648 39584 14700 39636
rect 16488 39627 16540 39636
rect 16488 39593 16497 39627
rect 16497 39593 16531 39627
rect 16531 39593 16540 39627
rect 16488 39584 16540 39593
rect 16948 39627 17000 39636
rect 16948 39593 16957 39627
rect 16957 39593 16991 39627
rect 16991 39593 17000 39627
rect 16948 39584 17000 39593
rect 18420 39584 18472 39636
rect 1860 39516 1912 39568
rect 1308 39448 1360 39500
rect 2504 39448 2556 39500
rect 6552 39448 6604 39500
rect 8484 39448 8536 39500
rect 8668 39448 8720 39500
rect 4620 39380 4672 39432
rect 5448 39423 5500 39432
rect 5448 39389 5457 39423
rect 5457 39389 5491 39423
rect 5491 39389 5500 39423
rect 5448 39380 5500 39389
rect 8208 39380 8260 39432
rect 9036 39380 9088 39432
rect 11244 39491 11296 39500
rect 11244 39457 11253 39491
rect 11253 39457 11287 39491
rect 11287 39457 11296 39491
rect 11244 39448 11296 39457
rect 14740 39516 14792 39568
rect 17776 39516 17828 39568
rect 37832 39584 37884 39636
rect 11888 39380 11940 39432
rect 12256 39423 12308 39432
rect 12256 39389 12265 39423
rect 12265 39389 12299 39423
rect 12299 39389 12308 39423
rect 12256 39380 12308 39389
rect 12900 39380 12952 39432
rect 14004 39448 14056 39500
rect 15200 39448 15252 39500
rect 15568 39448 15620 39500
rect 17592 39491 17644 39500
rect 17592 39457 17601 39491
rect 17601 39457 17635 39491
rect 17635 39457 17644 39491
rect 17592 39448 17644 39457
rect 19800 39516 19852 39568
rect 21732 39516 21784 39568
rect 19708 39448 19760 39500
rect 21916 39448 21968 39500
rect 22100 39491 22152 39500
rect 22100 39457 22109 39491
rect 22109 39457 22143 39491
rect 22143 39457 22152 39491
rect 22100 39448 22152 39457
rect 22744 39491 22796 39500
rect 22744 39457 22753 39491
rect 22753 39457 22787 39491
rect 22787 39457 22796 39491
rect 22744 39448 22796 39457
rect 23296 39448 23348 39500
rect 5816 39244 5868 39296
rect 8668 39312 8720 39364
rect 12072 39312 12124 39364
rect 19984 39380 20036 39432
rect 24308 39380 24360 39432
rect 20352 39312 20404 39364
rect 21272 39312 21324 39364
rect 24584 39312 24636 39364
rect 8576 39244 8628 39296
rect 9128 39287 9180 39296
rect 9128 39253 9137 39287
rect 9137 39253 9171 39287
rect 9171 39253 9180 39287
rect 9128 39244 9180 39253
rect 9496 39287 9548 39296
rect 9496 39253 9505 39287
rect 9505 39253 9539 39287
rect 9539 39253 9548 39287
rect 9496 39244 9548 39253
rect 12624 39244 12676 39296
rect 14188 39244 14240 39296
rect 14464 39244 14516 39296
rect 15200 39287 15252 39296
rect 15200 39253 15209 39287
rect 15209 39253 15243 39287
rect 15243 39253 15252 39287
rect 15200 39244 15252 39253
rect 15292 39287 15344 39296
rect 15292 39253 15301 39287
rect 15301 39253 15335 39287
rect 15335 39253 15344 39287
rect 15292 39244 15344 39253
rect 17224 39244 17276 39296
rect 18420 39244 18472 39296
rect 21640 39244 21692 39296
rect 22192 39287 22244 39296
rect 22192 39253 22201 39287
rect 22201 39253 22235 39287
rect 22235 39253 22244 39287
rect 22192 39244 22244 39253
rect 23572 39287 23624 39296
rect 23572 39253 23581 39287
rect 23581 39253 23615 39287
rect 23615 39253 23624 39287
rect 23572 39244 23624 39253
rect 23756 39244 23808 39296
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 27950 39142 28002 39194
rect 28014 39142 28066 39194
rect 28078 39142 28130 39194
rect 28142 39142 28194 39194
rect 28206 39142 28258 39194
rect 37950 39142 38002 39194
rect 38014 39142 38066 39194
rect 38078 39142 38130 39194
rect 38142 39142 38194 39194
rect 38206 39142 38258 39194
rect 47950 39142 48002 39194
rect 48014 39142 48066 39194
rect 48078 39142 48130 39194
rect 48142 39142 48194 39194
rect 48206 39142 48258 39194
rect 5724 39040 5776 39092
rect 7288 38972 7340 39024
rect 8208 38972 8260 39024
rect 10140 39040 10192 39092
rect 12532 39040 12584 39092
rect 13176 39040 13228 39092
rect 11704 38972 11756 39024
rect 12716 38972 12768 39024
rect 14188 39083 14240 39092
rect 14188 39049 14197 39083
rect 14197 39049 14231 39083
rect 14231 39049 14240 39083
rect 14188 39040 14240 39049
rect 15016 39040 15068 39092
rect 16948 39040 17000 39092
rect 17776 39040 17828 39092
rect 19984 39040 20036 39092
rect 5264 38904 5316 38956
rect 8484 38947 8536 38956
rect 8484 38913 8493 38947
rect 8493 38913 8527 38947
rect 8527 38913 8536 38947
rect 8484 38904 8536 38913
rect 12532 38947 12584 38956
rect 12532 38913 12541 38947
rect 12541 38913 12575 38947
rect 12575 38913 12584 38947
rect 12532 38904 12584 38913
rect 13084 38904 13136 38956
rect 14004 38947 14056 38956
rect 14004 38913 14013 38947
rect 14013 38913 14047 38947
rect 14047 38913 14056 38947
rect 14004 38904 14056 38913
rect 15476 38904 15528 38956
rect 16028 38904 16080 38956
rect 21272 38972 21324 39024
rect 16856 38904 16908 38956
rect 18236 38904 18288 38956
rect 4988 38836 5040 38888
rect 6460 38836 6512 38888
rect 7196 38836 7248 38888
rect 9128 38836 9180 38888
rect 11888 38836 11940 38888
rect 12992 38836 13044 38888
rect 13452 38879 13504 38888
rect 13452 38845 13461 38879
rect 13461 38845 13495 38879
rect 13495 38845 13504 38879
rect 13452 38836 13504 38845
rect 13636 38879 13688 38888
rect 13636 38845 13645 38879
rect 13645 38845 13679 38879
rect 13679 38845 13688 38879
rect 13636 38836 13688 38845
rect 14740 38879 14792 38888
rect 14740 38845 14749 38879
rect 14749 38845 14783 38879
rect 14783 38845 14792 38879
rect 14740 38836 14792 38845
rect 5632 38768 5684 38820
rect 8484 38768 8536 38820
rect 11152 38811 11204 38820
rect 11152 38777 11161 38811
rect 11161 38777 11195 38811
rect 11195 38777 11204 38811
rect 11152 38768 11204 38777
rect 5356 38700 5408 38752
rect 6092 38700 6144 38752
rect 8944 38700 8996 38752
rect 9772 38700 9824 38752
rect 11244 38700 11296 38752
rect 14280 38768 14332 38820
rect 14004 38700 14056 38752
rect 15660 38700 15712 38752
rect 18696 38836 18748 38888
rect 19248 38836 19300 38888
rect 19892 38836 19944 38888
rect 20168 38836 20220 38888
rect 23848 39083 23900 39092
rect 23848 39049 23857 39083
rect 23857 39049 23891 39083
rect 23891 39049 23900 39083
rect 23848 39040 23900 39049
rect 23480 38904 23532 38956
rect 22560 38836 22612 38888
rect 23296 38836 23348 38888
rect 48872 38836 48924 38888
rect 21640 38768 21692 38820
rect 18420 38700 18472 38752
rect 19156 38700 19208 38752
rect 19248 38700 19300 38752
rect 22100 38700 22152 38752
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 32950 38598 33002 38650
rect 33014 38598 33066 38650
rect 33078 38598 33130 38650
rect 33142 38598 33194 38650
rect 33206 38598 33258 38650
rect 42950 38598 43002 38650
rect 43014 38598 43066 38650
rect 43078 38598 43130 38650
rect 43142 38598 43194 38650
rect 43206 38598 43258 38650
rect 4620 38539 4672 38548
rect 4620 38505 4629 38539
rect 4629 38505 4663 38539
rect 4663 38505 4672 38539
rect 4620 38496 4672 38505
rect 5264 38539 5316 38548
rect 5264 38505 5273 38539
rect 5273 38505 5307 38539
rect 5307 38505 5316 38539
rect 5264 38496 5316 38505
rect 5724 38496 5776 38548
rect 6920 38496 6972 38548
rect 9496 38496 9548 38548
rect 11980 38496 12032 38548
rect 8300 38428 8352 38480
rect 9312 38428 9364 38480
rect 1308 38360 1360 38412
rect 5540 38360 5592 38412
rect 6736 38360 6788 38412
rect 8852 38360 8904 38412
rect 9404 38360 9456 38412
rect 9496 38360 9548 38412
rect 9772 38403 9824 38412
rect 9772 38369 9781 38403
rect 9781 38369 9815 38403
rect 9815 38369 9824 38403
rect 9772 38360 9824 38369
rect 10968 38403 11020 38412
rect 10968 38369 10977 38403
rect 10977 38369 11011 38403
rect 11011 38369 11020 38403
rect 10968 38360 11020 38369
rect 15108 38496 15160 38548
rect 19064 38496 19116 38548
rect 22744 38496 22796 38548
rect 17868 38428 17920 38480
rect 5908 38292 5960 38344
rect 6828 38335 6880 38344
rect 6828 38301 6837 38335
rect 6837 38301 6871 38335
rect 6871 38301 6880 38335
rect 6828 38292 6880 38301
rect 8208 38292 8260 38344
rect 8392 38292 8444 38344
rect 14556 38360 14608 38412
rect 16488 38403 16540 38412
rect 16488 38369 16497 38403
rect 16497 38369 16531 38403
rect 16531 38369 16540 38403
rect 16488 38360 16540 38369
rect 18328 38360 18380 38412
rect 21456 38360 21508 38412
rect 23940 38360 23992 38412
rect 11980 38335 12032 38344
rect 11980 38301 11989 38335
rect 11989 38301 12023 38335
rect 12023 38301 12032 38335
rect 11980 38292 12032 38301
rect 14280 38335 14332 38344
rect 14280 38301 14289 38335
rect 14289 38301 14323 38335
rect 14323 38301 14332 38335
rect 14280 38292 14332 38301
rect 20536 38335 20588 38344
rect 20536 38301 20545 38335
rect 20545 38301 20579 38335
rect 20579 38301 20588 38335
rect 20536 38292 20588 38301
rect 22836 38292 22888 38344
rect 23572 38335 23624 38344
rect 23572 38301 23581 38335
rect 23581 38301 23615 38335
rect 23615 38301 23624 38335
rect 23572 38292 23624 38301
rect 24400 38292 24452 38344
rect 7380 38224 7432 38276
rect 5448 38156 5500 38208
rect 6644 38156 6696 38208
rect 9864 38224 9916 38276
rect 9956 38224 10008 38276
rect 8852 38156 8904 38208
rect 9772 38156 9824 38208
rect 10876 38199 10928 38208
rect 10876 38165 10885 38199
rect 10885 38165 10919 38199
rect 10919 38165 10928 38199
rect 10876 38156 10928 38165
rect 11060 38156 11112 38208
rect 12532 38156 12584 38208
rect 12716 38224 12768 38276
rect 14832 38224 14884 38276
rect 13084 38156 13136 38208
rect 14464 38156 14516 38208
rect 16672 38224 16724 38276
rect 17224 38224 17276 38276
rect 15568 38156 15620 38208
rect 16120 38156 16172 38208
rect 21272 38224 21324 38276
rect 22284 38156 22336 38208
rect 22376 38156 22428 38208
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 27950 38054 28002 38106
rect 28014 38054 28066 38106
rect 28078 38054 28130 38106
rect 28142 38054 28194 38106
rect 28206 38054 28258 38106
rect 37950 38054 38002 38106
rect 38014 38054 38066 38106
rect 38078 38054 38130 38106
rect 38142 38054 38194 38106
rect 38206 38054 38258 38106
rect 47950 38054 48002 38106
rect 48014 38054 48066 38106
rect 48078 38054 48130 38106
rect 48142 38054 48194 38106
rect 48206 38054 48258 38106
rect 4344 37995 4396 38004
rect 4344 37961 4353 37995
rect 4353 37961 4387 37995
rect 4387 37961 4396 37995
rect 4344 37952 4396 37961
rect 5908 37952 5960 38004
rect 5724 37884 5776 37936
rect 7288 37952 7340 38004
rect 7472 37952 7524 38004
rect 8576 37995 8628 38004
rect 8576 37961 8585 37995
rect 8585 37961 8619 37995
rect 8619 37961 8628 37995
rect 8576 37952 8628 37961
rect 8944 37952 8996 38004
rect 9588 37995 9640 38004
rect 9588 37961 9597 37995
rect 9597 37961 9631 37995
rect 9631 37961 9640 37995
rect 9588 37952 9640 37961
rect 9864 37952 9916 38004
rect 11612 37952 11664 38004
rect 12164 37952 12216 38004
rect 12716 37952 12768 38004
rect 14464 37952 14516 38004
rect 8208 37816 8260 37868
rect 8392 37816 8444 37868
rect 1308 37748 1360 37800
rect 4528 37748 4580 37800
rect 4896 37748 4948 37800
rect 5448 37748 5500 37800
rect 5908 37791 5960 37800
rect 5908 37757 5917 37791
rect 5917 37757 5951 37791
rect 5951 37757 5960 37791
rect 5908 37748 5960 37757
rect 6828 37791 6880 37800
rect 6828 37757 6837 37791
rect 6837 37757 6871 37791
rect 6871 37757 6880 37791
rect 6828 37748 6880 37757
rect 8300 37748 8352 37800
rect 9864 37791 9916 37800
rect 9864 37757 9873 37791
rect 9873 37757 9907 37791
rect 9907 37757 9916 37791
rect 10968 37884 11020 37936
rect 13820 37927 13872 37936
rect 13820 37893 13829 37927
rect 13829 37893 13863 37927
rect 13863 37893 13872 37927
rect 13820 37884 13872 37893
rect 17868 37952 17920 38004
rect 22284 37952 22336 38004
rect 23388 37952 23440 38004
rect 15384 37884 15436 37936
rect 17224 37884 17276 37936
rect 18604 37884 18656 37936
rect 18788 37884 18840 37936
rect 20720 37884 20772 37936
rect 22008 37884 22060 37936
rect 12624 37816 12676 37868
rect 14556 37859 14608 37868
rect 14556 37825 14565 37859
rect 14565 37825 14599 37859
rect 14599 37825 14608 37859
rect 14556 37816 14608 37825
rect 16488 37816 16540 37868
rect 9864 37748 9916 37757
rect 10140 37748 10192 37800
rect 8116 37680 8168 37732
rect 9496 37680 9548 37732
rect 12992 37791 13044 37800
rect 12992 37757 13001 37791
rect 13001 37757 13035 37791
rect 13035 37757 13044 37791
rect 12992 37748 13044 37757
rect 13084 37791 13136 37800
rect 13084 37757 13093 37791
rect 13093 37757 13127 37791
rect 13127 37757 13136 37791
rect 13084 37748 13136 37757
rect 13728 37748 13780 37800
rect 14096 37748 14148 37800
rect 15200 37748 15252 37800
rect 16120 37748 16172 37800
rect 17592 37748 17644 37800
rect 18788 37748 18840 37800
rect 20168 37748 20220 37800
rect 20536 37748 20588 37800
rect 23296 37791 23348 37800
rect 23296 37757 23305 37791
rect 23305 37757 23339 37791
rect 23339 37757 23348 37791
rect 23296 37748 23348 37757
rect 14556 37680 14608 37732
rect 8392 37612 8444 37664
rect 9220 37655 9272 37664
rect 9220 37621 9229 37655
rect 9229 37621 9263 37655
rect 9263 37621 9272 37655
rect 9220 37612 9272 37621
rect 14832 37612 14884 37664
rect 16672 37612 16724 37664
rect 21364 37612 21416 37664
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 32950 37510 33002 37562
rect 33014 37510 33066 37562
rect 33078 37510 33130 37562
rect 33142 37510 33194 37562
rect 33206 37510 33258 37562
rect 42950 37510 43002 37562
rect 43014 37510 43066 37562
rect 43078 37510 43130 37562
rect 43142 37510 43194 37562
rect 43206 37510 43258 37562
rect 5908 37408 5960 37460
rect 5632 37315 5684 37324
rect 5632 37281 5641 37315
rect 5641 37281 5675 37315
rect 5675 37281 5684 37315
rect 5632 37272 5684 37281
rect 8024 37340 8076 37392
rect 6644 37272 6696 37324
rect 7380 37272 7432 37324
rect 8300 37408 8352 37460
rect 11060 37408 11112 37460
rect 13728 37451 13780 37460
rect 13728 37417 13737 37451
rect 13737 37417 13771 37451
rect 13771 37417 13780 37451
rect 13728 37408 13780 37417
rect 18788 37451 18840 37460
rect 18788 37417 18797 37451
rect 18797 37417 18831 37451
rect 18831 37417 18840 37451
rect 18788 37408 18840 37417
rect 22284 37451 22336 37460
rect 22284 37417 22293 37451
rect 22293 37417 22327 37451
rect 22327 37417 22336 37451
rect 22284 37408 22336 37417
rect 23940 37408 23992 37460
rect 7656 37204 7708 37256
rect 9864 37340 9916 37392
rect 10232 37340 10284 37392
rect 9680 37272 9732 37324
rect 13544 37272 13596 37324
rect 14280 37272 14332 37324
rect 15568 37272 15620 37324
rect 16120 37272 16172 37324
rect 18880 37272 18932 37324
rect 21456 37272 21508 37324
rect 23296 37315 23348 37324
rect 23296 37281 23305 37315
rect 23305 37281 23339 37315
rect 23339 37281 23348 37315
rect 23296 37272 23348 37281
rect 8668 37204 8720 37256
rect 9036 37204 9088 37256
rect 11060 37247 11112 37256
rect 11060 37213 11069 37247
rect 11069 37213 11103 37247
rect 11103 37213 11112 37247
rect 11060 37204 11112 37213
rect 11980 37247 12032 37256
rect 11980 37213 11989 37247
rect 11989 37213 12023 37247
rect 12023 37213 12032 37247
rect 11980 37204 12032 37213
rect 5540 37111 5592 37120
rect 5540 37077 5549 37111
rect 5549 37077 5583 37111
rect 5583 37077 5592 37111
rect 5540 37068 5592 37077
rect 7196 37136 7248 37188
rect 7472 37136 7524 37188
rect 6736 37111 6788 37120
rect 6736 37077 6745 37111
rect 6745 37077 6779 37111
rect 6779 37077 6788 37111
rect 6736 37068 6788 37077
rect 7564 37111 7616 37120
rect 7564 37077 7573 37111
rect 7573 37077 7607 37111
rect 7607 37077 7616 37111
rect 7564 37068 7616 37077
rect 7840 37136 7892 37188
rect 9496 37136 9548 37188
rect 12716 37136 12768 37188
rect 14464 37136 14516 37188
rect 15384 37136 15436 37188
rect 8208 37068 8260 37120
rect 10416 37068 10468 37120
rect 15936 37068 15988 37120
rect 18696 37204 18748 37256
rect 20168 37204 20220 37256
rect 22836 37204 22888 37256
rect 23572 37204 23624 37256
rect 17224 37136 17276 37188
rect 17408 37136 17460 37188
rect 17776 37136 17828 37188
rect 18788 37136 18840 37188
rect 20812 37179 20864 37188
rect 20812 37145 20821 37179
rect 20821 37145 20855 37179
rect 20855 37145 20864 37179
rect 20812 37136 20864 37145
rect 18696 37068 18748 37120
rect 20720 37068 20772 37120
rect 21272 37136 21324 37188
rect 21180 37068 21232 37120
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 27950 36966 28002 37018
rect 28014 36966 28066 37018
rect 28078 36966 28130 37018
rect 28142 36966 28194 37018
rect 28206 36966 28258 37018
rect 37950 36966 38002 37018
rect 38014 36966 38066 37018
rect 38078 36966 38130 37018
rect 38142 36966 38194 37018
rect 38206 36966 38258 37018
rect 47950 36966 48002 37018
rect 48014 36966 48066 37018
rect 48078 36966 48130 37018
rect 48142 36966 48194 37018
rect 48206 36966 48258 37018
rect 6184 36864 6236 36916
rect 7104 36864 7156 36916
rect 7380 36864 7432 36916
rect 7656 36864 7708 36916
rect 8392 36907 8444 36916
rect 8392 36873 8401 36907
rect 8401 36873 8435 36907
rect 8435 36873 8444 36907
rect 8392 36864 8444 36873
rect 9220 36864 9272 36916
rect 9588 36907 9640 36916
rect 9588 36873 9597 36907
rect 9597 36873 9631 36907
rect 9631 36873 9640 36907
rect 9588 36864 9640 36873
rect 10600 36864 10652 36916
rect 5080 36796 5132 36848
rect 6736 36796 6788 36848
rect 8944 36796 8996 36848
rect 1768 36771 1820 36780
rect 1768 36737 1777 36771
rect 1777 36737 1811 36771
rect 1811 36737 1820 36771
rect 1768 36728 1820 36737
rect 6828 36728 6880 36780
rect 1308 36660 1360 36712
rect 3516 36660 3568 36712
rect 6552 36660 6604 36712
rect 7104 36703 7156 36712
rect 7104 36669 7113 36703
rect 7113 36669 7147 36703
rect 7147 36669 7156 36703
rect 7104 36660 7156 36669
rect 7380 36728 7432 36780
rect 11796 36728 11848 36780
rect 7656 36660 7708 36712
rect 8668 36703 8720 36712
rect 8668 36669 8677 36703
rect 8677 36669 8711 36703
rect 8711 36669 8720 36703
rect 8668 36660 8720 36669
rect 9128 36660 9180 36712
rect 9588 36660 9640 36712
rect 10600 36660 10652 36712
rect 11336 36660 11388 36712
rect 3424 36592 3476 36644
rect 7472 36592 7524 36644
rect 9864 36592 9916 36644
rect 9956 36592 10008 36644
rect 12624 36864 12676 36916
rect 15108 36864 15160 36916
rect 15476 36907 15528 36916
rect 15476 36873 15485 36907
rect 15485 36873 15519 36907
rect 15519 36873 15528 36907
rect 15476 36864 15528 36873
rect 16396 36864 16448 36916
rect 16580 36864 16632 36916
rect 22376 36907 22428 36916
rect 22376 36873 22385 36907
rect 22385 36873 22419 36907
rect 22419 36873 22428 36907
rect 22376 36864 22428 36873
rect 22652 36864 22704 36916
rect 12072 36796 12124 36848
rect 14280 36796 14332 36848
rect 12348 36728 12400 36780
rect 13820 36728 13872 36780
rect 18052 36796 18104 36848
rect 18880 36796 18932 36848
rect 19340 36796 19392 36848
rect 20720 36796 20772 36848
rect 15200 36728 15252 36780
rect 16856 36771 16908 36780
rect 16856 36737 16865 36771
rect 16865 36737 16899 36771
rect 16899 36737 16908 36771
rect 16856 36728 16908 36737
rect 16948 36728 17000 36780
rect 18604 36728 18656 36780
rect 18696 36728 18748 36780
rect 14832 36703 14884 36712
rect 14832 36669 14841 36703
rect 14841 36669 14875 36703
rect 14875 36669 14884 36703
rect 14832 36660 14884 36669
rect 16028 36703 16080 36712
rect 16028 36669 16037 36703
rect 16037 36669 16071 36703
rect 16071 36669 16080 36703
rect 16028 36660 16080 36669
rect 17408 36703 17460 36712
rect 17408 36669 17417 36703
rect 17417 36669 17451 36703
rect 17451 36669 17460 36703
rect 17408 36660 17460 36669
rect 15292 36592 15344 36644
rect 18788 36660 18840 36712
rect 18880 36660 18932 36712
rect 23572 36728 23624 36780
rect 4712 36567 4764 36576
rect 4712 36533 4721 36567
rect 4721 36533 4755 36567
rect 4755 36533 4764 36567
rect 4712 36524 4764 36533
rect 5816 36524 5868 36576
rect 7932 36524 7984 36576
rect 8300 36524 8352 36576
rect 11336 36524 11388 36576
rect 17684 36524 17736 36576
rect 17776 36567 17828 36576
rect 17776 36533 17785 36567
rect 17785 36533 17819 36567
rect 17819 36533 17828 36567
rect 17776 36524 17828 36533
rect 18052 36524 18104 36576
rect 18972 36524 19024 36576
rect 21548 36592 21600 36644
rect 20812 36524 20864 36576
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 32950 36422 33002 36474
rect 33014 36422 33066 36474
rect 33078 36422 33130 36474
rect 33142 36422 33194 36474
rect 33206 36422 33258 36474
rect 42950 36422 43002 36474
rect 43014 36422 43066 36474
rect 43078 36422 43130 36474
rect 43142 36422 43194 36474
rect 43206 36422 43258 36474
rect 5540 36320 5592 36372
rect 6552 36252 6604 36304
rect 10600 36320 10652 36372
rect 11796 36363 11848 36372
rect 11796 36329 11805 36363
rect 11805 36329 11839 36363
rect 11839 36329 11848 36363
rect 11796 36320 11848 36329
rect 12808 36320 12860 36372
rect 14740 36320 14792 36372
rect 17408 36320 17460 36372
rect 22192 36320 22244 36372
rect 19064 36252 19116 36304
rect 19340 36252 19392 36304
rect 21916 36295 21968 36304
rect 21916 36261 21925 36295
rect 21925 36261 21959 36295
rect 21959 36261 21968 36295
rect 21916 36252 21968 36261
rect 6460 36184 6512 36236
rect 7104 36184 7156 36236
rect 7932 36184 7984 36236
rect 8484 36227 8536 36236
rect 8484 36193 8493 36227
rect 8493 36193 8527 36227
rect 8527 36193 8536 36227
rect 8484 36184 8536 36193
rect 8944 36184 8996 36236
rect 4068 36116 4120 36168
rect 6368 36116 6420 36168
rect 6644 36116 6696 36168
rect 6920 36116 6972 36168
rect 9036 36116 9088 36168
rect 13728 36184 13780 36236
rect 16028 36184 16080 36236
rect 16856 36184 16908 36236
rect 20168 36227 20220 36236
rect 20168 36193 20177 36227
rect 20177 36193 20211 36227
rect 20211 36193 20220 36227
rect 20168 36184 20220 36193
rect 13912 36116 13964 36168
rect 14280 36116 14332 36168
rect 18420 36116 18472 36168
rect 2780 36091 2832 36100
rect 2780 36057 2789 36091
rect 2789 36057 2823 36091
rect 2823 36057 2832 36091
rect 2780 36048 2832 36057
rect 6276 36048 6328 36100
rect 6460 36048 6512 36100
rect 7012 36091 7064 36100
rect 7012 36057 7021 36091
rect 7021 36057 7055 36091
rect 7055 36057 7064 36091
rect 7012 36048 7064 36057
rect 7380 36048 7432 36100
rect 7656 36048 7708 36100
rect 10416 36048 10468 36100
rect 11244 36048 11296 36100
rect 5724 35980 5776 36032
rect 6828 35980 6880 36032
rect 7932 35980 7984 36032
rect 12808 36023 12860 36032
rect 12808 35989 12817 36023
rect 12817 35989 12851 36023
rect 12851 35989 12860 36023
rect 12808 35980 12860 35989
rect 13360 35980 13412 36032
rect 15384 36048 15436 36100
rect 16212 35980 16264 36032
rect 20444 36091 20496 36100
rect 20444 36057 20453 36091
rect 20453 36057 20487 36091
rect 20487 36057 20496 36091
rect 20444 36048 20496 36057
rect 20720 36048 20772 36100
rect 23388 36048 23440 36100
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 27950 35878 28002 35930
rect 28014 35878 28066 35930
rect 28078 35878 28130 35930
rect 28142 35878 28194 35930
rect 28206 35878 28258 35930
rect 37950 35878 38002 35930
rect 38014 35878 38066 35930
rect 38078 35878 38130 35930
rect 38142 35878 38194 35930
rect 38206 35878 38258 35930
rect 47950 35878 48002 35930
rect 48014 35878 48066 35930
rect 48078 35878 48130 35930
rect 48142 35878 48194 35930
rect 48206 35878 48258 35930
rect 5724 35776 5776 35828
rect 7748 35776 7800 35828
rect 6000 35708 6052 35760
rect 5356 35640 5408 35692
rect 4804 35504 4856 35556
rect 6552 35572 6604 35624
rect 8484 35708 8536 35760
rect 9772 35776 9824 35828
rect 10048 35776 10100 35828
rect 13544 35776 13596 35828
rect 16580 35776 16632 35828
rect 17776 35776 17828 35828
rect 10140 35708 10192 35760
rect 11520 35708 11572 35760
rect 12716 35708 12768 35760
rect 14464 35708 14516 35760
rect 7564 35640 7616 35692
rect 14096 35640 14148 35692
rect 19432 35776 19484 35828
rect 22284 35776 22336 35828
rect 7472 35615 7524 35624
rect 7472 35581 7481 35615
rect 7481 35581 7515 35615
rect 7515 35581 7524 35615
rect 7472 35572 7524 35581
rect 8576 35615 8628 35624
rect 8576 35581 8585 35615
rect 8585 35581 8619 35615
rect 8619 35581 8628 35615
rect 8576 35572 8628 35581
rect 8668 35572 8720 35624
rect 10508 35572 10560 35624
rect 12348 35572 12400 35624
rect 11244 35504 11296 35556
rect 6736 35436 6788 35488
rect 9128 35436 9180 35488
rect 9220 35479 9272 35488
rect 9220 35445 9229 35479
rect 9229 35445 9263 35479
rect 9263 35445 9272 35479
rect 9220 35436 9272 35445
rect 13544 35572 13596 35624
rect 14648 35572 14700 35624
rect 17408 35572 17460 35624
rect 17776 35572 17828 35624
rect 17868 35572 17920 35624
rect 15844 35504 15896 35556
rect 17040 35504 17092 35556
rect 20720 35708 20772 35760
rect 22008 35751 22060 35760
rect 22008 35717 22017 35751
rect 22017 35717 22051 35751
rect 22051 35717 22060 35751
rect 22008 35708 22060 35717
rect 19340 35504 19392 35556
rect 24124 35572 24176 35624
rect 14280 35436 14332 35488
rect 17316 35436 17368 35488
rect 18420 35436 18472 35488
rect 19708 35436 19760 35488
rect 21548 35436 21600 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 32950 35334 33002 35386
rect 33014 35334 33066 35386
rect 33078 35334 33130 35386
rect 33142 35334 33194 35386
rect 33206 35334 33258 35386
rect 42950 35334 43002 35386
rect 43014 35334 43066 35386
rect 43078 35334 43130 35386
rect 43142 35334 43194 35386
rect 43206 35334 43258 35386
rect 7840 35275 7892 35284
rect 7840 35241 7849 35275
rect 7849 35241 7883 35275
rect 7883 35241 7892 35275
rect 7840 35232 7892 35241
rect 10508 35232 10560 35284
rect 12808 35232 12860 35284
rect 13452 35232 13504 35284
rect 16304 35232 16356 35284
rect 17408 35232 17460 35284
rect 7656 35164 7708 35216
rect 8208 35164 8260 35216
rect 9312 35164 9364 35216
rect 10968 35164 11020 35216
rect 17040 35164 17092 35216
rect 19340 35164 19392 35216
rect 23756 35164 23808 35216
rect 1308 35096 1360 35148
rect 5908 35139 5960 35148
rect 5908 35105 5917 35139
rect 5917 35105 5951 35139
rect 5951 35105 5960 35139
rect 5908 35096 5960 35105
rect 3976 35028 4028 35080
rect 5816 35071 5868 35080
rect 5816 35037 5825 35071
rect 5825 35037 5859 35071
rect 5859 35037 5868 35071
rect 5816 35028 5868 35037
rect 6736 35096 6788 35148
rect 7196 35139 7248 35148
rect 7196 35105 7205 35139
rect 7205 35105 7239 35139
rect 7239 35105 7248 35139
rect 7196 35096 7248 35105
rect 7748 35096 7800 35148
rect 12072 35096 12124 35148
rect 13544 35139 13596 35148
rect 13544 35105 13553 35139
rect 13553 35105 13587 35139
rect 13587 35105 13596 35139
rect 13544 35096 13596 35105
rect 14924 35139 14976 35148
rect 14924 35105 14933 35139
rect 14933 35105 14967 35139
rect 14967 35105 14976 35139
rect 14924 35096 14976 35105
rect 16672 35096 16724 35148
rect 19708 35096 19760 35148
rect 20628 35139 20680 35148
rect 20628 35105 20637 35139
rect 20637 35105 20671 35139
rect 20671 35105 20680 35139
rect 20628 35096 20680 35105
rect 21732 35139 21784 35148
rect 21732 35105 21741 35139
rect 21741 35105 21775 35139
rect 21775 35105 21784 35139
rect 21732 35096 21784 35105
rect 21824 35139 21876 35148
rect 21824 35105 21833 35139
rect 21833 35105 21867 35139
rect 21867 35105 21876 35139
rect 21824 35096 21876 35105
rect 8300 35028 8352 35080
rect 13360 35071 13412 35080
rect 13360 35037 13369 35071
rect 13369 35037 13403 35071
rect 13403 35037 13412 35071
rect 13360 35028 13412 35037
rect 14648 35028 14700 35080
rect 16212 35028 16264 35080
rect 21180 35028 21232 35080
rect 21640 35071 21692 35080
rect 21640 35037 21649 35071
rect 21649 35037 21683 35071
rect 21683 35037 21692 35071
rect 21640 35028 21692 35037
rect 7196 34960 7248 35012
rect 8116 34960 8168 35012
rect 6920 34892 6972 34944
rect 7012 34892 7064 34944
rect 8208 34935 8260 34944
rect 8208 34901 8217 34935
rect 8217 34901 8251 34935
rect 8251 34901 8260 34935
rect 8208 34892 8260 34901
rect 10232 34960 10284 35012
rect 10416 34960 10468 35012
rect 12808 34960 12860 35012
rect 8392 34892 8444 34944
rect 9680 34892 9732 34944
rect 15936 34935 15988 34944
rect 15936 34901 15945 34935
rect 15945 34901 15979 34935
rect 15979 34901 15988 34935
rect 15936 34892 15988 34901
rect 16212 34892 16264 34944
rect 17316 34960 17368 35012
rect 17868 34960 17920 35012
rect 21364 34960 21416 35012
rect 17500 34892 17552 34944
rect 18328 34892 18380 34944
rect 21272 34935 21324 34944
rect 21272 34901 21281 34935
rect 21281 34901 21315 34935
rect 21315 34901 21324 34935
rect 21272 34892 21324 34901
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 27950 34790 28002 34842
rect 28014 34790 28066 34842
rect 28078 34790 28130 34842
rect 28142 34790 28194 34842
rect 28206 34790 28258 34842
rect 37950 34790 38002 34842
rect 38014 34790 38066 34842
rect 38078 34790 38130 34842
rect 38142 34790 38194 34842
rect 38206 34790 38258 34842
rect 47950 34790 48002 34842
rect 48014 34790 48066 34842
rect 48078 34790 48130 34842
rect 48142 34790 48194 34842
rect 48206 34790 48258 34842
rect 8392 34688 8444 34740
rect 8760 34731 8812 34740
rect 8760 34697 8769 34731
rect 8769 34697 8803 34731
rect 8803 34697 8812 34731
rect 8760 34688 8812 34697
rect 10968 34688 11020 34740
rect 6644 34620 6696 34672
rect 12348 34663 12400 34672
rect 12348 34629 12357 34663
rect 12357 34629 12391 34663
rect 12391 34629 12400 34663
rect 12348 34620 12400 34629
rect 12624 34620 12676 34672
rect 14004 34620 14056 34672
rect 7288 34552 7340 34604
rect 2044 34527 2096 34536
rect 2044 34493 2053 34527
rect 2053 34493 2087 34527
rect 2087 34493 2096 34527
rect 2044 34484 2096 34493
rect 8668 34552 8720 34604
rect 9956 34552 10008 34604
rect 11888 34552 11940 34604
rect 12072 34595 12124 34604
rect 12072 34561 12081 34595
rect 12081 34561 12115 34595
rect 12115 34561 12124 34595
rect 12072 34552 12124 34561
rect 13636 34552 13688 34604
rect 16120 34688 16172 34740
rect 17500 34688 17552 34740
rect 21824 34688 21876 34740
rect 15384 34620 15436 34672
rect 16212 34620 16264 34672
rect 17224 34620 17276 34672
rect 17408 34620 17460 34672
rect 17960 34620 18012 34672
rect 20720 34620 20772 34672
rect 19708 34595 19760 34604
rect 19708 34561 19717 34595
rect 19717 34561 19751 34595
rect 19751 34561 19760 34595
rect 19708 34552 19760 34561
rect 7288 34416 7340 34468
rect 7104 34348 7156 34400
rect 8208 34416 8260 34468
rect 10232 34484 10284 34536
rect 10508 34527 10560 34536
rect 10508 34493 10517 34527
rect 10517 34493 10551 34527
rect 10551 34493 10560 34527
rect 10508 34484 10560 34493
rect 13544 34484 13596 34536
rect 14280 34484 14332 34536
rect 14832 34527 14884 34536
rect 14832 34493 14841 34527
rect 14841 34493 14875 34527
rect 14875 34493 14884 34527
rect 14832 34484 14884 34493
rect 16672 34484 16724 34536
rect 9404 34416 9456 34468
rect 14004 34416 14056 34468
rect 14372 34416 14424 34468
rect 17316 34416 17368 34468
rect 21548 34484 21600 34536
rect 7564 34391 7616 34400
rect 7564 34357 7573 34391
rect 7573 34357 7607 34391
rect 7607 34357 7616 34391
rect 7564 34348 7616 34357
rect 9956 34391 10008 34400
rect 9956 34357 9965 34391
rect 9965 34357 9999 34391
rect 9999 34357 10008 34391
rect 9956 34348 10008 34357
rect 10048 34348 10100 34400
rect 12072 34348 12124 34400
rect 12164 34348 12216 34400
rect 15200 34348 15252 34400
rect 16488 34348 16540 34400
rect 18788 34348 18840 34400
rect 22560 34416 22612 34468
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 32950 34246 33002 34298
rect 33014 34246 33066 34298
rect 33078 34246 33130 34298
rect 33142 34246 33194 34298
rect 33206 34246 33258 34298
rect 42950 34246 43002 34298
rect 43014 34246 43066 34298
rect 43078 34246 43130 34298
rect 43142 34246 43194 34298
rect 43206 34246 43258 34298
rect 7196 34144 7248 34196
rect 7840 34144 7892 34196
rect 10324 34144 10376 34196
rect 7748 34076 7800 34128
rect 9036 34008 9088 34060
rect 12072 34144 12124 34196
rect 11060 33940 11112 33992
rect 11428 33940 11480 33992
rect 12440 34008 12492 34060
rect 12992 34008 13044 34060
rect 13912 34144 13964 34196
rect 15936 34144 15988 34196
rect 21456 34144 21508 34196
rect 14648 34008 14700 34060
rect 19064 34008 19116 34060
rect 13544 33940 13596 33992
rect 14280 33983 14332 33992
rect 14280 33949 14289 33983
rect 14289 33949 14323 33983
rect 14323 33949 14332 33983
rect 14280 33940 14332 33949
rect 16672 33983 16724 33992
rect 16672 33949 16681 33983
rect 16681 33949 16715 33983
rect 16715 33949 16724 33983
rect 16672 33940 16724 33949
rect 6552 33872 6604 33924
rect 7104 33872 7156 33924
rect 10324 33872 10376 33924
rect 12164 33872 12216 33924
rect 12256 33872 12308 33924
rect 12900 33872 12952 33924
rect 12992 33915 13044 33924
rect 12992 33881 13001 33915
rect 13001 33881 13035 33915
rect 13035 33881 13044 33915
rect 12992 33872 13044 33881
rect 13912 33872 13964 33924
rect 14648 33872 14700 33924
rect 16120 33872 16172 33924
rect 16488 33872 16540 33924
rect 17408 33872 17460 33924
rect 19708 33872 19760 33924
rect 20812 33872 20864 33924
rect 9680 33804 9732 33856
rect 10784 33804 10836 33856
rect 11428 33847 11480 33856
rect 11428 33813 11437 33847
rect 11437 33813 11471 33847
rect 11471 33813 11480 33847
rect 11428 33804 11480 33813
rect 12072 33804 12124 33856
rect 13360 33804 13412 33856
rect 17776 33804 17828 33856
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 27950 33702 28002 33754
rect 28014 33702 28066 33754
rect 28078 33702 28130 33754
rect 28142 33702 28194 33754
rect 28206 33702 28258 33754
rect 37950 33702 38002 33754
rect 38014 33702 38066 33754
rect 38078 33702 38130 33754
rect 38142 33702 38194 33754
rect 38206 33702 38258 33754
rect 47950 33702 48002 33754
rect 48014 33702 48066 33754
rect 48078 33702 48130 33754
rect 48142 33702 48194 33754
rect 48206 33702 48258 33754
rect 7196 33600 7248 33652
rect 7380 33600 7432 33652
rect 7564 33600 7616 33652
rect 6644 33575 6696 33584
rect 6644 33541 6653 33575
rect 6653 33541 6687 33575
rect 6687 33541 6696 33575
rect 6644 33532 6696 33541
rect 6828 33532 6880 33584
rect 6092 33464 6144 33516
rect 1308 33396 1360 33448
rect 7472 33396 7524 33448
rect 10324 33532 10376 33584
rect 9036 33507 9088 33516
rect 9036 33473 9045 33507
rect 9045 33473 9079 33507
rect 9079 33473 9088 33507
rect 9036 33464 9088 33473
rect 12900 33600 12952 33652
rect 15660 33600 15712 33652
rect 16764 33600 16816 33652
rect 18328 33600 18380 33652
rect 18512 33600 18564 33652
rect 21272 33600 21324 33652
rect 10784 33532 10836 33584
rect 11060 33507 11112 33516
rect 11060 33473 11069 33507
rect 11069 33473 11103 33507
rect 11103 33473 11112 33507
rect 11060 33464 11112 33473
rect 12256 33464 12308 33516
rect 8300 33328 8352 33380
rect 10048 33396 10100 33448
rect 13636 33532 13688 33584
rect 14280 33532 14332 33584
rect 16672 33532 16724 33584
rect 14004 33464 14056 33516
rect 14004 33328 14056 33380
rect 14740 33464 14792 33516
rect 15384 33507 15436 33516
rect 15384 33473 15393 33507
rect 15393 33473 15427 33507
rect 15427 33473 15436 33507
rect 15384 33464 15436 33473
rect 16488 33464 16540 33516
rect 17592 33507 17644 33516
rect 17592 33473 17601 33507
rect 17601 33473 17635 33507
rect 17635 33473 17644 33507
rect 17592 33464 17644 33473
rect 18788 33507 18840 33516
rect 18788 33473 18797 33507
rect 18797 33473 18831 33507
rect 18831 33473 18840 33507
rect 18788 33464 18840 33473
rect 15108 33396 15160 33448
rect 19432 33464 19484 33516
rect 20444 33464 20496 33516
rect 19064 33439 19116 33448
rect 19064 33405 19073 33439
rect 19073 33405 19107 33439
rect 19107 33405 19116 33439
rect 19064 33396 19116 33405
rect 18420 33328 18472 33380
rect 5632 33260 5684 33312
rect 10416 33260 10468 33312
rect 17132 33260 17184 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 32950 33158 33002 33210
rect 33014 33158 33066 33210
rect 33078 33158 33130 33210
rect 33142 33158 33194 33210
rect 33206 33158 33258 33210
rect 42950 33158 43002 33210
rect 43014 33158 43066 33210
rect 43078 33158 43130 33210
rect 43142 33158 43194 33210
rect 43206 33158 43258 33210
rect 7564 33056 7616 33108
rect 12348 33056 12400 33108
rect 14004 33056 14056 33108
rect 19156 33056 19208 33108
rect 9772 32988 9824 33040
rect 1308 32920 1360 32972
rect 7748 32920 7800 32972
rect 10876 32920 10928 32972
rect 4712 32852 4764 32904
rect 6920 32852 6972 32904
rect 9220 32852 9272 32904
rect 9864 32852 9916 32904
rect 10600 32852 10652 32904
rect 19248 32920 19300 32972
rect 11704 32895 11756 32904
rect 11704 32861 11713 32895
rect 11713 32861 11747 32895
rect 11747 32861 11756 32895
rect 11704 32852 11756 32861
rect 16488 32852 16540 32904
rect 22008 33056 22060 33108
rect 5448 32827 5500 32836
rect 5448 32793 5457 32827
rect 5457 32793 5491 32827
rect 5491 32793 5500 32827
rect 5448 32784 5500 32793
rect 7656 32784 7708 32836
rect 10692 32784 10744 32836
rect 11980 32827 12032 32836
rect 11980 32793 11989 32827
rect 11989 32793 12023 32827
rect 12023 32793 12032 32827
rect 11980 32784 12032 32793
rect 12716 32784 12768 32836
rect 5540 32759 5592 32768
rect 5540 32725 5549 32759
rect 5549 32725 5583 32759
rect 5583 32725 5592 32759
rect 5540 32716 5592 32725
rect 9312 32759 9364 32768
rect 9312 32725 9321 32759
rect 9321 32725 9355 32759
rect 9355 32725 9364 32759
rect 9312 32716 9364 32725
rect 10968 32759 11020 32768
rect 10968 32725 10977 32759
rect 10977 32725 11011 32759
rect 11011 32725 11020 32759
rect 10968 32716 11020 32725
rect 13820 32716 13872 32768
rect 14924 32716 14976 32768
rect 16856 32784 16908 32836
rect 17868 32784 17920 32836
rect 19524 32827 19576 32836
rect 19524 32793 19533 32827
rect 19533 32793 19567 32827
rect 19567 32793 19576 32827
rect 19524 32784 19576 32793
rect 15476 32759 15528 32768
rect 15476 32725 15485 32759
rect 15485 32725 15519 32759
rect 15519 32725 15528 32759
rect 15476 32716 15528 32725
rect 16028 32716 16080 32768
rect 18972 32716 19024 32768
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 27950 32614 28002 32666
rect 28014 32614 28066 32666
rect 28078 32614 28130 32666
rect 28142 32614 28194 32666
rect 28206 32614 28258 32666
rect 37950 32614 38002 32666
rect 38014 32614 38066 32666
rect 38078 32614 38130 32666
rect 38142 32614 38194 32666
rect 38206 32614 38258 32666
rect 47950 32614 48002 32666
rect 48014 32614 48066 32666
rect 48078 32614 48130 32666
rect 48142 32614 48194 32666
rect 48206 32614 48258 32666
rect 8852 32555 8904 32564
rect 8852 32521 8861 32555
rect 8861 32521 8895 32555
rect 8895 32521 8904 32555
rect 8852 32512 8904 32521
rect 9220 32555 9272 32564
rect 9220 32521 9229 32555
rect 9229 32521 9263 32555
rect 9263 32521 9272 32555
rect 9220 32512 9272 32521
rect 9680 32512 9732 32564
rect 10416 32555 10468 32564
rect 10416 32521 10425 32555
rect 10425 32521 10459 32555
rect 10459 32521 10468 32555
rect 10416 32512 10468 32521
rect 11704 32512 11756 32564
rect 5448 32444 5500 32496
rect 6920 32240 6972 32292
rect 7472 32240 7524 32292
rect 7840 32240 7892 32292
rect 9128 32376 9180 32428
rect 11888 32419 11940 32428
rect 11888 32385 11897 32419
rect 11897 32385 11931 32419
rect 11931 32385 11940 32419
rect 11888 32376 11940 32385
rect 14280 32512 14332 32564
rect 14464 32512 14516 32564
rect 14648 32512 14700 32564
rect 14832 32512 14884 32564
rect 12716 32444 12768 32496
rect 17408 32444 17460 32496
rect 18420 32512 18472 32564
rect 19064 32512 19116 32564
rect 20628 32512 20680 32564
rect 14464 32376 14516 32428
rect 20720 32376 20772 32428
rect 8944 32308 8996 32360
rect 11336 32240 11388 32292
rect 7656 32215 7708 32224
rect 7656 32181 7665 32215
rect 7665 32181 7699 32215
rect 7699 32181 7708 32215
rect 7656 32172 7708 32181
rect 11244 32172 11296 32224
rect 12624 32351 12676 32360
rect 12624 32317 12633 32351
rect 12633 32317 12667 32351
rect 12667 32317 12676 32351
rect 12624 32308 12676 32317
rect 13360 32308 13412 32360
rect 13820 32308 13872 32360
rect 12624 32172 12676 32224
rect 13820 32172 13872 32224
rect 14924 32308 14976 32360
rect 14924 32172 14976 32224
rect 16948 32172 17000 32224
rect 17500 32308 17552 32360
rect 17868 32308 17920 32360
rect 17868 32172 17920 32224
rect 21456 32308 21508 32360
rect 19708 32172 19760 32224
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 32950 32070 33002 32122
rect 33014 32070 33066 32122
rect 33078 32070 33130 32122
rect 33142 32070 33194 32122
rect 33206 32070 33258 32122
rect 42950 32070 43002 32122
rect 43014 32070 43066 32122
rect 43078 32070 43130 32122
rect 43142 32070 43194 32122
rect 43206 32070 43258 32122
rect 1308 31832 1360 31884
rect 6920 31875 6972 31884
rect 6920 31841 6929 31875
rect 6929 31841 6963 31875
rect 6963 31841 6972 31875
rect 6920 31832 6972 31841
rect 10600 31968 10652 32020
rect 10876 32011 10928 32020
rect 10876 31977 10885 32011
rect 10885 31977 10919 32011
rect 10919 31977 10928 32011
rect 10876 31968 10928 31977
rect 13728 31968 13780 32020
rect 14924 32011 14976 32020
rect 14924 31977 14933 32011
rect 14933 31977 14967 32011
rect 14967 31977 14976 32011
rect 14924 31968 14976 31977
rect 11980 31900 12032 31952
rect 10140 31832 10192 31884
rect 12348 31832 12400 31884
rect 15292 31832 15344 31884
rect 16028 31832 16080 31884
rect 16764 31968 16816 32020
rect 17500 31968 17552 32020
rect 17684 31968 17736 32020
rect 17776 31832 17828 31884
rect 5632 31764 5684 31816
rect 11704 31764 11756 31816
rect 7104 31628 7156 31680
rect 7748 31628 7800 31680
rect 10416 31696 10468 31748
rect 12532 31696 12584 31748
rect 12716 31696 12768 31748
rect 15660 31696 15712 31748
rect 10232 31628 10284 31680
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 27950 31526 28002 31578
rect 28014 31526 28066 31578
rect 28078 31526 28130 31578
rect 28142 31526 28194 31578
rect 28206 31526 28258 31578
rect 37950 31526 38002 31578
rect 38014 31526 38066 31578
rect 38078 31526 38130 31578
rect 38142 31526 38194 31578
rect 38206 31526 38258 31578
rect 47950 31526 48002 31578
rect 48014 31526 48066 31578
rect 48078 31526 48130 31578
rect 48142 31526 48194 31578
rect 48206 31526 48258 31578
rect 12716 31424 12768 31476
rect 10416 31356 10468 31408
rect 10692 31356 10744 31408
rect 12532 31356 12584 31408
rect 13544 31356 13596 31408
rect 15108 31424 15160 31476
rect 19432 31467 19484 31476
rect 19432 31433 19441 31467
rect 19441 31433 19475 31467
rect 19475 31433 19484 31467
rect 19432 31424 19484 31433
rect 14924 31356 14976 31408
rect 5540 31288 5592 31340
rect 16764 31288 16816 31340
rect 17868 31356 17920 31408
rect 18420 31356 18472 31408
rect 1308 31220 1360 31272
rect 8392 31220 8444 31272
rect 11336 31220 11388 31272
rect 11704 31263 11756 31272
rect 11704 31229 11713 31263
rect 11713 31229 11747 31263
rect 11747 31229 11756 31263
rect 11704 31220 11756 31229
rect 13544 31220 13596 31272
rect 14556 31263 14608 31272
rect 14556 31229 14565 31263
rect 14565 31229 14599 31263
rect 14599 31229 14608 31263
rect 14556 31220 14608 31229
rect 14832 31263 14884 31272
rect 14832 31229 14841 31263
rect 14841 31229 14875 31263
rect 14875 31229 14884 31263
rect 14832 31220 14884 31229
rect 17500 31220 17552 31272
rect 18328 31220 18380 31272
rect 20628 31220 20680 31272
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 32950 30982 33002 31034
rect 33014 30982 33066 31034
rect 33078 30982 33130 31034
rect 33142 30982 33194 31034
rect 33206 30982 33258 31034
rect 42950 30982 43002 31034
rect 43014 30982 43066 31034
rect 43078 30982 43130 31034
rect 43142 30982 43194 31034
rect 43206 30982 43258 31034
rect 9772 30880 9824 30932
rect 14924 30880 14976 30932
rect 15660 30880 15712 30932
rect 16856 30880 16908 30932
rect 7748 30812 7800 30864
rect 7840 30744 7892 30796
rect 10140 30744 10192 30796
rect 11704 30744 11756 30796
rect 14556 30744 14608 30796
rect 16764 30744 16816 30796
rect 7656 30676 7708 30728
rect 9496 30719 9548 30728
rect 9496 30685 9505 30719
rect 9505 30685 9539 30719
rect 9539 30685 9548 30719
rect 9496 30676 9548 30685
rect 14464 30719 14516 30728
rect 14464 30685 14473 30719
rect 14473 30685 14507 30719
rect 14507 30685 14516 30719
rect 14464 30676 14516 30685
rect 11060 30608 11112 30660
rect 11612 30608 11664 30660
rect 11888 30540 11940 30592
rect 12624 30583 12676 30592
rect 12624 30549 12633 30583
rect 12633 30549 12667 30583
rect 12667 30549 12676 30583
rect 12624 30540 12676 30549
rect 15108 30608 15160 30660
rect 15660 30608 15712 30660
rect 15384 30540 15436 30592
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 27950 30438 28002 30490
rect 28014 30438 28066 30490
rect 28078 30438 28130 30490
rect 28142 30438 28194 30490
rect 28206 30438 28258 30490
rect 37950 30438 38002 30490
rect 38014 30438 38066 30490
rect 38078 30438 38130 30490
rect 38142 30438 38194 30490
rect 38206 30438 38258 30490
rect 47950 30438 48002 30490
rect 48014 30438 48066 30490
rect 48078 30438 48130 30490
rect 48142 30438 48194 30490
rect 48206 30438 48258 30490
rect 10416 30336 10468 30388
rect 11060 30336 11112 30388
rect 11704 30336 11756 30388
rect 10048 30311 10100 30320
rect 10048 30277 10057 30311
rect 10057 30277 10091 30311
rect 10091 30277 10100 30311
rect 10048 30268 10100 30277
rect 11612 30268 11664 30320
rect 12532 30268 12584 30320
rect 1768 30243 1820 30252
rect 1768 30209 1777 30243
rect 1777 30209 1811 30243
rect 1811 30209 1820 30243
rect 1768 30200 1820 30209
rect 9588 30200 9640 30252
rect 11796 30243 11848 30252
rect 11796 30209 11805 30243
rect 11805 30209 11839 30243
rect 11839 30209 11848 30243
rect 11796 30200 11848 30209
rect 1308 30132 1360 30184
rect 9680 30132 9732 30184
rect 12624 30132 12676 30184
rect 13544 30175 13596 30184
rect 13544 30141 13553 30175
rect 13553 30141 13587 30175
rect 13587 30141 13596 30175
rect 13544 30132 13596 30141
rect 13820 30132 13872 30184
rect 17316 30132 17368 30184
rect 14096 30064 14148 30116
rect 8392 29996 8444 30048
rect 9036 29996 9088 30048
rect 14648 29996 14700 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 32950 29894 33002 29946
rect 33014 29894 33066 29946
rect 33078 29894 33130 29946
rect 33142 29894 33194 29946
rect 33206 29894 33258 29946
rect 42950 29894 43002 29946
rect 43014 29894 43066 29946
rect 43078 29894 43130 29946
rect 43142 29894 43194 29946
rect 43206 29894 43258 29946
rect 1768 29792 1820 29844
rect 9036 29792 9088 29844
rect 11152 29792 11204 29844
rect 11336 29792 11388 29844
rect 14372 29792 14424 29844
rect 10048 29656 10100 29708
rect 11796 29656 11848 29708
rect 13268 29656 13320 29708
rect 13728 29656 13780 29708
rect 16120 29656 16172 29708
rect 11888 29631 11940 29640
rect 11888 29597 11897 29631
rect 11897 29597 11931 29631
rect 11931 29597 11940 29631
rect 11888 29588 11940 29597
rect 14464 29588 14516 29640
rect 14740 29588 14792 29640
rect 1308 29520 1360 29572
rect 10048 29520 10100 29572
rect 10416 29520 10468 29572
rect 13728 29520 13780 29572
rect 10600 29452 10652 29504
rect 14740 29495 14792 29504
rect 14740 29461 14749 29495
rect 14749 29461 14783 29495
rect 14783 29461 14792 29495
rect 14740 29452 14792 29461
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 27950 29350 28002 29402
rect 28014 29350 28066 29402
rect 28078 29350 28130 29402
rect 28142 29350 28194 29402
rect 28206 29350 28258 29402
rect 37950 29350 38002 29402
rect 38014 29350 38066 29402
rect 38078 29350 38130 29402
rect 38142 29350 38194 29402
rect 38206 29350 38258 29402
rect 47950 29350 48002 29402
rect 48014 29350 48066 29402
rect 48078 29350 48130 29402
rect 48142 29350 48194 29402
rect 48206 29350 48258 29402
rect 8392 29248 8444 29300
rect 9588 29248 9640 29300
rect 9956 29248 10008 29300
rect 15016 29248 15068 29300
rect 7748 29223 7800 29232
rect 7748 29189 7757 29223
rect 7757 29189 7791 29223
rect 7791 29189 7800 29223
rect 7748 29180 7800 29189
rect 10048 29180 10100 29232
rect 12624 29180 12676 29232
rect 10600 29112 10652 29164
rect 9680 29044 9732 29096
rect 10692 29087 10744 29096
rect 10692 29053 10701 29087
rect 10701 29053 10735 29087
rect 10735 29053 10744 29087
rect 10692 29044 10744 29053
rect 12532 29044 12584 29096
rect 12808 29044 12860 29096
rect 13360 29087 13412 29096
rect 13360 29053 13369 29087
rect 13369 29053 13403 29087
rect 13403 29053 13412 29087
rect 13360 29044 13412 29053
rect 12072 28976 12124 29028
rect 8208 28908 8260 28960
rect 12808 28908 12860 28960
rect 14004 28908 14056 28960
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 32950 28806 33002 28858
rect 33014 28806 33066 28858
rect 33078 28806 33130 28858
rect 33142 28806 33194 28858
rect 33206 28806 33258 28858
rect 42950 28806 43002 28858
rect 43014 28806 43066 28858
rect 43078 28806 43130 28858
rect 43142 28806 43194 28858
rect 43206 28806 43258 28858
rect 7840 28747 7892 28756
rect 7840 28713 7849 28747
rect 7849 28713 7883 28747
rect 7883 28713 7892 28747
rect 7840 28704 7892 28713
rect 10692 28704 10744 28756
rect 13360 28704 13412 28756
rect 13544 28704 13596 28756
rect 7472 28636 7524 28688
rect 1308 28568 1360 28620
rect 7564 28568 7616 28620
rect 11612 28636 11664 28688
rect 10232 28568 10284 28620
rect 1768 28543 1820 28552
rect 1768 28509 1777 28543
rect 1777 28509 1811 28543
rect 1811 28509 1820 28543
rect 1768 28500 1820 28509
rect 7748 28500 7800 28552
rect 8208 28543 8260 28552
rect 8208 28509 8217 28543
rect 8217 28509 8251 28543
rect 8251 28509 8260 28543
rect 8208 28500 8260 28509
rect 11428 28500 11480 28552
rect 11704 28611 11756 28620
rect 11704 28577 11713 28611
rect 11713 28577 11747 28611
rect 11747 28577 11756 28611
rect 11704 28568 11756 28577
rect 11980 28500 12032 28552
rect 12440 28568 12492 28620
rect 15292 28500 15344 28552
rect 10232 28475 10284 28484
rect 10232 28441 10241 28475
rect 10241 28441 10275 28475
rect 10275 28441 10284 28475
rect 10232 28432 10284 28441
rect 14740 28432 14792 28484
rect 12716 28407 12768 28416
rect 12716 28373 12725 28407
rect 12725 28373 12759 28407
rect 12759 28373 12768 28407
rect 12716 28364 12768 28373
rect 19892 28364 19944 28416
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 27950 28262 28002 28314
rect 28014 28262 28066 28314
rect 28078 28262 28130 28314
rect 28142 28262 28194 28314
rect 28206 28262 28258 28314
rect 37950 28262 38002 28314
rect 38014 28262 38066 28314
rect 38078 28262 38130 28314
rect 38142 28262 38194 28314
rect 38206 28262 38258 28314
rect 47950 28262 48002 28314
rect 48014 28262 48066 28314
rect 48078 28262 48130 28314
rect 48142 28262 48194 28314
rect 48206 28262 48258 28314
rect 9772 28203 9824 28212
rect 9772 28169 9781 28203
rect 9781 28169 9815 28203
rect 9815 28169 9824 28203
rect 9772 28160 9824 28169
rect 9864 28203 9916 28212
rect 9864 28169 9873 28203
rect 9873 28169 9907 28203
rect 9907 28169 9916 28203
rect 9864 28160 9916 28169
rect 12808 28160 12860 28212
rect 12624 28092 12676 28144
rect 20996 28024 21048 28076
rect 1308 27956 1360 28008
rect 9680 27888 9732 27940
rect 13636 27956 13688 28008
rect 9404 27863 9456 27872
rect 9404 27829 9413 27863
rect 9413 27829 9447 27863
rect 9447 27829 9456 27863
rect 9404 27820 9456 27829
rect 15108 27820 15160 27872
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 32950 27718 33002 27770
rect 33014 27718 33066 27770
rect 33078 27718 33130 27770
rect 33142 27718 33194 27770
rect 33206 27718 33258 27770
rect 42950 27718 43002 27770
rect 43014 27718 43066 27770
rect 43078 27718 43130 27770
rect 43142 27718 43194 27770
rect 43206 27718 43258 27770
rect 11520 27548 11572 27600
rect 12348 27523 12400 27532
rect 12348 27489 12357 27523
rect 12357 27489 12391 27523
rect 12391 27489 12400 27523
rect 12348 27480 12400 27489
rect 14188 27412 14240 27464
rect 1676 27276 1728 27328
rect 18696 27344 18748 27396
rect 17132 27276 17184 27328
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 27950 27174 28002 27226
rect 28014 27174 28066 27226
rect 28078 27174 28130 27226
rect 28142 27174 28194 27226
rect 28206 27174 28258 27226
rect 37950 27174 38002 27226
rect 38014 27174 38066 27226
rect 38078 27174 38130 27226
rect 38142 27174 38194 27226
rect 38206 27174 38258 27226
rect 47950 27174 48002 27226
rect 48014 27174 48066 27226
rect 48078 27174 48130 27226
rect 48142 27174 48194 27226
rect 48206 27174 48258 27226
rect 12072 27115 12124 27124
rect 12072 27081 12081 27115
rect 12081 27081 12115 27115
rect 12115 27081 12124 27115
rect 12072 27072 12124 27081
rect 6460 27004 6512 27056
rect 9312 27004 9364 27056
rect 940 26936 992 26988
rect 11336 26936 11388 26988
rect 16212 26732 16264 26784
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 32950 26630 33002 26682
rect 33014 26630 33066 26682
rect 33078 26630 33130 26682
rect 33142 26630 33194 26682
rect 33206 26630 33258 26682
rect 42950 26630 43002 26682
rect 43014 26630 43066 26682
rect 43078 26630 43130 26682
rect 43142 26630 43194 26682
rect 43206 26630 43258 26682
rect 1860 26435 1912 26444
rect 1860 26401 1869 26435
rect 1869 26401 1903 26435
rect 1903 26401 1912 26435
rect 1860 26392 1912 26401
rect 1584 26367 1636 26376
rect 1584 26333 1593 26367
rect 1593 26333 1627 26367
rect 1627 26333 1636 26367
rect 1584 26324 1636 26333
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 27950 26086 28002 26138
rect 28014 26086 28066 26138
rect 28078 26086 28130 26138
rect 28142 26086 28194 26138
rect 28206 26086 28258 26138
rect 37950 26086 38002 26138
rect 38014 26086 38066 26138
rect 38078 26086 38130 26138
rect 38142 26086 38194 26138
rect 38206 26086 38258 26138
rect 47950 26086 48002 26138
rect 48014 26086 48066 26138
rect 48078 26086 48130 26138
rect 48142 26086 48194 26138
rect 48206 26086 48258 26138
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 32950 25542 33002 25594
rect 33014 25542 33066 25594
rect 33078 25542 33130 25594
rect 33142 25542 33194 25594
rect 33206 25542 33258 25594
rect 42950 25542 43002 25594
rect 43014 25542 43066 25594
rect 43078 25542 43130 25594
rect 43142 25542 43194 25594
rect 43206 25542 43258 25594
rect 12532 25440 12584 25492
rect 4988 25304 5040 25356
rect 10876 25347 10928 25356
rect 10876 25313 10885 25347
rect 10885 25313 10919 25347
rect 10919 25313 10928 25347
rect 10876 25304 10928 25313
rect 940 25236 992 25288
rect 10324 25100 10376 25152
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 27950 24998 28002 25050
rect 28014 24998 28066 25050
rect 28078 24998 28130 25050
rect 28142 24998 28194 25050
rect 28206 24998 28258 25050
rect 37950 24998 38002 25050
rect 38014 24998 38066 25050
rect 38078 24998 38130 25050
rect 38142 24998 38194 25050
rect 38206 24998 38258 25050
rect 47950 24998 48002 25050
rect 48014 24998 48066 25050
rect 48078 24998 48130 25050
rect 48142 24998 48194 25050
rect 48206 24998 48258 25050
rect 1584 24896 1636 24948
rect 10324 24896 10376 24948
rect 940 24760 992 24812
rect 4896 24760 4948 24812
rect 33692 24760 33744 24812
rect 24124 24692 24176 24744
rect 24676 24692 24728 24744
rect 26424 24624 26476 24676
rect 34336 24735 34388 24744
rect 34336 24701 34345 24735
rect 34345 24701 34379 24735
rect 34379 24701 34388 24735
rect 34336 24692 34388 24701
rect 47860 24692 47912 24744
rect 10784 24556 10836 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 13912 24352 13964 24404
rect 14832 24216 14884 24268
rect 10784 24191 10836 24200
rect 10784 24157 10793 24191
rect 10793 24157 10827 24191
rect 10827 24157 10836 24191
rect 10784 24148 10836 24157
rect 12440 24191 12492 24200
rect 12440 24157 12449 24191
rect 12449 24157 12483 24191
rect 12483 24157 12492 24191
rect 12440 24148 12492 24157
rect 12808 24148 12860 24200
rect 13820 24148 13872 24200
rect 10876 24055 10928 24064
rect 10876 24021 10885 24055
rect 10885 24021 10919 24055
rect 10919 24021 10928 24055
rect 10876 24012 10928 24021
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 18788 23808 18840 23860
rect 3516 23672 3568 23724
rect 940 23604 992 23656
rect 12532 23647 12584 23656
rect 12532 23613 12541 23647
rect 12541 23613 12575 23647
rect 12575 23613 12584 23647
rect 12532 23604 12584 23613
rect 17408 23604 17460 23656
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 17592 23264 17644 23316
rect 5908 23128 5960 23180
rect 18328 23128 18380 23180
rect 940 23060 992 23112
rect 12440 22992 12492 23044
rect 12348 22967 12400 22976
rect 12348 22933 12357 22967
rect 12357 22933 12391 22967
rect 12391 22933 12400 22967
rect 12348 22924 12400 22933
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 3424 22040 3476 22092
rect 940 21972 992 22024
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 4804 21496 4856 21548
rect 940 21428 992 21480
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 19156 21020 19208 21072
rect 9404 20884 9456 20936
rect 15108 20884 15160 20936
rect 18604 20748 18656 20800
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 7104 20408 7156 20460
rect 16212 20451 16264 20460
rect 16212 20417 16221 20451
rect 16221 20417 16255 20451
rect 16255 20417 16264 20451
rect 16212 20408 16264 20417
rect 25872 20408 25924 20460
rect 940 20340 992 20392
rect 18696 20204 18748 20256
rect 23572 20204 23624 20256
rect 34336 20204 34388 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 1860 19975 1912 19984
rect 1860 19941 1869 19975
rect 1869 19941 1903 19975
rect 1903 19941 1912 19975
rect 1860 19932 1912 19941
rect 940 19728 992 19780
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 8392 18912 8444 18964
rect 940 18708 992 18760
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 8668 18368 8720 18420
rect 1768 18275 1820 18284
rect 1768 18241 1777 18275
rect 1777 18241 1811 18275
rect 1811 18241 1820 18275
rect 1768 18232 1820 18241
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 25412 17731 25464 17740
rect 25412 17697 25421 17731
rect 25421 17697 25455 17731
rect 25455 17697 25464 17731
rect 25412 17688 25464 17697
rect 26148 17688 26200 17740
rect 24952 17663 25004 17672
rect 24952 17629 24961 17663
rect 24961 17629 24995 17663
rect 24995 17629 25004 17663
rect 24952 17620 25004 17629
rect 27252 17663 27304 17672
rect 27252 17629 27261 17663
rect 27261 17629 27295 17663
rect 27295 17629 27304 17663
rect 27252 17620 27304 17629
rect 25136 17595 25188 17604
rect 25136 17561 25145 17595
rect 25145 17561 25179 17595
rect 25179 17561 25188 17595
rect 25136 17552 25188 17561
rect 24492 17484 24544 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 26424 17323 26476 17332
rect 26424 17289 26433 17323
rect 26433 17289 26467 17323
rect 26467 17289 26476 17323
rect 26424 17280 26476 17289
rect 20720 17212 20772 17264
rect 30748 17255 30800 17264
rect 30748 17221 30757 17255
rect 30757 17221 30791 17255
rect 30791 17221 30800 17255
rect 30748 17212 30800 17221
rect 940 17144 992 17196
rect 17132 17187 17184 17196
rect 17132 17153 17141 17187
rect 17141 17153 17175 17187
rect 17175 17153 17184 17187
rect 17132 17144 17184 17153
rect 1860 17119 1912 17128
rect 1860 17085 1869 17119
rect 1869 17085 1903 17119
rect 1903 17085 1912 17119
rect 1860 17076 1912 17085
rect 15844 17076 15896 17128
rect 23572 17144 23624 17196
rect 24676 17187 24728 17196
rect 24676 17153 24685 17187
rect 24685 17153 24719 17187
rect 24719 17153 24728 17187
rect 24676 17144 24728 17153
rect 28908 17119 28960 17128
rect 28908 17085 28917 17119
rect 28917 17085 28951 17119
rect 28951 17085 28960 17119
rect 28908 17076 28960 17085
rect 29092 17119 29144 17128
rect 29092 17085 29101 17119
rect 29101 17085 29135 17119
rect 29135 17085 29144 17119
rect 29092 17076 29144 17085
rect 24676 17008 24728 17060
rect 17776 16983 17828 16992
rect 17776 16949 17785 16983
rect 17785 16949 17819 16983
rect 17819 16949 17828 16983
rect 17776 16940 17828 16949
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 1952 16668 2004 16720
rect 31024 16643 31076 16652
rect 31024 16609 31033 16643
rect 31033 16609 31067 16643
rect 31067 16609 31076 16643
rect 31024 16600 31076 16609
rect 23572 16575 23624 16584
rect 23572 16541 23616 16575
rect 23616 16541 23624 16575
rect 23572 16532 23624 16541
rect 25136 16532 25188 16584
rect 32864 16575 32916 16584
rect 32864 16541 32873 16575
rect 32873 16541 32907 16575
rect 32907 16541 32916 16575
rect 32864 16532 32916 16541
rect 940 16464 992 16516
rect 31208 16507 31260 16516
rect 31208 16473 31217 16507
rect 31217 16473 31251 16507
rect 31251 16473 31260 16507
rect 31208 16464 31260 16473
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 26424 15648 26476 15700
rect 7656 15580 7708 15632
rect 25872 15487 25924 15496
rect 25872 15453 25881 15487
rect 25881 15453 25915 15487
rect 25915 15453 25924 15487
rect 25872 15444 25924 15453
rect 940 15376 992 15428
rect 25964 15308 26016 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 24492 15104 24544 15156
rect 6920 14968 6972 15020
rect 17868 14968 17920 15020
rect 25964 14968 26016 15020
rect 940 14900 992 14952
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 25044 14356 25096 14408
rect 29092 14220 29144 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 1676 14016 1728 14068
rect 20904 14016 20956 14068
rect 24676 14016 24728 14068
rect 31208 14016 31260 14068
rect 20720 13948 20772 14000
rect 940 13880 992 13932
rect 18604 13923 18656 13932
rect 18604 13889 18613 13923
rect 18613 13889 18647 13923
rect 18647 13889 18656 13923
rect 18604 13880 18656 13889
rect 19708 13923 19760 13932
rect 19708 13889 19717 13923
rect 19717 13889 19751 13923
rect 19751 13889 19760 13923
rect 19708 13880 19760 13889
rect 26700 13880 26752 13932
rect 17224 13812 17276 13864
rect 17868 13812 17920 13864
rect 20628 13676 20680 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 24676 13515 24728 13524
rect 24676 13481 24685 13515
rect 24685 13481 24719 13515
rect 24719 13481 24728 13515
rect 24676 13472 24728 13481
rect 940 13268 992 13320
rect 23388 13268 23440 13320
rect 25872 13268 25924 13320
rect 12716 13132 12768 13184
rect 19340 13132 19392 13184
rect 25044 13175 25096 13184
rect 25044 13141 25053 13175
rect 25053 13141 25087 13175
rect 25087 13141 25096 13175
rect 25044 13132 25096 13141
rect 45560 13132 45612 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 18696 12860 18748 12912
rect 19156 12835 19208 12844
rect 19156 12801 19165 12835
rect 19165 12801 19199 12835
rect 19199 12801 19208 12835
rect 19156 12792 19208 12801
rect 19340 12767 19392 12776
rect 19340 12733 19349 12767
rect 19349 12733 19383 12767
rect 19383 12733 19392 12767
rect 19340 12724 19392 12733
rect 21364 12724 21416 12776
rect 22652 12656 22704 12708
rect 24124 12588 24176 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 21364 12384 21416 12436
rect 26700 12384 26752 12436
rect 940 12112 992 12164
rect 11980 12044 12032 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 940 11704 992 11756
rect 10968 11500 11020 11552
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 20628 11296 20680 11348
rect 21364 11160 21416 11212
rect 23388 11092 23440 11144
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 940 10616 992 10668
rect 12808 10412 12860 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 940 9936 992 9988
rect 10692 9868 10744 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 1584 9163 1636 9172
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 940 8916 992 8968
rect 17776 8916 17828 8968
rect 19432 8848 19484 8900
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 1768 8483 1820 8492
rect 1768 8449 1777 8483
rect 1777 8449 1811 8483
rect 1811 8449 1820 8483
rect 1768 8440 1820 8449
rect 10876 8304 10928 8356
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 6920 8032 6972 8084
rect 9588 7896 9640 7948
rect 20720 7896 20772 7948
rect 15844 7828 15896 7880
rect 10692 7803 10744 7812
rect 10692 7769 10701 7803
rect 10701 7769 10735 7803
rect 10735 7769 10744 7803
rect 10692 7760 10744 7769
rect 20628 7760 20680 7812
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 940 7352 992 7404
rect 10232 7148 10284 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 7748 6808 7800 6860
rect 17224 6740 17276 6792
rect 20904 6783 20956 6792
rect 20904 6749 20913 6783
rect 20913 6749 20947 6783
rect 20947 6749 20956 6783
rect 20904 6740 20956 6749
rect 22652 6783 22704 6792
rect 22652 6749 22661 6783
rect 22661 6749 22695 6783
rect 22695 6749 22704 6783
rect 22652 6740 22704 6749
rect 940 6672 992 6724
rect 15292 6672 15344 6724
rect 22192 6672 22244 6724
rect 23480 6672 23532 6724
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 19340 6332 19392 6384
rect 24124 6332 24176 6384
rect 28816 6128 28868 6180
rect 15200 6060 15252 6112
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 21364 5652 21416 5704
rect 940 5584 992 5636
rect 11520 5516 11572 5568
rect 18328 5516 18380 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 9220 5244 9272 5296
rect 940 5176 992 5228
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 940 4020 992 4072
rect 12348 4020 12400 4072
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 940 3476 992 3528
rect 12532 3476 12584 3528
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 28816 3043 28868 3052
rect 28816 3009 28825 3043
rect 28825 3009 28859 3043
rect 28859 3009 28868 3043
rect 28816 3000 28868 3009
rect 48596 3000 48648 3052
rect 28724 2932 28776 2984
rect 19524 2796 19576 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 31024 2592 31076 2644
rect 24952 2524 25004 2576
rect 5540 2456 5592 2508
rect 8852 2456 8904 2508
rect 12164 2456 12216 2508
rect 2228 2388 2280 2440
rect 6920 2388 6972 2440
rect 15200 2456 15252 2508
rect 15476 2499 15528 2508
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 18788 2456 18840 2508
rect 22100 2456 22152 2508
rect 25412 2456 25464 2508
rect 28908 2524 28960 2576
rect 45560 2635 45612 2644
rect 45560 2601 45569 2635
rect 45569 2601 45603 2635
rect 45603 2601 45612 2635
rect 45560 2592 45612 2601
rect 18328 2388 18380 2440
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 22192 2431 22244 2440
rect 22192 2397 22201 2431
rect 22201 2397 22235 2431
rect 22235 2397 22244 2431
rect 22192 2388 22244 2397
rect 23480 2388 23532 2440
rect 32036 2388 32088 2440
rect 35348 2388 35400 2440
rect 15292 2320 15344 2372
rect 27252 2320 27304 2372
rect 38660 2431 38712 2440
rect 38660 2397 38669 2431
rect 38669 2397 38703 2431
rect 38703 2397 38712 2431
rect 38660 2388 38712 2397
rect 41972 2388 42024 2440
rect 45284 2320 45336 2372
rect 10692 2252 10744 2304
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
<< metal2 >>
rect 1582 56200 1638 57000
rect 2226 56200 2282 57000
rect 2870 56200 2926 57000
rect 3514 56200 3570 57000
rect 4158 56200 4214 57000
rect 4802 56200 4858 57000
rect 5446 56200 5502 57000
rect 6090 56200 6146 57000
rect 6734 56200 6790 57000
rect 7378 56200 7434 57000
rect 8022 56200 8078 57000
rect 8666 56200 8722 57000
rect 9310 56200 9366 57000
rect 9954 56200 10010 57000
rect 10598 56200 10654 57000
rect 11242 56200 11298 57000
rect 11886 56200 11942 57000
rect 12530 56200 12586 57000
rect 13174 56200 13230 57000
rect 13818 56200 13874 57000
rect 14462 56200 14518 57000
rect 15106 56200 15162 57000
rect 15750 56200 15806 57000
rect 16394 56200 16450 57000
rect 17038 56200 17094 57000
rect 17682 56200 17738 57000
rect 18326 56200 18382 57000
rect 18970 56200 19026 57000
rect 19614 56200 19670 57000
rect 20258 56200 20314 57000
rect 20902 56200 20958 57000
rect 21546 56200 21602 57000
rect 22190 56200 22246 57000
rect 22834 56200 22890 57000
rect 23478 56200 23534 57000
rect 24122 56200 24178 57000
rect 24766 56200 24822 57000
rect 25410 56200 25466 57000
rect 26054 56200 26110 57000
rect 26698 56200 26754 57000
rect 27342 56200 27398 57000
rect 27986 56200 28042 57000
rect 28630 56200 28686 57000
rect 29274 56200 29330 57000
rect 29918 56200 29974 57000
rect 30024 56222 30328 56250
rect 1596 52562 1624 56200
rect 2240 53038 2268 56200
rect 2320 54188 2372 54194
rect 2320 54130 2372 54136
rect 2228 53032 2280 53038
rect 2228 52974 2280 52980
rect 1584 52556 1636 52562
rect 1584 52498 1636 52504
rect 1308 51468 1360 51474
rect 1308 51410 1360 51416
rect 1320 51377 1348 51410
rect 1306 51368 1362 51377
rect 1306 51303 1362 51312
rect 1308 50856 1360 50862
rect 1308 50798 1360 50804
rect 1320 50561 1348 50798
rect 1306 50552 1362 50561
rect 1306 50487 1362 50496
rect 1584 50448 1636 50454
rect 1584 50390 1636 50396
rect 1308 49768 1360 49774
rect 1306 49736 1308 49745
rect 1360 49736 1362 49745
rect 1306 49671 1362 49680
rect 1308 49292 1360 49298
rect 1308 49234 1360 49240
rect 1320 48929 1348 49234
rect 1306 48920 1362 48929
rect 1306 48855 1362 48864
rect 1308 48204 1360 48210
rect 1308 48146 1360 48152
rect 1320 48113 1348 48146
rect 1306 48104 1362 48113
rect 1306 48039 1362 48048
rect 1308 47592 1360 47598
rect 1308 47534 1360 47540
rect 1320 47297 1348 47534
rect 1306 47288 1362 47297
rect 1306 47223 1362 47232
rect 1308 46504 1360 46510
rect 1306 46472 1308 46481
rect 1360 46472 1362 46481
rect 1306 46407 1362 46416
rect 1308 46028 1360 46034
rect 1308 45970 1360 45976
rect 1320 45665 1348 45970
rect 1306 45656 1362 45665
rect 1306 45591 1362 45600
rect 1308 44940 1360 44946
rect 1308 44882 1360 44888
rect 1320 44849 1348 44882
rect 1306 44840 1362 44849
rect 1306 44775 1362 44784
rect 1308 43240 1360 43246
rect 1306 43208 1308 43217
rect 1360 43208 1362 43217
rect 1306 43143 1362 43152
rect 1308 42764 1360 42770
rect 1308 42706 1360 42712
rect 1320 42401 1348 42706
rect 1596 42702 1624 50390
rect 2332 46714 2360 54130
rect 2778 53816 2834 53825
rect 2778 53751 2834 53760
rect 2688 53100 2740 53106
rect 2688 53042 2740 53048
rect 2320 46708 2372 46714
rect 2320 46650 2372 46656
rect 2700 45558 2728 53042
rect 2792 52698 2820 53751
rect 2884 53650 2912 56200
rect 3422 54632 3478 54641
rect 3422 54567 3478 54576
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 2872 53644 2924 53650
rect 2872 53586 2924 53592
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 2780 52692 2832 52698
rect 2780 52634 2832 52640
rect 3330 52184 3386 52193
rect 3330 52119 3386 52128
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 3344 51474 3372 52119
rect 3332 51468 3384 51474
rect 3332 51410 3384 51416
rect 3436 51074 3464 54567
rect 3528 54262 3556 56200
rect 3516 54256 3568 54262
rect 3516 54198 3568 54204
rect 3606 53000 3662 53009
rect 3606 52935 3662 52944
rect 3436 51046 3556 51074
rect 3332 50924 3384 50930
rect 3332 50866 3384 50872
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 3344 46170 3372 50866
rect 3424 49224 3476 49230
rect 3424 49166 3476 49172
rect 3332 46164 3384 46170
rect 3332 46106 3384 46112
rect 2688 45552 2740 45558
rect 2688 45494 2740 45500
rect 2504 45484 2556 45490
rect 2504 45426 2556 45432
rect 2044 44328 2096 44334
rect 2044 44270 2096 44276
rect 2056 44033 2084 44270
rect 2042 44024 2098 44033
rect 2042 43959 2098 43968
rect 1584 42696 1636 42702
rect 1584 42638 1636 42644
rect 1306 42392 1362 42401
rect 1306 42327 1362 42336
rect 1768 41744 1820 41750
rect 1768 41686 1820 41692
rect 1308 41676 1360 41682
rect 1308 41618 1360 41624
rect 1320 41585 1348 41618
rect 1306 41576 1362 41585
rect 1306 41511 1362 41520
rect 1308 41064 1360 41070
rect 1308 41006 1360 41012
rect 1320 40769 1348 41006
rect 1306 40760 1362 40769
rect 1306 40695 1362 40704
rect 1308 39500 1360 39506
rect 1308 39442 1360 39448
rect 1320 39137 1348 39442
rect 1306 39128 1362 39137
rect 1306 39063 1362 39072
rect 1308 38412 1360 38418
rect 1308 38354 1360 38360
rect 1320 38321 1348 38354
rect 1306 38312 1362 38321
rect 1306 38247 1362 38256
rect 1308 37800 1360 37806
rect 1308 37742 1360 37748
rect 1320 37505 1348 37742
rect 1306 37496 1362 37505
rect 1306 37431 1362 37440
rect 1780 36786 1808 41686
rect 2044 39976 2096 39982
rect 2042 39944 2044 39953
rect 2096 39944 2098 39953
rect 2042 39879 2098 39888
rect 1860 39568 1912 39574
rect 1860 39510 1912 39516
rect 1768 36780 1820 36786
rect 1768 36722 1820 36728
rect 1308 36712 1360 36718
rect 1306 36680 1308 36689
rect 1360 36680 1362 36689
rect 1306 36615 1362 36624
rect 1308 35148 1360 35154
rect 1308 35090 1360 35096
rect 1320 35057 1348 35090
rect 1306 35048 1362 35057
rect 1306 34983 1362 34992
rect 1308 33448 1360 33454
rect 1306 33416 1308 33425
rect 1360 33416 1362 33425
rect 1306 33351 1362 33360
rect 1308 32972 1360 32978
rect 1308 32914 1360 32920
rect 1320 32609 1348 32914
rect 1306 32600 1362 32609
rect 1306 32535 1362 32544
rect 1308 31884 1360 31890
rect 1308 31826 1360 31832
rect 1320 31793 1348 31826
rect 1306 31784 1362 31793
rect 1306 31719 1362 31728
rect 1308 31272 1360 31278
rect 1308 31214 1360 31220
rect 1320 30977 1348 31214
rect 1306 30968 1362 30977
rect 1306 30903 1362 30912
rect 1768 30252 1820 30258
rect 1768 30194 1820 30200
rect 1308 30184 1360 30190
rect 1306 30152 1308 30161
rect 1360 30152 1362 30161
rect 1306 30087 1362 30096
rect 1780 29850 1808 30194
rect 1768 29844 1820 29850
rect 1768 29786 1820 29792
rect 1308 29572 1360 29578
rect 1308 29514 1360 29520
rect 1320 29345 1348 29514
rect 1306 29336 1362 29345
rect 1306 29271 1362 29280
rect 1766 28656 1822 28665
rect 1308 28620 1360 28626
rect 1766 28591 1822 28600
rect 1308 28562 1360 28568
rect 1320 28529 1348 28562
rect 1780 28558 1808 28591
rect 1768 28552 1820 28558
rect 1306 28520 1362 28529
rect 1768 28494 1820 28500
rect 1306 28455 1362 28464
rect 1308 28008 1360 28014
rect 1308 27950 1360 27956
rect 1320 27713 1348 27950
rect 1306 27704 1362 27713
rect 1306 27639 1362 27648
rect 1676 27328 1728 27334
rect 1676 27270 1728 27276
rect 940 26988 992 26994
rect 940 26930 992 26936
rect 952 26897 980 26930
rect 938 26888 994 26897
rect 938 26823 994 26832
rect 1584 26376 1636 26382
rect 1584 26318 1636 26324
rect 1596 26081 1624 26318
rect 1582 26072 1638 26081
rect 1582 26007 1638 26016
rect 940 25288 992 25294
rect 938 25256 940 25265
rect 992 25256 994 25265
rect 938 25191 994 25200
rect 1584 24948 1636 24954
rect 1584 24890 1636 24896
rect 940 24812 992 24818
rect 940 24754 992 24760
rect 952 24449 980 24754
rect 938 24440 994 24449
rect 938 24375 994 24384
rect 940 23656 992 23662
rect 938 23624 940 23633
rect 992 23624 994 23633
rect 938 23559 994 23568
rect 940 23112 992 23118
rect 940 23054 992 23060
rect 952 22817 980 23054
rect 938 22808 994 22817
rect 938 22743 994 22752
rect 940 22024 992 22030
rect 938 21992 940 22001
rect 992 21992 994 22001
rect 938 21927 994 21936
rect 940 21480 992 21486
rect 940 21422 992 21428
rect 952 21185 980 21422
rect 938 21176 994 21185
rect 938 21111 994 21120
rect 940 20392 992 20398
rect 938 20360 940 20369
rect 992 20360 994 20369
rect 938 20295 994 20304
rect 940 19780 992 19786
rect 940 19722 992 19728
rect 952 19553 980 19722
rect 938 19544 994 19553
rect 938 19479 994 19488
rect 940 18760 992 18766
rect 938 18728 940 18737
rect 992 18728 994 18737
rect 938 18663 994 18672
rect 940 17196 992 17202
rect 940 17138 992 17144
rect 952 17105 980 17138
rect 938 17096 994 17105
rect 938 17031 994 17040
rect 940 16516 992 16522
rect 940 16458 992 16464
rect 952 16289 980 16458
rect 938 16280 994 16289
rect 938 16215 994 16224
rect 938 15464 994 15473
rect 938 15399 940 15408
rect 992 15399 994 15408
rect 940 15370 992 15376
rect 940 14952 992 14958
rect 940 14894 992 14900
rect 952 14657 980 14894
rect 938 14648 994 14657
rect 938 14583 994 14592
rect 940 13932 992 13938
rect 940 13874 992 13880
rect 952 13841 980 13874
rect 938 13832 994 13841
rect 938 13767 994 13776
rect 940 13320 992 13326
rect 940 13262 992 13268
rect 952 13025 980 13262
rect 938 13016 994 13025
rect 938 12951 994 12960
rect 938 12200 994 12209
rect 938 12135 940 12144
rect 992 12135 994 12144
rect 940 12106 992 12112
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 952 11393 980 11698
rect 938 11384 994 11393
rect 938 11319 994 11328
rect 940 10668 992 10674
rect 940 10610 992 10616
rect 952 10577 980 10610
rect 938 10568 994 10577
rect 938 10503 994 10512
rect 940 9988 992 9994
rect 940 9930 992 9936
rect 952 9761 980 9930
rect 938 9752 994 9761
rect 938 9687 994 9696
rect 1596 9178 1624 24890
rect 1688 14074 1716 27270
rect 1872 26450 1900 39510
rect 2516 39506 2544 45426
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 3436 45082 3464 49166
rect 3528 45529 3556 51046
rect 3620 49298 3648 52935
rect 4172 52562 4200 56200
rect 4712 53576 4764 53582
rect 4712 53518 4764 53524
rect 4160 52556 4212 52562
rect 4160 52498 4212 52504
rect 4252 52488 4304 52494
rect 4252 52430 4304 52436
rect 3608 49292 3660 49298
rect 3608 49234 3660 49240
rect 3884 48136 3936 48142
rect 3884 48078 3936 48084
rect 3700 45960 3752 45966
rect 3700 45902 3752 45908
rect 3514 45520 3570 45529
rect 3514 45455 3570 45464
rect 3424 45076 3476 45082
rect 3424 45018 3476 45024
rect 3516 44396 3568 44402
rect 3516 44338 3568 44344
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 2504 39500 2556 39506
rect 2504 39442 2556 39448
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 3528 36718 3556 44338
rect 3712 42770 3740 45902
rect 3896 45558 3924 48078
rect 4160 47660 4212 47666
rect 4160 47602 4212 47608
rect 3884 45552 3936 45558
rect 3884 45494 3936 45500
rect 4172 44538 4200 47602
rect 4160 44532 4212 44538
rect 4160 44474 4212 44480
rect 4264 44470 4292 52430
rect 4620 49836 4672 49842
rect 4620 49778 4672 49784
rect 4528 46572 4580 46578
rect 4528 46514 4580 46520
rect 4436 46504 4488 46510
rect 4436 46446 4488 46452
rect 4344 44872 4396 44878
rect 4344 44814 4396 44820
rect 4252 44464 4304 44470
rect 4252 44406 4304 44412
rect 4160 44328 4212 44334
rect 4160 44270 4212 44276
rect 3700 42764 3752 42770
rect 3700 42706 3752 42712
rect 4172 42362 4200 44270
rect 4160 42356 4212 42362
rect 4160 42298 4212 42304
rect 4356 41818 4384 44814
rect 4448 43994 4476 46446
rect 4436 43988 4488 43994
rect 4436 43930 4488 43936
rect 4344 41812 4396 41818
rect 4344 41754 4396 41760
rect 4344 40112 4396 40118
rect 4344 40054 4396 40060
rect 3976 39908 4028 39914
rect 3976 39850 4028 39856
rect 3516 36712 3568 36718
rect 3516 36654 3568 36660
rect 3424 36644 3476 36650
rect 3424 36586 3476 36592
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 2780 36100 2832 36106
rect 2780 36042 2832 36048
rect 2792 35873 2820 36042
rect 2778 35864 2834 35873
rect 2778 35799 2834 35808
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 2044 34536 2096 34542
rect 2044 34478 2096 34484
rect 2056 34241 2084 34478
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 2042 34232 2098 34241
rect 2950 34235 3258 34244
rect 2042 34167 2098 34176
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 1860 26444 1912 26450
rect 1860 26386 1912 26392
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 3436 22098 3464 36586
rect 3528 23730 3556 36654
rect 3988 35086 4016 39850
rect 4068 39840 4120 39846
rect 4068 39782 4120 39788
rect 4080 36174 4108 39782
rect 4356 38010 4384 40054
rect 4344 38004 4396 38010
rect 4344 37946 4396 37952
rect 4540 37806 4568 46514
rect 4632 45558 4660 49778
rect 4620 45552 4672 45558
rect 4620 45494 4672 45500
rect 4724 45082 4752 53518
rect 4816 53038 4844 56200
rect 4896 54188 4948 54194
rect 4896 54130 4948 54136
rect 4804 53032 4856 53038
rect 4804 52974 4856 52980
rect 4908 52086 4936 54130
rect 5460 54126 5488 56200
rect 5448 54120 5500 54126
rect 5448 54062 5500 54068
rect 6104 53650 6132 56200
rect 6092 53644 6144 53650
rect 6092 53586 6144 53592
rect 5540 53576 5592 53582
rect 5540 53518 5592 53524
rect 4896 52080 4948 52086
rect 4896 52022 4948 52028
rect 5552 51542 5580 53518
rect 5816 53100 5868 53106
rect 5816 53042 5868 53048
rect 5828 52154 5856 53042
rect 6748 52562 6776 56200
rect 7392 55214 7420 56200
rect 8036 55214 8064 56200
rect 7392 55186 7604 55214
rect 7380 53576 7432 53582
rect 7380 53518 7432 53524
rect 6736 52556 6788 52562
rect 6736 52498 6788 52504
rect 5816 52148 5868 52154
rect 5816 52090 5868 52096
rect 7392 51610 7420 53518
rect 7576 53038 7604 55186
rect 7852 55186 8064 55214
rect 7748 54188 7800 54194
rect 7748 54130 7800 54136
rect 7564 53032 7616 53038
rect 7564 52974 7616 52980
rect 7380 51604 7432 51610
rect 7380 51546 7432 51552
rect 5540 51536 5592 51542
rect 5540 51478 5592 51484
rect 5172 51400 5224 51406
rect 5172 51342 5224 51348
rect 5184 46714 5212 51342
rect 7760 51066 7788 54130
rect 7852 53650 7880 55186
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 8680 54262 8708 56200
rect 8668 54256 8720 54262
rect 8668 54198 8720 54204
rect 7840 53644 7892 53650
rect 7840 53586 7892 53592
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 9036 53100 9088 53106
rect 9036 53042 9088 53048
rect 8484 52624 8536 52630
rect 8484 52566 8536 52572
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 8392 52012 8444 52018
rect 8392 51954 8444 51960
rect 7840 51400 7892 51406
rect 7840 51342 7892 51348
rect 7748 51060 7800 51066
rect 7748 51002 7800 51008
rect 7656 50924 7708 50930
rect 7656 50866 7708 50872
rect 5356 49768 5408 49774
rect 5356 49710 5408 49716
rect 5172 46708 5224 46714
rect 5172 46650 5224 46656
rect 4712 45076 4764 45082
rect 4712 45018 4764 45024
rect 4988 44804 5040 44810
rect 4988 44746 5040 44752
rect 4620 39432 4672 39438
rect 4620 39374 4672 39380
rect 4632 38554 4660 39374
rect 5000 38894 5028 44746
rect 5368 43314 5396 49710
rect 5448 45892 5500 45898
rect 5448 45834 5500 45840
rect 5460 45082 5488 45834
rect 5724 45484 5776 45490
rect 5724 45426 5776 45432
rect 6828 45484 6880 45490
rect 6828 45426 6880 45432
rect 5448 45076 5500 45082
rect 5448 45018 5500 45024
rect 5356 43308 5408 43314
rect 5356 43250 5408 43256
rect 5080 43240 5132 43246
rect 5080 43182 5132 43188
rect 4988 38888 5040 38894
rect 4988 38830 5040 38836
rect 4620 38548 4672 38554
rect 4620 38490 4672 38496
rect 4528 37800 4580 37806
rect 4528 37742 4580 37748
rect 4896 37800 4948 37806
rect 4896 37742 4948 37748
rect 4712 36576 4764 36582
rect 4712 36518 4764 36524
rect 4068 36168 4120 36174
rect 4068 36110 4120 36116
rect 3976 35080 4028 35086
rect 3976 35022 4028 35028
rect 4724 32910 4752 36518
rect 4804 35556 4856 35562
rect 4804 35498 4856 35504
rect 4712 32904 4764 32910
rect 4712 32846 4764 32852
rect 3516 23724 3568 23730
rect 3516 23666 3568 23672
rect 3424 22092 3476 22098
rect 3424 22034 3476 22040
rect 4816 21554 4844 35498
rect 4908 24818 4936 37742
rect 5000 25362 5028 38830
rect 5092 36854 5120 43182
rect 5460 39438 5488 45018
rect 5632 44804 5684 44810
rect 5632 44746 5684 44752
rect 5540 44736 5592 44742
rect 5540 44678 5592 44684
rect 5552 44470 5580 44678
rect 5540 44464 5592 44470
rect 5540 44406 5592 44412
rect 5644 42702 5672 44746
rect 5632 42696 5684 42702
rect 5632 42638 5684 42644
rect 5540 41472 5592 41478
rect 5540 41414 5592 41420
rect 5448 39432 5500 39438
rect 5448 39374 5500 39380
rect 5264 38956 5316 38962
rect 5264 38898 5316 38904
rect 5276 38554 5304 38898
rect 5356 38752 5408 38758
rect 5356 38694 5408 38700
rect 5264 38548 5316 38554
rect 5264 38490 5316 38496
rect 5080 36848 5132 36854
rect 5080 36790 5132 36796
rect 5368 35698 5396 38694
rect 5552 38418 5580 41414
rect 5736 39098 5764 45426
rect 6184 45416 6236 45422
rect 6184 45358 6236 45364
rect 5816 44872 5868 44878
rect 5816 44814 5868 44820
rect 5828 43994 5856 44814
rect 5816 43988 5868 43994
rect 5816 43930 5868 43936
rect 5828 41414 5856 43930
rect 6000 42696 6052 42702
rect 6000 42638 6052 42644
rect 5828 41386 5948 41414
rect 5816 39296 5868 39302
rect 5816 39238 5868 39244
rect 5724 39092 5776 39098
rect 5724 39034 5776 39040
rect 5632 38820 5684 38826
rect 5632 38762 5684 38768
rect 5540 38412 5592 38418
rect 5540 38354 5592 38360
rect 5448 38208 5500 38214
rect 5448 38150 5500 38156
rect 5460 37806 5488 38150
rect 5448 37800 5500 37806
rect 5448 37742 5500 37748
rect 5644 37330 5672 38762
rect 5724 38548 5776 38554
rect 5724 38490 5776 38496
rect 5736 37942 5764 38490
rect 5724 37936 5776 37942
rect 5724 37878 5776 37884
rect 5632 37324 5684 37330
rect 5632 37266 5684 37272
rect 5540 37120 5592 37126
rect 5828 37108 5856 39238
rect 5920 38350 5948 41386
rect 5908 38344 5960 38350
rect 5908 38286 5960 38292
rect 5920 38010 5948 38286
rect 5908 38004 5960 38010
rect 5908 37946 5960 37952
rect 5908 37800 5960 37806
rect 5908 37742 5960 37748
rect 5920 37466 5948 37742
rect 5908 37460 5960 37466
rect 5908 37402 5960 37408
rect 5828 37080 5948 37108
rect 5540 37062 5592 37068
rect 5552 36378 5580 37062
rect 5816 36576 5868 36582
rect 5816 36518 5868 36524
rect 5540 36372 5592 36378
rect 5540 36314 5592 36320
rect 5724 36032 5776 36038
rect 5724 35974 5776 35980
rect 5736 35834 5764 35974
rect 5724 35828 5776 35834
rect 5724 35770 5776 35776
rect 5356 35692 5408 35698
rect 5356 35634 5408 35640
rect 5828 35086 5856 36518
rect 5920 35154 5948 37080
rect 6012 35766 6040 42638
rect 6092 38752 6144 38758
rect 6092 38694 6144 38700
rect 6000 35760 6052 35766
rect 6000 35702 6052 35708
rect 5908 35148 5960 35154
rect 5908 35090 5960 35096
rect 5816 35080 5868 35086
rect 5816 35022 5868 35028
rect 6104 33522 6132 38694
rect 6196 36922 6224 45358
rect 6368 44736 6420 44742
rect 6368 44678 6420 44684
rect 6274 37360 6330 37369
rect 6274 37295 6330 37304
rect 6184 36916 6236 36922
rect 6184 36858 6236 36864
rect 6288 36106 6316 37295
rect 6380 36174 6408 44678
rect 6840 44538 6868 45426
rect 7668 45354 7696 50866
rect 7852 46170 7880 51342
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 8404 47530 8432 51954
rect 8392 47524 8444 47530
rect 8392 47466 8444 47472
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 7840 46164 7892 46170
rect 7840 46106 7892 46112
rect 7748 45960 7800 45966
rect 7748 45902 7800 45908
rect 7656 45348 7708 45354
rect 7656 45290 7708 45296
rect 7012 45280 7064 45286
rect 7012 45222 7064 45228
rect 6828 44532 6880 44538
rect 6828 44474 6880 44480
rect 7024 43790 7052 45222
rect 7288 43852 7340 43858
rect 7288 43794 7340 43800
rect 7012 43784 7064 43790
rect 7012 43726 7064 43732
rect 7012 42560 7064 42566
rect 7012 42502 7064 42508
rect 7024 41614 7052 42502
rect 7104 42084 7156 42090
rect 7104 42026 7156 42032
rect 7012 41608 7064 41614
rect 7012 41550 7064 41556
rect 6920 40996 6972 41002
rect 6920 40938 6972 40944
rect 6552 39500 6604 39506
rect 6552 39442 6604 39448
rect 6460 38888 6512 38894
rect 6460 38830 6512 38836
rect 6472 36242 6500 38830
rect 6564 36718 6592 39442
rect 6932 38554 6960 40938
rect 6920 38548 6972 38554
rect 6920 38490 6972 38496
rect 6736 38412 6788 38418
rect 6736 38354 6788 38360
rect 6644 38208 6696 38214
rect 6644 38150 6696 38156
rect 6656 37330 6684 38150
rect 6748 37618 6776 38354
rect 6828 38344 6880 38350
rect 6880 38292 6960 38298
rect 6828 38286 6960 38292
rect 6840 38270 6960 38286
rect 6828 37800 6880 37806
rect 6932 37754 6960 38270
rect 6880 37748 6960 37754
rect 6828 37742 6960 37748
rect 6840 37726 6960 37742
rect 6748 37590 6868 37618
rect 6644 37324 6696 37330
rect 6644 37266 6696 37272
rect 6552 36712 6604 36718
rect 6552 36654 6604 36660
rect 6564 36310 6592 36654
rect 6552 36304 6604 36310
rect 6552 36246 6604 36252
rect 6460 36236 6512 36242
rect 6460 36178 6512 36184
rect 6368 36168 6420 36174
rect 6368 36110 6420 36116
rect 6276 36100 6328 36106
rect 6276 36042 6328 36048
rect 6460 36100 6512 36106
rect 6460 36042 6512 36048
rect 6092 33516 6144 33522
rect 6092 33458 6144 33464
rect 5632 33312 5684 33318
rect 5632 33254 5684 33260
rect 5448 32836 5500 32842
rect 5448 32778 5500 32784
rect 5460 32502 5488 32778
rect 5540 32768 5592 32774
rect 5540 32710 5592 32716
rect 5448 32496 5500 32502
rect 5448 32438 5500 32444
rect 5552 31346 5580 32710
rect 5644 31822 5672 33254
rect 5632 31816 5684 31822
rect 5632 31758 5684 31764
rect 6288 31754 6316 36042
rect 5920 31726 6316 31754
rect 5540 31340 5592 31346
rect 5540 31282 5592 31288
rect 4988 25356 5040 25362
rect 4988 25298 5040 25304
rect 4896 24812 4948 24818
rect 4896 24754 4948 24760
rect 5920 23186 5948 31726
rect 6472 27062 6500 36042
rect 6564 35630 6592 36246
rect 6656 36174 6684 37266
rect 6736 37120 6788 37126
rect 6736 37062 6788 37068
rect 6748 36854 6776 37062
rect 6736 36848 6788 36854
rect 6736 36790 6788 36796
rect 6840 36786 6868 37590
rect 6828 36780 6880 36786
rect 6828 36722 6880 36728
rect 6932 36174 6960 37726
rect 6644 36168 6696 36174
rect 6644 36110 6696 36116
rect 6920 36168 6972 36174
rect 6920 36110 6972 36116
rect 7024 36106 7052 41550
rect 7116 36922 7144 42026
rect 7300 39030 7328 43794
rect 7656 43784 7708 43790
rect 7656 43726 7708 43732
rect 7472 43648 7524 43654
rect 7472 43590 7524 43596
rect 7288 39024 7340 39030
rect 7288 38966 7340 38972
rect 7196 38888 7248 38894
rect 7196 38830 7248 38836
rect 7208 37194 7236 38830
rect 7380 38276 7432 38282
rect 7380 38218 7432 38224
rect 7288 38004 7340 38010
rect 7288 37946 7340 37952
rect 7196 37188 7248 37194
rect 7196 37130 7248 37136
rect 7104 36916 7156 36922
rect 7104 36858 7156 36864
rect 7104 36712 7156 36718
rect 7102 36680 7104 36689
rect 7156 36680 7158 36689
rect 7102 36615 7158 36624
rect 7104 36236 7156 36242
rect 7104 36178 7156 36184
rect 7012 36100 7064 36106
rect 7012 36042 7064 36048
rect 6828 36032 6880 36038
rect 6828 35974 6880 35980
rect 6552 35624 6604 35630
rect 6552 35566 6604 35572
rect 6564 33930 6592 35566
rect 6736 35488 6788 35494
rect 6736 35430 6788 35436
rect 6748 35154 6776 35430
rect 6736 35148 6788 35154
rect 6736 35090 6788 35096
rect 6644 34672 6696 34678
rect 6644 34614 6696 34620
rect 6552 33924 6604 33930
rect 6552 33866 6604 33872
rect 6656 33590 6684 34614
rect 6840 33590 6868 35974
rect 6920 34944 6972 34950
rect 6920 34886 6972 34892
rect 7012 34944 7064 34950
rect 7012 34886 7064 34892
rect 6644 33584 6696 33590
rect 6644 33526 6696 33532
rect 6828 33584 6880 33590
rect 6828 33526 6880 33532
rect 6932 32910 6960 34886
rect 6920 32904 6972 32910
rect 6920 32846 6972 32852
rect 6920 32292 6972 32298
rect 6920 32234 6972 32240
rect 6932 31890 6960 32234
rect 6920 31884 6972 31890
rect 6920 31826 6972 31832
rect 6460 27056 6512 27062
rect 6460 26998 6512 27004
rect 7024 26234 7052 34886
rect 7116 34406 7144 36178
rect 7196 35148 7248 35154
rect 7196 35090 7248 35096
rect 7208 35018 7236 35090
rect 7196 35012 7248 35018
rect 7196 34954 7248 34960
rect 7104 34400 7156 34406
rect 7104 34342 7156 34348
rect 7208 34202 7236 34954
rect 7300 34610 7328 37946
rect 7392 37505 7420 38218
rect 7484 38010 7512 43590
rect 7564 42628 7616 42634
rect 7564 42570 7616 42576
rect 7576 39642 7604 42570
rect 7564 39636 7616 39642
rect 7564 39578 7616 39584
rect 7472 38004 7524 38010
rect 7472 37946 7524 37952
rect 7378 37496 7434 37505
rect 7378 37431 7434 37440
rect 7380 37324 7432 37330
rect 7380 37266 7432 37272
rect 7392 36922 7420 37266
rect 7668 37262 7696 43726
rect 7760 40730 7788 45902
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 8496 42566 8524 52566
rect 9048 51066 9076 53042
rect 9324 52562 9352 56200
rect 9968 55214 9996 56200
rect 9968 55186 10088 55214
rect 9956 53100 10008 53106
rect 9956 53042 10008 53048
rect 9312 52556 9364 52562
rect 9312 52498 9364 52504
rect 9220 52488 9272 52494
rect 9220 52430 9272 52436
rect 9680 52488 9732 52494
rect 9680 52430 9732 52436
rect 9232 51610 9260 52430
rect 9692 52154 9720 52430
rect 9968 52154 9996 53042
rect 10060 53038 10088 55186
rect 10416 54732 10468 54738
rect 10416 54674 10468 54680
rect 10048 53032 10100 53038
rect 10048 52974 10100 52980
rect 9680 52148 9732 52154
rect 9680 52090 9732 52096
rect 9956 52148 10008 52154
rect 9956 52090 10008 52096
rect 9864 52012 9916 52018
rect 9864 51954 9916 51960
rect 9220 51604 9272 51610
rect 9220 51546 9272 51552
rect 9036 51060 9088 51066
rect 9036 51002 9088 51008
rect 9220 50924 9272 50930
rect 9220 50866 9272 50872
rect 9232 48890 9260 50866
rect 9772 49156 9824 49162
rect 9772 49098 9824 49104
rect 9220 48884 9272 48890
rect 9220 48826 9272 48832
rect 8760 47184 8812 47190
rect 8760 47126 8812 47132
rect 8772 44402 8800 47126
rect 9588 46572 9640 46578
rect 9588 46514 9640 46520
rect 9128 45484 9180 45490
rect 9128 45426 9180 45432
rect 8760 44396 8812 44402
rect 8760 44338 8812 44344
rect 8944 42900 8996 42906
rect 8944 42842 8996 42848
rect 8760 42628 8812 42634
rect 8760 42570 8812 42576
rect 8484 42560 8536 42566
rect 8484 42502 8536 42508
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 8496 42022 8524 42502
rect 8772 42226 8800 42570
rect 8760 42220 8812 42226
rect 8760 42162 8812 42168
rect 8772 42106 8800 42162
rect 8588 42078 8800 42106
rect 8484 42016 8536 42022
rect 8484 41958 8536 41964
rect 8300 41608 8352 41614
rect 8300 41550 8352 41556
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 7840 41132 7892 41138
rect 7840 41074 7892 41080
rect 7748 40724 7800 40730
rect 7748 40666 7800 40672
rect 7748 40384 7800 40390
rect 7748 40326 7800 40332
rect 7656 37256 7708 37262
rect 7656 37198 7708 37204
rect 7472 37188 7524 37194
rect 7472 37130 7524 37136
rect 7380 36916 7432 36922
rect 7380 36858 7432 36864
rect 7484 36825 7512 37130
rect 7564 37120 7616 37126
rect 7564 37062 7616 37068
rect 7470 36816 7526 36825
rect 7380 36780 7432 36786
rect 7470 36751 7526 36760
rect 7380 36722 7432 36728
rect 7392 36106 7420 36722
rect 7484 36650 7512 36751
rect 7472 36644 7524 36650
rect 7472 36586 7524 36592
rect 7380 36100 7432 36106
rect 7380 36042 7432 36048
rect 7288 34604 7340 34610
rect 7288 34546 7340 34552
rect 7288 34468 7340 34474
rect 7288 34410 7340 34416
rect 7196 34196 7248 34202
rect 7196 34138 7248 34144
rect 7104 33924 7156 33930
rect 7104 33866 7156 33872
rect 7116 31686 7144 33866
rect 7196 33652 7248 33658
rect 7196 33594 7248 33600
rect 7104 31680 7156 31686
rect 7104 31622 7156 31628
rect 7208 26234 7236 33594
rect 6932 26206 7052 26234
rect 7116 26206 7236 26234
rect 7300 26234 7328 34410
rect 7392 33658 7420 36042
rect 7576 35698 7604 37062
rect 7656 36916 7708 36922
rect 7656 36858 7708 36864
rect 7668 36718 7696 36858
rect 7656 36712 7708 36718
rect 7656 36654 7708 36660
rect 7668 36106 7696 36654
rect 7656 36100 7708 36106
rect 7656 36042 7708 36048
rect 7668 35714 7696 36042
rect 7760 35834 7788 40326
rect 7852 37194 7880 41074
rect 8208 40928 8260 40934
rect 8208 40870 8260 40876
rect 8220 40372 8248 40870
rect 8312 40526 8340 41550
rect 8484 41132 8536 41138
rect 8484 41074 8536 41080
rect 8496 40526 8524 41074
rect 8588 41070 8616 42078
rect 8668 42016 8720 42022
rect 8668 41958 8720 41964
rect 8576 41064 8628 41070
rect 8576 41006 8628 41012
rect 8300 40520 8352 40526
rect 8300 40462 8352 40468
rect 8484 40520 8536 40526
rect 8484 40462 8536 40468
rect 8392 40384 8444 40390
rect 8220 40344 8340 40372
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 8312 40118 8340 40344
rect 8392 40326 8444 40332
rect 8300 40112 8352 40118
rect 8300 40054 8352 40060
rect 8404 39982 8432 40326
rect 8496 40050 8524 40462
rect 8484 40044 8536 40050
rect 8484 39986 8536 39992
rect 8392 39976 8444 39982
rect 8392 39918 8444 39924
rect 8208 39636 8260 39642
rect 8208 39578 8260 39584
rect 8220 39438 8248 39578
rect 8484 39500 8536 39506
rect 8588 39488 8616 41006
rect 8680 39506 8708 41958
rect 8760 40452 8812 40458
rect 8760 40394 8812 40400
rect 8536 39460 8616 39488
rect 8668 39500 8720 39506
rect 8484 39442 8536 39448
rect 8668 39442 8720 39448
rect 8208 39432 8260 39438
rect 8208 39374 8260 39380
rect 8220 39284 8248 39374
rect 8220 39256 8340 39284
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 8208 39024 8260 39030
rect 8312 39012 8340 39256
rect 8260 38984 8340 39012
rect 8208 38966 8260 38972
rect 8220 38350 8248 38966
rect 8496 38962 8524 39442
rect 8668 39364 8720 39370
rect 8668 39306 8720 39312
rect 8576 39296 8628 39302
rect 8576 39238 8628 39244
rect 8484 38956 8536 38962
rect 8484 38898 8536 38904
rect 8484 38820 8536 38826
rect 8484 38762 8536 38768
rect 8300 38480 8352 38486
rect 8300 38422 8352 38428
rect 8208 38344 8260 38350
rect 8208 38286 8260 38292
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 8208 37868 8260 37874
rect 8208 37810 8260 37816
rect 8116 37732 8168 37738
rect 8116 37674 8168 37680
rect 8128 37618 8156 37674
rect 8036 37590 8156 37618
rect 8036 37398 8064 37590
rect 8024 37392 8076 37398
rect 8024 37334 8076 37340
rect 7840 37188 7892 37194
rect 7840 37130 7892 37136
rect 8220 37126 8248 37810
rect 8312 37806 8340 38422
rect 8392 38344 8444 38350
rect 8392 38286 8444 38292
rect 8404 37874 8432 38286
rect 8392 37868 8444 37874
rect 8392 37810 8444 37816
rect 8300 37800 8352 37806
rect 8300 37742 8352 37748
rect 8392 37664 8444 37670
rect 8392 37606 8444 37612
rect 8300 37460 8352 37466
rect 8300 37402 8352 37408
rect 8208 37120 8260 37126
rect 8208 37062 8260 37068
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 8312 36904 8340 37402
rect 8404 36922 8432 37606
rect 8220 36876 8340 36904
rect 8392 36916 8444 36922
rect 8220 36689 8248 36876
rect 8392 36858 8444 36864
rect 8206 36680 8262 36689
rect 8206 36615 8262 36624
rect 7932 36576 7984 36582
rect 7932 36518 7984 36524
rect 8300 36576 8352 36582
rect 8300 36518 8352 36524
rect 7944 36242 7972 36518
rect 7932 36236 7984 36242
rect 7932 36178 7984 36184
rect 7932 36032 7984 36038
rect 7852 35992 7932 36020
rect 7748 35828 7800 35834
rect 7748 35770 7800 35776
rect 7564 35692 7616 35698
rect 7668 35686 7788 35714
rect 7564 35634 7616 35640
rect 7472 35624 7524 35630
rect 7472 35566 7524 35572
rect 7380 33652 7432 33658
rect 7380 33594 7432 33600
rect 7484 33454 7512 35566
rect 7656 35216 7708 35222
rect 7656 35158 7708 35164
rect 7564 34400 7616 34406
rect 7564 34342 7616 34348
rect 7576 33658 7604 34342
rect 7564 33652 7616 33658
rect 7564 33594 7616 33600
rect 7472 33448 7524 33454
rect 7472 33390 7524 33396
rect 7564 33108 7616 33114
rect 7564 33050 7616 33056
rect 7472 32292 7524 32298
rect 7472 32234 7524 32240
rect 7484 28694 7512 32234
rect 7472 28688 7524 28694
rect 7472 28630 7524 28636
rect 7576 28626 7604 33050
rect 7668 32842 7696 35158
rect 7760 35154 7788 35686
rect 7852 35290 7880 35992
rect 7932 35974 7984 35980
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 7840 35284 7892 35290
rect 7840 35226 7892 35232
rect 8208 35216 8260 35222
rect 8208 35158 8260 35164
rect 7748 35148 7800 35154
rect 7748 35090 7800 35096
rect 7760 34134 7788 35090
rect 8114 35048 8170 35057
rect 8114 34983 8116 34992
rect 8168 34983 8170 34992
rect 8116 34954 8168 34960
rect 8220 34950 8248 35158
rect 8312 35086 8340 36518
rect 8496 36242 8524 38762
rect 8588 38010 8616 39238
rect 8576 38004 8628 38010
rect 8576 37946 8628 37952
rect 8484 36236 8536 36242
rect 8484 36178 8536 36184
rect 8484 35760 8536 35766
rect 8484 35702 8536 35708
rect 8300 35080 8352 35086
rect 8300 35022 8352 35028
rect 8208 34944 8260 34950
rect 8208 34886 8260 34892
rect 8392 34944 8444 34950
rect 8392 34886 8444 34892
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 8404 34746 8432 34886
rect 8392 34740 8444 34746
rect 8392 34682 8444 34688
rect 8208 34468 8260 34474
rect 8208 34410 8260 34416
rect 7840 34196 7892 34202
rect 7840 34138 7892 34144
rect 7748 34128 7800 34134
rect 7748 34070 7800 34076
rect 7748 32972 7800 32978
rect 7748 32914 7800 32920
rect 7656 32836 7708 32842
rect 7656 32778 7708 32784
rect 7656 32224 7708 32230
rect 7656 32166 7708 32172
rect 7668 30734 7696 32166
rect 7760 31686 7788 32914
rect 7852 32298 7880 34138
rect 8220 33844 8248 34410
rect 8220 33816 8340 33844
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 8312 33386 8340 33816
rect 8300 33380 8352 33386
rect 8300 33322 8352 33328
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 7840 32292 7892 32298
rect 7840 32234 7892 32240
rect 7748 31680 7800 31686
rect 7748 31622 7800 31628
rect 7760 30870 7788 31622
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 8392 31272 8444 31278
rect 8392 31214 8444 31220
rect 7748 30864 7800 30870
rect 7748 30806 7800 30812
rect 7656 30728 7708 30734
rect 7656 30670 7708 30676
rect 7760 29238 7788 30806
rect 7840 30796 7892 30802
rect 7840 30738 7892 30744
rect 7748 29232 7800 29238
rect 7748 29174 7800 29180
rect 7852 28762 7880 30738
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 8404 30054 8432 31214
rect 8392 30048 8444 30054
rect 8392 29990 8444 29996
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 8404 29306 8432 29990
rect 8392 29300 8444 29306
rect 8392 29242 8444 29248
rect 8208 28960 8260 28966
rect 8208 28902 8260 28908
rect 7840 28756 7892 28762
rect 7840 28698 7892 28704
rect 7564 28620 7616 28626
rect 7564 28562 7616 28568
rect 8220 28558 8248 28902
rect 7748 28552 7800 28558
rect 7748 28494 7800 28500
rect 8208 28552 8260 28558
rect 8208 28494 8260 28500
rect 7300 26206 7696 26234
rect 5908 23180 5960 23186
rect 5908 23122 5960 23128
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 1858 20360 1914 20369
rect 1858 20295 1914 20304
rect 1872 19990 1900 20295
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 1860 19984 1912 19990
rect 1860 19926 1912 19932
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1780 17921 1808 18226
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 1766 17912 1822 17921
rect 2950 17915 3258 17924
rect 1766 17847 1822 17856
rect 1950 17776 2006 17785
rect 1950 17711 2006 17720
rect 1860 17128 1912 17134
rect 1858 17096 1860 17105
rect 1912 17096 1914 17105
rect 1858 17031 1914 17040
rect 1964 16726 1992 17711
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 1952 16720 2004 16726
rect 1952 16662 2004 16668
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 6932 15026 6960 26206
rect 7116 20466 7144 26206
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7668 15638 7696 26206
rect 7656 15632 7708 15638
rect 7656 15574 7708 15580
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 940 8968 992 8974
rect 938 8936 940 8945
rect 992 8936 994 8945
rect 938 8871 994 8880
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1780 8129 1808 8434
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 1766 8120 1822 8129
rect 2950 8123 3258 8132
rect 1766 8055 1822 8064
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 940 7404 992 7410
rect 940 7346 992 7352
rect 952 7313 980 7346
rect 938 7304 994 7313
rect 938 7239 994 7248
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 940 6724 992 6730
rect 940 6666 992 6672
rect 952 6497 980 6666
rect 938 6488 994 6497
rect 938 6423 994 6432
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 938 5672 994 5681
rect 938 5607 940 5616
rect 992 5607 994 5616
rect 940 5578 992 5584
rect 940 5228 992 5234
rect 940 5170 992 5176
rect 952 4865 980 5170
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 938 4856 994 4865
rect 2950 4859 3258 4868
rect 938 4791 994 4800
rect 940 4072 992 4078
rect 938 4040 940 4049
rect 992 4040 994 4049
rect 938 3975 994 3984
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 940 3528 992 3534
rect 940 3470 992 3476
rect 952 3233 980 3470
rect 938 3224 994 3233
rect 938 3159 994 3168
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2240 800 2268 2382
rect 5552 800 5580 2450
rect 6932 2446 6960 8026
rect 7760 6866 7788 28494
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 8496 26234 8524 35702
rect 8588 35630 8616 37946
rect 8680 37262 8708 39306
rect 8668 37256 8720 37262
rect 8668 37198 8720 37204
rect 8668 36712 8720 36718
rect 8668 36654 8720 36660
rect 8680 35630 8708 36654
rect 8576 35624 8628 35630
rect 8576 35566 8628 35572
rect 8668 35624 8720 35630
rect 8668 35566 8720 35572
rect 8772 34746 8800 40394
rect 8852 40180 8904 40186
rect 8852 40122 8904 40128
rect 8864 38418 8892 40122
rect 8956 38758 8984 42842
rect 9036 42152 9088 42158
rect 9036 42094 9088 42100
rect 9048 40594 9076 42094
rect 9140 40730 9168 45426
rect 9404 44192 9456 44198
rect 9404 44134 9456 44140
rect 9220 43308 9272 43314
rect 9220 43250 9272 43256
rect 9232 43217 9260 43250
rect 9218 43208 9274 43217
rect 9218 43143 9274 43152
rect 9220 43104 9272 43110
rect 9220 43046 9272 43052
rect 9232 41206 9260 43046
rect 9312 42696 9364 42702
rect 9312 42638 9364 42644
rect 9324 42362 9352 42638
rect 9312 42356 9364 42362
rect 9312 42298 9364 42304
rect 9416 41682 9444 44134
rect 9600 43110 9628 46514
rect 9680 43920 9732 43926
rect 9680 43862 9732 43868
rect 9588 43104 9640 43110
rect 9588 43046 9640 43052
rect 9404 41676 9456 41682
rect 9404 41618 9456 41624
rect 9220 41200 9272 41206
rect 9220 41142 9272 41148
rect 9128 40724 9180 40730
rect 9128 40666 9180 40672
rect 9036 40588 9088 40594
rect 9036 40530 9088 40536
rect 9312 40588 9364 40594
rect 9312 40530 9364 40536
rect 9048 39642 9076 40530
rect 9036 39636 9088 39642
rect 9036 39578 9088 39584
rect 9036 39432 9088 39438
rect 9036 39374 9088 39380
rect 8944 38752 8996 38758
rect 8944 38694 8996 38700
rect 8852 38412 8904 38418
rect 8852 38354 8904 38360
rect 8852 38208 8904 38214
rect 8852 38150 8904 38156
rect 8760 34740 8812 34746
rect 8760 34682 8812 34688
rect 8668 34604 8720 34610
rect 8668 34546 8720 34552
rect 8404 26206 8524 26234
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 8404 18970 8432 26206
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 8680 18426 8708 34546
rect 8864 32570 8892 38150
rect 8944 38004 8996 38010
rect 8944 37946 8996 37952
rect 8956 36854 8984 37946
rect 9048 37369 9076 39374
rect 9128 39296 9180 39302
rect 9128 39238 9180 39244
rect 9140 38894 9168 39238
rect 9128 38888 9180 38894
rect 9128 38830 9180 38836
rect 9126 38720 9182 38729
rect 9126 38655 9182 38664
rect 9034 37360 9090 37369
rect 9034 37295 9090 37304
rect 9036 37256 9088 37262
rect 9036 37198 9088 37204
rect 8944 36848 8996 36854
rect 8944 36790 8996 36796
rect 8944 36236 8996 36242
rect 8944 36178 8996 36184
rect 8852 32564 8904 32570
rect 8852 32506 8904 32512
rect 8956 32366 8984 36178
rect 9048 36174 9076 37198
rect 9140 36718 9168 38655
rect 9324 38486 9352 40530
rect 9496 39296 9548 39302
rect 9496 39238 9548 39244
rect 9508 38554 9536 39238
rect 9496 38548 9548 38554
rect 9496 38490 9548 38496
rect 9312 38480 9364 38486
rect 9312 38422 9364 38428
rect 9404 38412 9456 38418
rect 9404 38354 9456 38360
rect 9496 38412 9548 38418
rect 9496 38354 9548 38360
rect 9220 37664 9272 37670
rect 9220 37606 9272 37612
rect 9232 36922 9260 37606
rect 9310 37496 9366 37505
rect 9310 37431 9366 37440
rect 9220 36916 9272 36922
rect 9220 36858 9272 36864
rect 9128 36712 9180 36718
rect 9128 36654 9180 36660
rect 9036 36168 9088 36174
rect 9036 36110 9088 36116
rect 9048 34066 9076 36110
rect 9128 35488 9180 35494
rect 9128 35430 9180 35436
rect 9220 35488 9272 35494
rect 9220 35430 9272 35436
rect 9036 34060 9088 34066
rect 9036 34002 9088 34008
rect 9048 33522 9076 34002
rect 9036 33516 9088 33522
rect 9036 33458 9088 33464
rect 9140 32434 9168 35430
rect 9232 32910 9260 35430
rect 9324 35222 9352 37431
rect 9312 35216 9364 35222
rect 9312 35158 9364 35164
rect 9416 34474 9444 38354
rect 9508 37738 9536 38354
rect 9600 38010 9628 43046
rect 9588 38004 9640 38010
rect 9588 37946 9640 37952
rect 9496 37732 9548 37738
rect 9496 37674 9548 37680
rect 9692 37505 9720 43862
rect 9784 43450 9812 49098
rect 9876 47802 9904 51954
rect 9956 49428 10008 49434
rect 9956 49370 10008 49376
rect 9864 47796 9916 47802
rect 9864 47738 9916 47744
rect 9864 47660 9916 47666
rect 9864 47602 9916 47608
rect 9876 43450 9904 47602
rect 9968 44878 9996 49370
rect 9956 44872 10008 44878
rect 9956 44814 10008 44820
rect 10428 44470 10456 54674
rect 10612 54262 10640 56200
rect 10600 54256 10652 54262
rect 10600 54198 10652 54204
rect 10876 54188 10928 54194
rect 10876 54130 10928 54136
rect 10600 54120 10652 54126
rect 10600 54062 10652 54068
rect 10508 52012 10560 52018
rect 10508 51954 10560 51960
rect 10520 47802 10548 51954
rect 10508 47796 10560 47802
rect 10508 47738 10560 47744
rect 10612 46186 10640 54062
rect 10692 51944 10744 51950
rect 10692 51886 10744 51892
rect 10704 47802 10732 51886
rect 10888 51610 10916 54130
rect 11256 53650 11284 56200
rect 11612 54596 11664 54602
rect 11612 54538 11664 54544
rect 11244 53644 11296 53650
rect 11244 53586 11296 53592
rect 10876 51604 10928 51610
rect 10876 51546 10928 51552
rect 10968 51400 11020 51406
rect 10968 51342 11020 51348
rect 11060 51400 11112 51406
rect 11060 51342 11112 51348
rect 10784 51332 10836 51338
rect 10784 51274 10836 51280
rect 10692 47796 10744 47802
rect 10692 47738 10744 47744
rect 10796 47258 10824 51274
rect 10784 47252 10836 47258
rect 10784 47194 10836 47200
rect 10980 46714 11008 51342
rect 10968 46708 11020 46714
rect 10968 46650 11020 46656
rect 10612 46158 10732 46186
rect 11072 46170 11100 51342
rect 11624 51074 11652 54538
rect 11704 53576 11756 53582
rect 11704 53518 11756 53524
rect 11532 51046 11652 51074
rect 11244 48748 11296 48754
rect 11244 48690 11296 48696
rect 9956 44464 10008 44470
rect 9956 44406 10008 44412
rect 10416 44464 10468 44470
rect 10416 44406 10468 44412
rect 9772 43444 9824 43450
rect 9772 43386 9824 43392
rect 9864 43444 9916 43450
rect 9864 43386 9916 43392
rect 9772 43172 9824 43178
rect 9772 43114 9824 43120
rect 9784 41614 9812 43114
rect 9772 41608 9824 41614
rect 9772 41550 9824 41556
rect 9862 40488 9918 40497
rect 9862 40423 9918 40432
rect 9772 38752 9824 38758
rect 9772 38694 9824 38700
rect 9784 38418 9812 38694
rect 9772 38412 9824 38418
rect 9772 38354 9824 38360
rect 9876 38282 9904 40423
rect 9968 38282 9996 44406
rect 10232 44396 10284 44402
rect 10232 44338 10284 44344
rect 10048 43308 10100 43314
rect 10048 43250 10100 43256
rect 9864 38276 9916 38282
rect 9864 38218 9916 38224
rect 9956 38276 10008 38282
rect 9956 38218 10008 38224
rect 9772 38208 9824 38214
rect 9772 38150 9824 38156
rect 9678 37496 9734 37505
rect 9678 37431 9734 37440
rect 9680 37324 9732 37330
rect 9680 37266 9732 37272
rect 9496 37188 9548 37194
rect 9496 37130 9548 37136
rect 9404 34468 9456 34474
rect 9404 34410 9456 34416
rect 9220 32904 9272 32910
rect 9220 32846 9272 32852
rect 9312 32768 9364 32774
rect 9312 32710 9364 32716
rect 9218 32600 9274 32609
rect 9218 32535 9220 32544
rect 9272 32535 9274 32544
rect 9220 32506 9272 32512
rect 9128 32428 9180 32434
rect 9128 32370 9180 32376
rect 8944 32360 8996 32366
rect 8944 32302 8996 32308
rect 9036 30048 9088 30054
rect 9036 29990 9088 29996
rect 9048 29850 9076 29990
rect 9036 29844 9088 29850
rect 9036 29786 9088 29792
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 9232 5302 9260 32506
rect 9324 27062 9352 32710
rect 9508 30734 9536 37130
rect 9586 36952 9642 36961
rect 9586 36887 9588 36896
rect 9640 36887 9642 36896
rect 9588 36858 9640 36864
rect 9588 36712 9640 36718
rect 9586 36680 9588 36689
rect 9640 36680 9642 36689
rect 9586 36615 9642 36624
rect 9692 34950 9720 37266
rect 9784 35834 9812 38150
rect 9876 38010 9904 38218
rect 9864 38004 9916 38010
rect 9864 37946 9916 37952
rect 9864 37800 9916 37806
rect 9864 37742 9916 37748
rect 9876 37398 9904 37742
rect 9864 37392 9916 37398
rect 9864 37334 9916 37340
rect 9864 36644 9916 36650
rect 9864 36586 9916 36592
rect 9956 36644 10008 36650
rect 9956 36586 10008 36592
rect 9772 35828 9824 35834
rect 9772 35770 9824 35776
rect 9680 34944 9732 34950
rect 9680 34886 9732 34892
rect 9680 33856 9732 33862
rect 9680 33798 9732 33804
rect 9692 32570 9720 33798
rect 9772 33040 9824 33046
rect 9772 32982 9824 32988
rect 9680 32564 9732 32570
rect 9680 32506 9732 32512
rect 9784 31090 9812 32982
rect 9876 32910 9904 36586
rect 9968 34610 9996 36586
rect 10060 35834 10088 43250
rect 10244 41414 10272 44338
rect 10324 42628 10376 42634
rect 10376 42588 10548 42616
rect 10324 42570 10376 42576
rect 10416 42152 10468 42158
rect 10416 42094 10468 42100
rect 10428 41682 10456 42094
rect 10520 42090 10548 42588
rect 10508 42084 10560 42090
rect 10508 42026 10560 42032
rect 10416 41676 10468 41682
rect 10416 41618 10468 41624
rect 10244 41386 10364 41414
rect 10336 41274 10364 41386
rect 10324 41268 10376 41274
rect 10324 41210 10376 41216
rect 10428 40458 10456 41618
rect 10416 40452 10468 40458
rect 10416 40394 10468 40400
rect 10140 40112 10192 40118
rect 10140 40054 10192 40060
rect 10152 39098 10180 40054
rect 10520 39545 10548 42026
rect 10600 41540 10652 41546
rect 10600 41482 10652 41488
rect 10506 39536 10562 39545
rect 10506 39471 10562 39480
rect 10140 39092 10192 39098
rect 10140 39034 10192 39040
rect 10140 37800 10192 37806
rect 10140 37742 10192 37748
rect 10048 35828 10100 35834
rect 10048 35770 10100 35776
rect 10152 35766 10180 37742
rect 10232 37392 10284 37398
rect 10232 37334 10284 37340
rect 10140 35760 10192 35766
rect 10140 35702 10192 35708
rect 10244 35018 10272 37334
rect 10416 37120 10468 37126
rect 10416 37062 10468 37068
rect 10428 36106 10456 37062
rect 10612 36922 10640 41482
rect 10704 40934 10732 46158
rect 11060 46164 11112 46170
rect 11060 46106 11112 46112
rect 10876 45348 10928 45354
rect 10876 45290 10928 45296
rect 10784 44192 10836 44198
rect 10784 44134 10836 44140
rect 10796 43450 10824 44134
rect 10784 43444 10836 43450
rect 10784 43386 10836 43392
rect 10888 41818 10916 45290
rect 11256 43994 11284 48690
rect 11336 46436 11388 46442
rect 11336 46378 11388 46384
rect 11244 43988 11296 43994
rect 11244 43930 11296 43936
rect 11348 43790 11376 46378
rect 11428 45960 11480 45966
rect 11428 45902 11480 45908
rect 11336 43784 11388 43790
rect 11336 43726 11388 43732
rect 11440 43450 11468 45902
rect 11428 43444 11480 43450
rect 11428 43386 11480 43392
rect 10968 43240 11020 43246
rect 10968 43182 11020 43188
rect 10876 41812 10928 41818
rect 10876 41754 10928 41760
rect 10980 41414 11008 43182
rect 11532 43178 11560 51046
rect 11716 50522 11744 53518
rect 11900 52562 11928 56200
rect 12544 55214 12572 56200
rect 12452 55186 12572 55214
rect 13188 55214 13216 56200
rect 13188 55186 13400 55214
rect 12348 53576 12400 53582
rect 12348 53518 12400 53524
rect 12164 53100 12216 53106
rect 12164 53042 12216 53048
rect 11888 52556 11940 52562
rect 11888 52498 11940 52504
rect 11796 52488 11848 52494
rect 11796 52430 11848 52436
rect 11704 50516 11756 50522
rect 11704 50458 11756 50464
rect 11808 49366 11836 52430
rect 11888 50312 11940 50318
rect 11888 50254 11940 50260
rect 11796 49360 11848 49366
rect 11796 49302 11848 49308
rect 11612 47728 11664 47734
rect 11612 47670 11664 47676
rect 11520 43172 11572 43178
rect 11440 43132 11520 43160
rect 11336 42628 11388 42634
rect 11336 42570 11388 42576
rect 11348 42344 11376 42570
rect 11072 42316 11376 42344
rect 11072 42226 11100 42316
rect 11060 42220 11112 42226
rect 11060 42162 11112 42168
rect 11152 42220 11204 42226
rect 11152 42162 11204 42168
rect 11164 41818 11192 42162
rect 11152 41812 11204 41818
rect 11152 41754 11204 41760
rect 10888 41386 11008 41414
rect 10782 41032 10838 41041
rect 10782 40967 10838 40976
rect 10692 40928 10744 40934
rect 10690 40896 10692 40905
rect 10744 40896 10746 40905
rect 10690 40831 10746 40840
rect 10692 40724 10744 40730
rect 10692 40666 10744 40672
rect 10704 38196 10732 40666
rect 10796 39642 10824 40967
rect 10888 40934 10916 41386
rect 11348 41206 11376 42316
rect 11336 41200 11388 41206
rect 11256 41160 11336 41188
rect 10876 40928 10928 40934
rect 10876 40870 10928 40876
rect 10888 39982 10916 40870
rect 11256 40458 11284 41160
rect 11336 41142 11388 41148
rect 11336 40996 11388 41002
rect 11336 40938 11388 40944
rect 11244 40452 11296 40458
rect 11244 40394 11296 40400
rect 11256 40186 11284 40394
rect 11244 40180 11296 40186
rect 11244 40122 11296 40128
rect 10966 40080 11022 40089
rect 10966 40015 11022 40024
rect 10876 39976 10928 39982
rect 10876 39918 10928 39924
rect 10784 39636 10836 39642
rect 10784 39578 10836 39584
rect 10980 38418 11008 40015
rect 11244 39500 11296 39506
rect 11244 39442 11296 39448
rect 11152 38820 11204 38826
rect 11152 38762 11204 38768
rect 10968 38412 11020 38418
rect 10968 38354 11020 38360
rect 10876 38208 10928 38214
rect 10704 38176 10876 38196
rect 10928 38176 10930 38185
rect 10704 38168 10874 38176
rect 10874 38111 10930 38120
rect 10980 37942 11008 38354
rect 11060 38208 11112 38214
rect 11060 38150 11112 38156
rect 10968 37936 11020 37942
rect 10968 37878 11020 37884
rect 11072 37466 11100 38150
rect 11060 37460 11112 37466
rect 11060 37402 11112 37408
rect 11060 37256 11112 37262
rect 11058 37224 11060 37233
rect 11112 37224 11114 37233
rect 11058 37159 11114 37168
rect 10600 36916 10652 36922
rect 10600 36858 10652 36864
rect 10600 36712 10652 36718
rect 10600 36654 10652 36660
rect 10612 36378 10640 36654
rect 10600 36372 10652 36378
rect 10600 36314 10652 36320
rect 10416 36100 10468 36106
rect 10416 36042 10468 36048
rect 10428 35018 10456 36042
rect 10508 35624 10560 35630
rect 10508 35566 10560 35572
rect 10520 35290 10548 35566
rect 10508 35284 10560 35290
rect 10508 35226 10560 35232
rect 10232 35012 10284 35018
rect 10416 35012 10468 35018
rect 10284 34972 10364 35000
rect 10232 34954 10284 34960
rect 9956 34604 10008 34610
rect 9956 34546 10008 34552
rect 10232 34536 10284 34542
rect 10232 34478 10284 34484
rect 9956 34400 10008 34406
rect 9956 34342 10008 34348
rect 10048 34400 10100 34406
rect 10048 34342 10100 34348
rect 9864 32904 9916 32910
rect 9864 32846 9916 32852
rect 9784 31062 9904 31090
rect 9772 30932 9824 30938
rect 9772 30874 9824 30880
rect 9496 30728 9548 30734
rect 9496 30670 9548 30676
rect 9588 30252 9640 30258
rect 9588 30194 9640 30200
rect 9600 29306 9628 30194
rect 9680 30184 9732 30190
rect 9680 30126 9732 30132
rect 9588 29300 9640 29306
rect 9588 29242 9640 29248
rect 9404 27872 9456 27878
rect 9404 27814 9456 27820
rect 9312 27056 9364 27062
rect 9312 26998 9364 27004
rect 9416 20942 9444 27814
rect 9404 20936 9456 20942
rect 9404 20878 9456 20884
rect 9600 7954 9628 29242
rect 9692 29102 9720 30126
rect 9680 29096 9732 29102
rect 9680 29038 9732 29044
rect 9692 27946 9720 29038
rect 9784 28218 9812 30874
rect 9876 28218 9904 31062
rect 9968 29306 9996 34342
rect 10060 33454 10088 34342
rect 10048 33448 10100 33454
rect 10048 33390 10100 33396
rect 10060 30326 10088 33390
rect 10140 31884 10192 31890
rect 10140 31826 10192 31832
rect 10152 30802 10180 31826
rect 10244 31686 10272 34478
rect 10336 34202 10364 34972
rect 10416 34954 10468 34960
rect 10324 34196 10376 34202
rect 10324 34138 10376 34144
rect 10324 33924 10376 33930
rect 10428 33912 10456 34954
rect 10520 34542 10548 35226
rect 10508 34536 10560 34542
rect 10508 34478 10560 34484
rect 10376 33884 10456 33912
rect 10324 33866 10376 33872
rect 10336 33590 10364 33866
rect 10324 33584 10376 33590
rect 10324 33526 10376 33532
rect 10336 31736 10364 33526
rect 10416 33312 10468 33318
rect 10416 33254 10468 33260
rect 10428 32570 10456 33254
rect 10612 32910 10640 36314
rect 10968 35216 11020 35222
rect 10968 35158 11020 35164
rect 10980 34746 11008 35158
rect 10968 34740 11020 34746
rect 10968 34682 11020 34688
rect 11072 33998 11100 37159
rect 11060 33992 11112 33998
rect 11060 33934 11112 33940
rect 10784 33856 10836 33862
rect 10784 33798 10836 33804
rect 10796 33590 10824 33798
rect 10784 33584 10836 33590
rect 10784 33526 10836 33532
rect 10690 33144 10746 33153
rect 10690 33079 10746 33088
rect 10600 32904 10652 32910
rect 10600 32846 10652 32852
rect 10612 32722 10640 32846
rect 10704 32842 10732 33079
rect 10692 32836 10744 32842
rect 10692 32778 10744 32784
rect 10612 32694 10732 32722
rect 10416 32564 10468 32570
rect 10416 32506 10468 32512
rect 10600 32020 10652 32026
rect 10600 31962 10652 31968
rect 10416 31748 10468 31754
rect 10336 31708 10416 31736
rect 10416 31690 10468 31696
rect 10232 31680 10284 31686
rect 10232 31622 10284 31628
rect 10140 30796 10192 30802
rect 10140 30738 10192 30744
rect 10048 30320 10100 30326
rect 10048 30262 10100 30268
rect 10152 29730 10180 30738
rect 10060 29714 10180 29730
rect 10048 29708 10180 29714
rect 10100 29702 10180 29708
rect 10048 29650 10100 29656
rect 10048 29572 10100 29578
rect 10048 29514 10100 29520
rect 9956 29300 10008 29306
rect 9956 29242 10008 29248
rect 10060 29238 10088 29514
rect 10048 29232 10100 29238
rect 10048 29174 10100 29180
rect 10244 28626 10272 31622
rect 10428 31414 10456 31690
rect 10416 31408 10468 31414
rect 10416 31350 10468 31356
rect 10428 30394 10456 31350
rect 10416 30388 10468 30394
rect 10416 30330 10468 30336
rect 10428 29578 10456 30330
rect 10416 29572 10468 29578
rect 10416 29514 10468 29520
rect 10612 29510 10640 31962
rect 10704 31414 10732 32694
rect 10692 31408 10744 31414
rect 10692 31350 10744 31356
rect 10600 29504 10652 29510
rect 10600 29446 10652 29452
rect 10612 29170 10640 29446
rect 10600 29164 10652 29170
rect 10600 29106 10652 29112
rect 10692 29096 10744 29102
rect 10692 29038 10744 29044
rect 10704 28762 10732 29038
rect 10692 28756 10744 28762
rect 10692 28698 10744 28704
rect 10232 28620 10284 28626
rect 10232 28562 10284 28568
rect 10232 28484 10284 28490
rect 10232 28426 10284 28432
rect 9772 28212 9824 28218
rect 9772 28154 9824 28160
rect 9864 28212 9916 28218
rect 9864 28154 9916 28160
rect 9680 27940 9732 27946
rect 9680 27882 9732 27888
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 10244 7206 10272 28426
rect 10796 26234 10824 33526
rect 11060 33516 11112 33522
rect 11060 33458 11112 33464
rect 10876 32972 10928 32978
rect 10876 32914 10928 32920
rect 10888 32026 10916 32914
rect 10968 32768 11020 32774
rect 10968 32710 11020 32716
rect 10876 32020 10928 32026
rect 10876 31962 10928 31968
rect 10874 28792 10930 28801
rect 10874 28727 10930 28736
rect 10704 26206 10824 26234
rect 10324 25152 10376 25158
rect 10324 25094 10376 25100
rect 10336 24954 10364 25094
rect 10324 24948 10376 24954
rect 10324 24890 10376 24896
rect 10704 9926 10732 26206
rect 10888 25362 10916 28727
rect 10876 25356 10928 25362
rect 10876 25298 10928 25304
rect 10784 24608 10836 24614
rect 10784 24550 10836 24556
rect 10796 24206 10824 24550
rect 10784 24200 10836 24206
rect 10784 24142 10836 24148
rect 10876 24064 10928 24070
rect 10876 24006 10928 24012
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10888 8362 10916 24006
rect 10980 11558 11008 32710
rect 11072 30666 11100 33458
rect 11060 30660 11112 30666
rect 11060 30602 11112 30608
rect 11072 30394 11100 30602
rect 11060 30388 11112 30394
rect 11060 30330 11112 30336
rect 11164 29850 11192 38762
rect 11256 38758 11284 39442
rect 11244 38752 11296 38758
rect 11244 38694 11296 38700
rect 11348 36718 11376 40938
rect 11336 36712 11388 36718
rect 11336 36654 11388 36660
rect 11336 36576 11388 36582
rect 11336 36518 11388 36524
rect 11244 36100 11296 36106
rect 11244 36042 11296 36048
rect 11256 35562 11284 36042
rect 11244 35556 11296 35562
rect 11244 35498 11296 35504
rect 11348 32298 11376 36518
rect 11440 33998 11468 43132
rect 11520 43114 11572 43120
rect 11624 42090 11652 47670
rect 11900 45082 11928 50254
rect 12176 49910 12204 53042
rect 12360 51066 12388 53518
rect 12452 53038 12480 55186
rect 12716 54664 12768 54670
rect 12716 54606 12768 54612
rect 12532 54188 12584 54194
rect 12532 54130 12584 54136
rect 12624 54188 12676 54194
rect 12624 54130 12676 54136
rect 12440 53032 12492 53038
rect 12440 52974 12492 52980
rect 12544 51066 12572 54130
rect 12348 51060 12400 51066
rect 12348 51002 12400 51008
rect 12532 51060 12584 51066
rect 12532 51002 12584 51008
rect 12348 50924 12400 50930
rect 12348 50866 12400 50872
rect 12164 49904 12216 49910
rect 12164 49846 12216 49852
rect 11980 49836 12032 49842
rect 11980 49778 12032 49784
rect 11888 45076 11940 45082
rect 11888 45018 11940 45024
rect 11992 44538 12020 49778
rect 12360 44810 12388 50866
rect 12636 49366 12664 54130
rect 12728 49910 12756 54606
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 13372 53650 13400 55186
rect 13832 54262 13860 56200
rect 13820 54256 13872 54262
rect 13820 54198 13872 54204
rect 13360 53644 13412 53650
rect 13360 53586 13412 53592
rect 13820 53576 13872 53582
rect 13820 53518 13872 53524
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 13360 51468 13412 51474
rect 13360 51410 13412 51416
rect 12808 50924 12860 50930
rect 12808 50866 12860 50872
rect 12716 49904 12768 49910
rect 12716 49846 12768 49852
rect 12624 49360 12676 49366
rect 12624 49302 12676 49308
rect 12716 49156 12768 49162
rect 12716 49098 12768 49104
rect 12728 48346 12756 49098
rect 12716 48340 12768 48346
rect 12716 48282 12768 48288
rect 12532 48136 12584 48142
rect 12532 48078 12584 48084
rect 12544 47802 12572 48078
rect 12624 48000 12676 48006
rect 12624 47942 12676 47948
rect 12532 47796 12584 47802
rect 12532 47738 12584 47744
rect 12532 47592 12584 47598
rect 12532 47534 12584 47540
rect 12544 47054 12572 47534
rect 12440 47048 12492 47054
rect 12440 46990 12492 46996
rect 12532 47048 12584 47054
rect 12532 46990 12584 46996
rect 12452 45082 12480 46990
rect 12532 46572 12584 46578
rect 12532 46514 12584 46520
rect 12440 45076 12492 45082
rect 12440 45018 12492 45024
rect 12544 44962 12572 46514
rect 12636 45558 12664 47942
rect 12716 47184 12768 47190
rect 12716 47126 12768 47132
rect 12624 45552 12676 45558
rect 12624 45494 12676 45500
rect 12728 45014 12756 47126
rect 12820 45286 12848 50866
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 13372 49230 13400 51410
rect 13636 50720 13688 50726
rect 13636 50662 13688 50668
rect 13648 50454 13676 50662
rect 13636 50448 13688 50454
rect 13636 50390 13688 50396
rect 13636 50244 13688 50250
rect 13636 50186 13688 50192
rect 13648 49994 13676 50186
rect 13648 49978 13768 49994
rect 13648 49972 13780 49978
rect 13648 49966 13728 49972
rect 13360 49224 13412 49230
rect 13360 49166 13412 49172
rect 13544 49088 13596 49094
rect 13544 49030 13596 49036
rect 13360 48544 13412 48550
rect 13360 48486 13412 48492
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 13268 48340 13320 48346
rect 13268 48282 13320 48288
rect 13280 47512 13308 48282
rect 13372 48142 13400 48486
rect 13360 48136 13412 48142
rect 13360 48078 13412 48084
rect 13280 47484 13400 47512
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 13372 47002 13400 47484
rect 13556 47258 13584 49030
rect 13648 48210 13676 49966
rect 13728 49914 13780 49920
rect 13832 49910 13860 53518
rect 14372 53168 14424 53174
rect 14372 53110 14424 53116
rect 14188 51400 14240 51406
rect 14188 51342 14240 51348
rect 14096 50856 14148 50862
rect 14096 50798 14148 50804
rect 14108 50318 14136 50798
rect 14096 50312 14148 50318
rect 14096 50254 14148 50260
rect 13820 49904 13872 49910
rect 13820 49846 13872 49852
rect 14108 49774 14136 50254
rect 14096 49768 14148 49774
rect 14096 49710 14148 49716
rect 13820 49360 13872 49366
rect 13820 49302 13872 49308
rect 13636 48204 13688 48210
rect 13636 48146 13688 48152
rect 13832 48142 13860 49302
rect 14108 48890 14136 49710
rect 14096 48884 14148 48890
rect 14096 48826 14148 48832
rect 14108 48210 14136 48826
rect 14096 48204 14148 48210
rect 14096 48146 14148 48152
rect 13820 48136 13872 48142
rect 13820 48078 13872 48084
rect 13728 47728 13780 47734
rect 13728 47670 13780 47676
rect 13636 47592 13688 47598
rect 13636 47534 13688 47540
rect 13544 47252 13596 47258
rect 13544 47194 13596 47200
rect 13648 47122 13676 47534
rect 13636 47116 13688 47122
rect 13636 47058 13688 47064
rect 12900 46980 12952 46986
rect 13372 46974 13492 47002
rect 12900 46922 12952 46928
rect 12912 46578 12940 46922
rect 13360 46912 13412 46918
rect 13360 46854 13412 46860
rect 12900 46572 12952 46578
rect 12900 46514 12952 46520
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 13372 46170 13400 46854
rect 13360 46164 13412 46170
rect 13360 46106 13412 46112
rect 12808 45280 12860 45286
rect 12808 45222 12860 45228
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 12716 45008 12768 45014
rect 12544 44934 12664 44962
rect 12716 44950 12768 44956
rect 13084 45008 13136 45014
rect 13084 44950 13136 44956
rect 12440 44872 12492 44878
rect 12440 44814 12492 44820
rect 12532 44872 12584 44878
rect 12532 44814 12584 44820
rect 12348 44804 12400 44810
rect 12348 44746 12400 44752
rect 11980 44532 12032 44538
rect 11980 44474 12032 44480
rect 12348 44192 12400 44198
rect 12348 44134 12400 44140
rect 11796 43852 11848 43858
rect 11796 43794 11848 43800
rect 11808 42906 11836 43794
rect 12360 43450 12388 44134
rect 12348 43444 12400 43450
rect 12348 43386 12400 43392
rect 12176 43302 12388 43330
rect 12176 43246 12204 43302
rect 12164 43240 12216 43246
rect 12164 43182 12216 43188
rect 12256 43240 12308 43246
rect 12256 43182 12308 43188
rect 11796 42900 11848 42906
rect 11796 42842 11848 42848
rect 12268 42344 12296 43182
rect 12084 42316 12296 42344
rect 11612 42084 11664 42090
rect 11612 42026 11664 42032
rect 11980 42016 12032 42022
rect 11980 41958 12032 41964
rect 11992 41750 12020 41958
rect 11980 41744 12032 41750
rect 11980 41686 12032 41692
rect 11888 41676 11940 41682
rect 11888 41618 11940 41624
rect 11900 41414 11928 41618
rect 11624 41386 11928 41414
rect 11520 41268 11572 41274
rect 11520 41210 11572 41216
rect 11532 39982 11560 41210
rect 11520 39976 11572 39982
rect 11520 39918 11572 39924
rect 11624 38010 11652 41386
rect 11704 41132 11756 41138
rect 11704 41074 11756 41080
rect 11716 40050 11744 41074
rect 11888 40928 11940 40934
rect 11888 40870 11940 40876
rect 11704 40044 11756 40050
rect 11704 39986 11756 39992
rect 11704 39840 11756 39846
rect 11704 39782 11756 39788
rect 11716 39030 11744 39782
rect 11900 39438 11928 40870
rect 11992 40730 12020 41686
rect 12084 41274 12112 42316
rect 12164 42220 12216 42226
rect 12164 42162 12216 42168
rect 12072 41268 12124 41274
rect 12072 41210 12124 41216
rect 12070 41168 12126 41177
rect 12070 41103 12126 41112
rect 11980 40724 12032 40730
rect 11980 40666 12032 40672
rect 12084 40118 12112 41103
rect 12176 40225 12204 42162
rect 12256 41472 12308 41478
rect 12256 41414 12308 41420
rect 12268 41070 12296 41414
rect 12256 41064 12308 41070
rect 12256 41006 12308 41012
rect 12268 40633 12296 41006
rect 12254 40624 12310 40633
rect 12254 40559 12310 40568
rect 12360 40338 12388 43302
rect 12452 42362 12480 44814
rect 12544 43790 12572 44814
rect 12532 43784 12584 43790
rect 12532 43726 12584 43732
rect 12532 43376 12584 43382
rect 12532 43318 12584 43324
rect 12440 42356 12492 42362
rect 12440 42298 12492 42304
rect 12544 40730 12572 43318
rect 12636 41818 12664 44934
rect 13096 44470 13124 44950
rect 13464 44826 13492 46974
rect 13544 46912 13596 46918
rect 13544 46854 13596 46860
rect 13372 44798 13492 44826
rect 13084 44464 13136 44470
rect 13084 44406 13136 44412
rect 12808 44396 12860 44402
rect 12808 44338 12860 44344
rect 12716 42628 12768 42634
rect 12716 42570 12768 42576
rect 12624 41812 12676 41818
rect 12624 41754 12676 41760
rect 12728 41614 12756 42570
rect 12716 41608 12768 41614
rect 12716 41550 12768 41556
rect 12728 41206 12756 41550
rect 12716 41200 12768 41206
rect 12622 41168 12678 41177
rect 12716 41142 12768 41148
rect 12622 41103 12678 41112
rect 12532 40724 12584 40730
rect 12532 40666 12584 40672
rect 12268 40310 12388 40338
rect 12162 40216 12218 40225
rect 12162 40151 12218 40160
rect 12072 40112 12124 40118
rect 12268 40066 12296 40310
rect 12346 40216 12402 40225
rect 12346 40151 12348 40160
rect 12400 40151 12402 40160
rect 12348 40122 12400 40128
rect 12072 40054 12124 40060
rect 12176 40038 12296 40066
rect 11980 39976 12032 39982
rect 11980 39918 12032 39924
rect 11888 39432 11940 39438
rect 11888 39374 11940 39380
rect 11704 39024 11756 39030
rect 11704 38966 11756 38972
rect 11888 38888 11940 38894
rect 11886 38856 11888 38865
rect 11940 38856 11942 38865
rect 11886 38791 11942 38800
rect 11992 38554 12020 39918
rect 12072 39364 12124 39370
rect 12072 39306 12124 39312
rect 12084 39001 12112 39306
rect 12070 38992 12126 39001
rect 12070 38927 12126 38936
rect 11980 38548 12032 38554
rect 11980 38490 12032 38496
rect 11980 38344 12032 38350
rect 11980 38286 12032 38292
rect 11612 38004 11664 38010
rect 11612 37946 11664 37952
rect 11992 37262 12020 38286
rect 12176 38010 12204 40038
rect 12254 39944 12310 39953
rect 12254 39879 12310 39888
rect 12268 39642 12296 39879
rect 12256 39636 12308 39642
rect 12256 39578 12308 39584
rect 12256 39432 12308 39438
rect 12256 39374 12308 39380
rect 12164 38004 12216 38010
rect 12164 37946 12216 37952
rect 11980 37256 12032 37262
rect 11980 37198 12032 37204
rect 11992 37074 12020 37198
rect 11992 37046 12112 37074
rect 12084 36854 12112 37046
rect 12072 36848 12124 36854
rect 12268 36825 12296 39374
rect 12072 36790 12124 36796
rect 12254 36816 12310 36825
rect 11796 36780 11848 36786
rect 11796 36722 11848 36728
rect 11808 36378 11836 36722
rect 11796 36372 11848 36378
rect 11796 36314 11848 36320
rect 11520 35760 11572 35766
rect 11520 35702 11572 35708
rect 11428 33992 11480 33998
rect 11428 33934 11480 33940
rect 11428 33856 11480 33862
rect 11428 33798 11480 33804
rect 11336 32292 11388 32298
rect 11336 32234 11388 32240
rect 11244 32224 11296 32230
rect 11244 32166 11296 32172
rect 11152 29844 11204 29850
rect 11152 29786 11204 29792
rect 11256 29073 11284 32166
rect 11336 31272 11388 31278
rect 11336 31214 11388 31220
rect 11348 29850 11376 31214
rect 11336 29844 11388 29850
rect 11336 29786 11388 29792
rect 11242 29064 11298 29073
rect 11242 28999 11298 29008
rect 11348 26994 11376 29786
rect 11440 28558 11468 33798
rect 11428 28552 11480 28558
rect 11428 28494 11480 28500
rect 11532 27606 11560 35702
rect 12084 35154 12112 36790
rect 12360 36786 12388 40122
rect 12440 39976 12492 39982
rect 12438 39944 12440 39953
rect 12492 39944 12494 39953
rect 12438 39879 12494 39888
rect 12636 39386 12664 41103
rect 12716 40520 12768 40526
rect 12716 40462 12768 40468
rect 12452 39358 12664 39386
rect 12254 36751 12310 36760
rect 12348 36780 12400 36786
rect 12348 36722 12400 36728
rect 12348 35624 12400 35630
rect 12348 35566 12400 35572
rect 12072 35148 12124 35154
rect 12072 35090 12124 35096
rect 12084 34610 12112 35090
rect 12360 34678 12388 35566
rect 12348 34672 12400 34678
rect 12348 34614 12400 34620
rect 11888 34604 11940 34610
rect 11888 34546 11940 34552
rect 12072 34604 12124 34610
rect 12072 34546 12124 34552
rect 11704 32904 11756 32910
rect 11704 32846 11756 32852
rect 11716 32570 11744 32846
rect 11704 32564 11756 32570
rect 11704 32506 11756 32512
rect 11900 32434 11928 34546
rect 12072 34400 12124 34406
rect 12072 34342 12124 34348
rect 12164 34400 12216 34406
rect 12164 34342 12216 34348
rect 12084 34202 12112 34342
rect 12072 34196 12124 34202
rect 12072 34138 12124 34144
rect 12176 33930 12204 34342
rect 12164 33924 12216 33930
rect 12164 33866 12216 33872
rect 12256 33924 12308 33930
rect 12256 33866 12308 33872
rect 12072 33856 12124 33862
rect 12072 33798 12124 33804
rect 11980 32836 12032 32842
rect 11980 32778 12032 32784
rect 11888 32428 11940 32434
rect 11888 32370 11940 32376
rect 11992 31958 12020 32778
rect 11980 31952 12032 31958
rect 11980 31894 12032 31900
rect 11704 31816 11756 31822
rect 11704 31758 11756 31764
rect 11716 31278 11744 31758
rect 12084 31754 12112 33798
rect 11992 31726 12112 31754
rect 11704 31272 11756 31278
rect 11704 31214 11756 31220
rect 11716 30802 11744 31214
rect 11704 30796 11756 30802
rect 11704 30738 11756 30744
rect 11612 30660 11664 30666
rect 11612 30602 11664 30608
rect 11624 30326 11652 30602
rect 11888 30592 11940 30598
rect 11888 30534 11940 30540
rect 11704 30388 11756 30394
rect 11704 30330 11756 30336
rect 11612 30320 11664 30326
rect 11612 30262 11664 30268
rect 11612 28688 11664 28694
rect 11612 28630 11664 28636
rect 11520 27600 11572 27606
rect 11520 27542 11572 27548
rect 11336 26988 11388 26994
rect 11336 26930 11388 26936
rect 11624 26234 11652 28630
rect 11716 28626 11744 30330
rect 11796 30252 11848 30258
rect 11796 30194 11848 30200
rect 11808 29714 11836 30194
rect 11796 29708 11848 29714
rect 11796 29650 11848 29656
rect 11900 29646 11928 30534
rect 11888 29640 11940 29646
rect 11888 29582 11940 29588
rect 11704 28620 11756 28626
rect 11704 28562 11756 28568
rect 11992 28558 12020 31726
rect 12072 29028 12124 29034
rect 12072 28970 12124 28976
rect 11980 28552 12032 28558
rect 11980 28494 12032 28500
rect 12084 27130 12112 28970
rect 12072 27124 12124 27130
rect 12072 27066 12124 27072
rect 12176 26234 12204 33866
rect 12268 33522 12296 33866
rect 12256 33516 12308 33522
rect 12256 33458 12308 33464
rect 12360 33114 12388 34614
rect 12452 34066 12480 39358
rect 12624 39296 12676 39302
rect 12530 39264 12586 39273
rect 12624 39238 12676 39244
rect 12530 39199 12586 39208
rect 12544 39098 12572 39199
rect 12532 39092 12584 39098
rect 12532 39034 12584 39040
rect 12532 38956 12584 38962
rect 12532 38898 12584 38904
rect 12544 38729 12572 38898
rect 12530 38720 12586 38729
rect 12530 38655 12586 38664
rect 12532 38208 12584 38214
rect 12636 38196 12664 39238
rect 12728 39030 12756 40462
rect 12716 39024 12768 39030
rect 12716 38966 12768 38972
rect 12716 38276 12768 38282
rect 12716 38218 12768 38224
rect 12584 38168 12664 38196
rect 12532 38150 12584 38156
rect 12728 38010 12756 38218
rect 12716 38004 12768 38010
rect 12716 37946 12768 37952
rect 12624 37868 12676 37874
rect 12624 37810 12676 37816
rect 12636 36922 12664 37810
rect 12728 37194 12756 37946
rect 12716 37188 12768 37194
rect 12716 37130 12768 37136
rect 12624 36916 12676 36922
rect 12624 36858 12676 36864
rect 12728 35766 12756 37130
rect 12820 36378 12848 44338
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 13372 43874 13400 44798
rect 13452 44736 13504 44742
rect 13452 44678 13504 44684
rect 13280 43846 13400 43874
rect 13280 43654 13308 43846
rect 13360 43716 13412 43722
rect 13360 43658 13412 43664
rect 13268 43648 13320 43654
rect 13268 43590 13320 43596
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 12990 40624 13046 40633
rect 12990 40559 12992 40568
rect 13044 40559 13046 40568
rect 12992 40530 13044 40536
rect 13268 40452 13320 40458
rect 13268 40394 13320 40400
rect 13280 39982 13308 40394
rect 13268 39976 13320 39982
rect 13268 39918 13320 39924
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 13372 39642 13400 43658
rect 13360 39636 13412 39642
rect 13360 39578 13412 39584
rect 12898 39536 12954 39545
rect 12898 39471 12954 39480
rect 13082 39536 13138 39545
rect 13082 39471 13138 39480
rect 12912 39438 12940 39471
rect 12900 39432 12952 39438
rect 12900 39374 12952 39380
rect 12990 39128 13046 39137
rect 12990 39063 13046 39072
rect 13004 38894 13032 39063
rect 13096 38962 13124 39471
rect 13464 39114 13492 44678
rect 13556 43450 13584 46854
rect 13636 45076 13688 45082
rect 13636 45018 13688 45024
rect 13544 43444 13596 43450
rect 13544 43386 13596 43392
rect 13648 42650 13676 45018
rect 13740 42786 13768 47670
rect 14004 47592 14056 47598
rect 14004 47534 14056 47540
rect 13912 47184 13964 47190
rect 13912 47126 13964 47132
rect 13924 46986 13952 47126
rect 14016 47054 14044 47534
rect 14004 47048 14056 47054
rect 14004 46990 14056 46996
rect 13912 46980 13964 46986
rect 13912 46922 13964 46928
rect 14004 46504 14056 46510
rect 14004 46446 14056 46452
rect 14016 46170 14044 46446
rect 14004 46164 14056 46170
rect 14004 46106 14056 46112
rect 14200 45354 14228 51342
rect 14384 50998 14412 53110
rect 14476 52562 14504 56200
rect 15120 52970 15148 56200
rect 15764 54262 15792 56200
rect 15752 54256 15804 54262
rect 15752 54198 15804 54204
rect 16408 53650 16436 56200
rect 16488 54052 16540 54058
rect 16488 53994 16540 54000
rect 16396 53644 16448 53650
rect 16396 53586 16448 53592
rect 15568 53100 15620 53106
rect 15568 53042 15620 53048
rect 15108 52964 15160 52970
rect 15108 52906 15160 52912
rect 14648 52692 14700 52698
rect 14648 52634 14700 52640
rect 14464 52556 14516 52562
rect 14464 52498 14516 52504
rect 14556 52488 14608 52494
rect 14556 52430 14608 52436
rect 14464 52012 14516 52018
rect 14464 51954 14516 51960
rect 14372 50992 14424 50998
rect 14372 50934 14424 50940
rect 14280 47456 14332 47462
rect 14280 47398 14332 47404
rect 14292 47122 14320 47398
rect 14280 47116 14332 47122
rect 14280 47058 14332 47064
rect 14476 46730 14504 51954
rect 14568 51610 14596 52430
rect 14660 51610 14688 52634
rect 15580 52154 15608 53042
rect 15568 52148 15620 52154
rect 15568 52090 15620 52096
rect 16304 51808 16356 51814
rect 16304 51750 16356 51756
rect 14556 51604 14608 51610
rect 14556 51546 14608 51552
rect 14648 51604 14700 51610
rect 14648 51546 14700 51552
rect 14660 49230 14688 51546
rect 16120 51468 16172 51474
rect 16120 51410 16172 51416
rect 15844 51400 15896 51406
rect 15844 51342 15896 51348
rect 15660 51332 15712 51338
rect 15660 51274 15712 51280
rect 15292 50992 15344 50998
rect 15212 50940 15292 50946
rect 15212 50934 15344 50940
rect 15212 50918 15332 50934
rect 15212 50250 15240 50918
rect 15200 50244 15252 50250
rect 15200 50186 15252 50192
rect 14832 49904 14884 49910
rect 14832 49846 14884 49852
rect 14844 49688 14872 49846
rect 15212 49688 15240 50186
rect 15568 50176 15620 50182
rect 15568 50118 15620 50124
rect 14752 49660 15240 49688
rect 14648 49224 14700 49230
rect 14648 49166 14700 49172
rect 14752 48822 14780 49660
rect 14924 49292 14976 49298
rect 14924 49234 14976 49240
rect 15016 49292 15068 49298
rect 15016 49234 15068 49240
rect 14936 49094 14964 49234
rect 14924 49088 14976 49094
rect 14924 49030 14976 49036
rect 14740 48816 14792 48822
rect 14740 48758 14792 48764
rect 14648 48544 14700 48550
rect 14648 48486 14700 48492
rect 14556 47116 14608 47122
rect 14556 47058 14608 47064
rect 14384 46702 14504 46730
rect 14188 45348 14240 45354
rect 14188 45290 14240 45296
rect 14384 45082 14412 46702
rect 14464 46572 14516 46578
rect 14464 46514 14516 46520
rect 14476 45354 14504 46514
rect 14568 46510 14596 47058
rect 14660 46986 14688 48486
rect 14752 47666 14780 48758
rect 15028 48686 15056 49234
rect 15016 48680 15068 48686
rect 15016 48622 15068 48628
rect 14924 48068 14976 48074
rect 14924 48010 14976 48016
rect 14740 47660 14792 47666
rect 14740 47602 14792 47608
rect 14740 47456 14792 47462
rect 14740 47398 14792 47404
rect 14648 46980 14700 46986
rect 14648 46922 14700 46928
rect 14556 46504 14608 46510
rect 14556 46446 14608 46452
rect 14568 45966 14596 46446
rect 14556 45960 14608 45966
rect 14556 45902 14608 45908
rect 14648 45484 14700 45490
rect 14648 45426 14700 45432
rect 14464 45348 14516 45354
rect 14464 45290 14516 45296
rect 14372 45076 14424 45082
rect 14372 45018 14424 45024
rect 14464 44872 14516 44878
rect 14464 44814 14516 44820
rect 13912 44532 13964 44538
rect 13912 44474 13964 44480
rect 13820 44260 13872 44266
rect 13820 44202 13872 44208
rect 13832 43858 13860 44202
rect 13820 43852 13872 43858
rect 13820 43794 13872 43800
rect 13924 43790 13952 44474
rect 14004 43852 14056 43858
rect 14004 43794 14056 43800
rect 13912 43784 13964 43790
rect 13912 43726 13964 43732
rect 14016 43314 14044 43794
rect 14004 43308 14056 43314
rect 14004 43250 14056 43256
rect 14188 42900 14240 42906
rect 14188 42842 14240 42848
rect 13740 42758 13952 42786
rect 13648 42622 13768 42650
rect 13636 42560 13688 42566
rect 13636 42502 13688 42508
rect 13544 42152 13596 42158
rect 13544 42094 13596 42100
rect 13556 39273 13584 42094
rect 13648 41070 13676 42502
rect 13740 42022 13768 42622
rect 13820 42628 13872 42634
rect 13820 42570 13872 42576
rect 13728 42016 13780 42022
rect 13728 41958 13780 41964
rect 13636 41064 13688 41070
rect 13636 41006 13688 41012
rect 13648 40934 13676 41006
rect 13636 40928 13688 40934
rect 13636 40870 13688 40876
rect 13832 40050 13860 42570
rect 13924 42566 13952 42758
rect 13912 42560 13964 42566
rect 13912 42502 13964 42508
rect 14096 41676 14148 41682
rect 14096 41618 14148 41624
rect 14108 41070 14136 41618
rect 14200 41414 14228 42842
rect 14280 42016 14332 42022
rect 14280 41958 14332 41964
rect 14292 41750 14320 41958
rect 14370 41848 14426 41857
rect 14370 41783 14426 41792
rect 14280 41744 14332 41750
rect 14280 41686 14332 41692
rect 14200 41386 14320 41414
rect 14096 41064 14148 41070
rect 14096 41006 14148 41012
rect 14188 41064 14240 41070
rect 14188 41006 14240 41012
rect 14108 40458 14136 41006
rect 14096 40452 14148 40458
rect 14096 40394 14148 40400
rect 14200 40390 14228 41006
rect 14188 40384 14240 40390
rect 14108 40332 14188 40338
rect 14108 40326 14240 40332
rect 14108 40310 14228 40326
rect 13820 40044 13872 40050
rect 13820 39986 13872 39992
rect 13912 40044 13964 40050
rect 13912 39986 13964 39992
rect 13636 39976 13688 39982
rect 13636 39918 13688 39924
rect 13542 39264 13598 39273
rect 13542 39199 13598 39208
rect 13648 39137 13676 39918
rect 13188 39098 13492 39114
rect 13176 39092 13492 39098
rect 13228 39086 13492 39092
rect 13634 39128 13690 39137
rect 13634 39063 13690 39072
rect 13176 39034 13228 39040
rect 13084 38956 13136 38962
rect 13084 38898 13136 38904
rect 12992 38888 13044 38894
rect 12992 38830 13044 38836
rect 13452 38888 13504 38894
rect 13452 38830 13504 38836
rect 13636 38888 13688 38894
rect 13636 38830 13688 38836
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 13084 38208 13136 38214
rect 13084 38150 13136 38156
rect 13096 37806 13124 38150
rect 12992 37800 13044 37806
rect 12990 37768 12992 37777
rect 13084 37800 13136 37806
rect 13044 37768 13046 37777
rect 13084 37742 13136 37748
rect 12990 37703 13046 37712
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 12808 36372 12860 36378
rect 12808 36314 12860 36320
rect 12808 36032 12860 36038
rect 12808 35974 12860 35980
rect 13360 36032 13412 36038
rect 13360 35974 13412 35980
rect 12716 35760 12768 35766
rect 12636 35720 12716 35748
rect 12636 34678 12664 35720
rect 12716 35702 12768 35708
rect 12820 35290 12848 35974
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 12808 35284 12860 35290
rect 12808 35226 12860 35232
rect 13372 35170 13400 35974
rect 13464 35290 13492 38830
rect 13648 37346 13676 38830
rect 13818 38040 13874 38049
rect 13818 37975 13874 37984
rect 13832 37942 13860 37975
rect 13820 37936 13872 37942
rect 13820 37878 13872 37884
rect 13728 37800 13780 37806
rect 13728 37742 13780 37748
rect 13740 37466 13768 37742
rect 13728 37460 13780 37466
rect 13728 37402 13780 37408
rect 13556 37330 13676 37346
rect 13544 37324 13676 37330
rect 13596 37318 13676 37324
rect 13544 37266 13596 37272
rect 13556 35834 13584 37266
rect 13820 36780 13872 36786
rect 13820 36722 13872 36728
rect 13728 36236 13780 36242
rect 13728 36178 13780 36184
rect 13544 35828 13596 35834
rect 13544 35770 13596 35776
rect 13544 35624 13596 35630
rect 13544 35566 13596 35572
rect 13452 35284 13504 35290
rect 13452 35226 13504 35232
rect 13280 35142 13400 35170
rect 13556 35154 13584 35566
rect 13544 35148 13596 35154
rect 12808 35012 12860 35018
rect 12808 34954 12860 34960
rect 12624 34672 12676 34678
rect 12624 34614 12676 34620
rect 12440 34060 12492 34066
rect 12440 34002 12492 34008
rect 12636 33969 12664 34614
rect 12622 33960 12678 33969
rect 12622 33895 12678 33904
rect 12348 33108 12400 33114
rect 12348 33050 12400 33056
rect 12636 32824 12664 33895
rect 12716 32836 12768 32842
rect 12636 32796 12716 32824
rect 12716 32778 12768 32784
rect 12728 32502 12756 32778
rect 12716 32496 12768 32502
rect 12452 32422 12664 32450
rect 12716 32438 12768 32444
rect 12348 31884 12400 31890
rect 12348 31826 12400 31832
rect 12360 27538 12388 31826
rect 12452 28626 12480 32422
rect 12636 32366 12664 32422
rect 12624 32360 12676 32366
rect 12624 32302 12676 32308
rect 12624 32224 12676 32230
rect 12624 32166 12676 32172
rect 12532 31748 12584 31754
rect 12532 31690 12584 31696
rect 12544 31414 12572 31690
rect 12532 31408 12584 31414
rect 12532 31350 12584 31356
rect 12544 30326 12572 31350
rect 12636 30598 12664 32166
rect 12728 31754 12756 32438
rect 12716 31748 12768 31754
rect 12716 31690 12768 31696
rect 12728 31482 12756 31690
rect 12716 31476 12768 31482
rect 12716 31418 12768 31424
rect 12624 30592 12676 30598
rect 12624 30534 12676 30540
rect 12532 30320 12584 30326
rect 12532 30262 12584 30268
rect 12636 30190 12664 30534
rect 12624 30184 12676 30190
rect 12624 30126 12676 30132
rect 12636 29238 12664 30126
rect 12624 29232 12676 29238
rect 12624 29174 12676 29180
rect 12820 29102 12848 34954
rect 13280 34388 13308 35142
rect 13544 35090 13596 35096
rect 13360 35080 13412 35086
rect 13358 35048 13360 35057
rect 13412 35048 13414 35057
rect 13358 34983 13414 34992
rect 13556 34542 13584 35090
rect 13636 34604 13688 34610
rect 13636 34546 13688 34552
rect 13544 34536 13596 34542
rect 13544 34478 13596 34484
rect 13280 34360 13492 34388
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 12992 34060 13044 34066
rect 12992 34002 13044 34008
rect 13004 33930 13032 34002
rect 12900 33924 12952 33930
rect 12900 33866 12952 33872
rect 12992 33924 13044 33930
rect 12992 33866 13044 33872
rect 12912 33658 12940 33866
rect 13360 33856 13412 33862
rect 13360 33798 13412 33804
rect 12900 33652 12952 33658
rect 12900 33594 12952 33600
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 13372 32366 13400 33798
rect 13360 32360 13412 32366
rect 13360 32302 13412 32308
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 13268 29708 13320 29714
rect 13268 29650 13320 29656
rect 12532 29096 12584 29102
rect 12808 29096 12860 29102
rect 12532 29038 12584 29044
rect 12622 29064 12678 29073
rect 12440 28620 12492 28626
rect 12440 28562 12492 28568
rect 12348 27532 12400 27538
rect 12348 27474 12400 27480
rect 11532 26206 11652 26234
rect 11992 26206 12204 26234
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 9220 5296 9272 5302
rect 9220 5238 9272 5244
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 8852 2508 8904 2514
rect 8852 2450 8904 2456
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 8864 800 8892 2450
rect 10704 2310 10732 7754
rect 11532 5574 11560 26206
rect 11992 12102 12020 26206
rect 12544 25498 12572 29038
rect 12808 29038 12860 29044
rect 13280 29017 13308 29650
rect 13464 29322 13492 34360
rect 13544 33992 13596 33998
rect 13544 33934 13596 33940
rect 13556 31414 13584 33934
rect 13648 33590 13676 34546
rect 13636 33584 13688 33590
rect 13636 33526 13688 33532
rect 13740 32586 13768 36178
rect 13832 32774 13860 36722
rect 13924 36174 13952 39986
rect 14004 39500 14056 39506
rect 14004 39442 14056 39448
rect 14016 38962 14044 39442
rect 14004 38956 14056 38962
rect 14004 38898 14056 38904
rect 14004 38752 14056 38758
rect 14004 38694 14056 38700
rect 13912 36168 13964 36174
rect 13912 36110 13964 36116
rect 14016 34678 14044 38694
rect 14108 37806 14136 40310
rect 14188 39296 14240 39302
rect 14188 39238 14240 39244
rect 14200 39098 14228 39238
rect 14188 39092 14240 39098
rect 14188 39034 14240 39040
rect 14186 38856 14242 38865
rect 14292 38826 14320 41386
rect 14186 38791 14242 38800
rect 14280 38820 14332 38826
rect 14096 37800 14148 37806
rect 14096 37742 14148 37748
rect 14096 35692 14148 35698
rect 14096 35634 14148 35640
rect 14004 34672 14056 34678
rect 14004 34614 14056 34620
rect 14004 34468 14056 34474
rect 14004 34410 14056 34416
rect 13912 34196 13964 34202
rect 13912 34138 13964 34144
rect 13924 33930 13952 34138
rect 13912 33924 13964 33930
rect 13912 33866 13964 33872
rect 13820 32768 13872 32774
rect 13820 32710 13872 32716
rect 13740 32558 13860 32586
rect 13832 32366 13860 32558
rect 13820 32360 13872 32366
rect 13740 32308 13820 32314
rect 13740 32302 13872 32308
rect 13740 32286 13860 32302
rect 13740 32026 13768 32286
rect 13820 32224 13872 32230
rect 13820 32166 13872 32172
rect 13728 32020 13780 32026
rect 13728 31962 13780 31968
rect 13832 31906 13860 32166
rect 13740 31878 13860 31906
rect 13544 31408 13596 31414
rect 13544 31350 13596 31356
rect 13544 31272 13596 31278
rect 13544 31214 13596 31220
rect 13556 30190 13584 31214
rect 13544 30184 13596 30190
rect 13544 30126 13596 30132
rect 13556 29458 13584 30126
rect 13740 29714 13768 31878
rect 13820 30184 13872 30190
rect 13820 30126 13872 30132
rect 13728 29708 13780 29714
rect 13728 29650 13780 29656
rect 13728 29572 13780 29578
rect 13728 29514 13780 29520
rect 13556 29430 13676 29458
rect 13464 29294 13584 29322
rect 13360 29096 13412 29102
rect 13360 29038 13412 29044
rect 12622 28999 12678 29008
rect 13266 29008 13322 29017
rect 12636 28150 12664 28999
rect 12808 28960 12860 28966
rect 13266 28943 13322 28952
rect 12808 28902 12860 28908
rect 12716 28416 12768 28422
rect 12716 28358 12768 28364
rect 12624 28144 12676 28150
rect 12624 28086 12676 28092
rect 12532 25492 12584 25498
rect 12532 25434 12584 25440
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 12452 23050 12480 24142
rect 12532 23656 12584 23662
rect 12532 23598 12584 23604
rect 12440 23044 12492 23050
rect 12440 22986 12492 22992
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 12360 4078 12388 22918
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 12544 3534 12572 23598
rect 12728 13190 12756 28358
rect 12820 28218 12848 28902
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 13372 28762 13400 29038
rect 13556 28762 13584 29294
rect 13360 28756 13412 28762
rect 13360 28698 13412 28704
rect 13544 28756 13596 28762
rect 13544 28698 13596 28704
rect 12808 28212 12860 28218
rect 12808 28154 12860 28160
rect 13648 28014 13676 29430
rect 13740 28914 13768 29514
rect 13832 29017 13860 30126
rect 13924 29209 13952 33866
rect 14016 33522 14044 34410
rect 14004 33516 14056 33522
rect 14004 33458 14056 33464
rect 14004 33380 14056 33386
rect 14004 33322 14056 33328
rect 14016 33114 14044 33322
rect 14004 33108 14056 33114
rect 14004 33050 14056 33056
rect 14108 30122 14136 35634
rect 14096 30116 14148 30122
rect 14096 30058 14148 30064
rect 13910 29200 13966 29209
rect 13910 29135 13966 29144
rect 13818 29008 13874 29017
rect 13818 28943 13874 28952
rect 14004 28960 14056 28966
rect 14002 28928 14004 28937
rect 14056 28928 14058 28937
rect 13740 28886 13952 28914
rect 13818 28792 13874 28801
rect 13818 28727 13874 28736
rect 13636 28008 13688 28014
rect 13636 27950 13688 27956
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 13832 24206 13860 28727
rect 13924 24410 13952 28886
rect 14002 28863 14058 28872
rect 14200 27470 14228 38791
rect 14280 38762 14332 38768
rect 14280 38344 14332 38350
rect 14280 38286 14332 38292
rect 14292 37330 14320 38286
rect 14280 37324 14332 37330
rect 14280 37266 14332 37272
rect 14292 36854 14320 37266
rect 14280 36848 14332 36854
rect 14280 36790 14332 36796
rect 14280 36168 14332 36174
rect 14280 36110 14332 36116
rect 14292 35494 14320 36110
rect 14280 35488 14332 35494
rect 14280 35430 14332 35436
rect 14292 34542 14320 35430
rect 14280 34536 14332 34542
rect 14280 34478 14332 34484
rect 14292 33998 14320 34478
rect 14384 34474 14412 41783
rect 14476 39302 14504 44814
rect 14556 42152 14608 42158
rect 14556 42094 14608 42100
rect 14568 41614 14596 42094
rect 14556 41608 14608 41614
rect 14556 41550 14608 41556
rect 14568 41274 14596 41550
rect 14556 41268 14608 41274
rect 14556 41210 14608 41216
rect 14568 40594 14596 41210
rect 14556 40588 14608 40594
rect 14556 40530 14608 40536
rect 14464 39296 14516 39302
rect 14464 39238 14516 39244
rect 14568 38418 14596 40530
rect 14660 39642 14688 45426
rect 14752 44946 14780 47398
rect 14936 46170 14964 48010
rect 15028 47598 15056 48622
rect 15200 48544 15252 48550
rect 15200 48486 15252 48492
rect 15016 47592 15068 47598
rect 15016 47534 15068 47540
rect 14924 46164 14976 46170
rect 14924 46106 14976 46112
rect 15108 45824 15160 45830
rect 15108 45766 15160 45772
rect 15016 45280 15068 45286
rect 15016 45222 15068 45228
rect 14740 44940 14792 44946
rect 14740 44882 14792 44888
rect 15028 43790 15056 45222
rect 15120 44146 15148 45766
rect 15212 45422 15240 48486
rect 15200 45416 15252 45422
rect 15200 45358 15252 45364
rect 15384 44804 15436 44810
rect 15384 44746 15436 44752
rect 15292 44736 15344 44742
rect 15292 44678 15344 44684
rect 15120 44118 15240 44146
rect 15212 43790 15240 44118
rect 15016 43784 15068 43790
rect 15016 43726 15068 43732
rect 15200 43784 15252 43790
rect 15200 43726 15252 43732
rect 14924 43308 14976 43314
rect 14924 43250 14976 43256
rect 14832 42152 14884 42158
rect 14832 42094 14884 42100
rect 14738 41712 14794 41721
rect 14738 41647 14740 41656
rect 14792 41647 14794 41656
rect 14740 41618 14792 41624
rect 14648 39636 14700 39642
rect 14648 39578 14700 39584
rect 14740 39568 14792 39574
rect 14844 39556 14872 42094
rect 14936 41041 14964 43250
rect 15200 42764 15252 42770
rect 15200 42706 15252 42712
rect 15212 42362 15240 42706
rect 15200 42356 15252 42362
rect 15200 42298 15252 42304
rect 15108 42288 15160 42294
rect 15304 42242 15332 44678
rect 15160 42236 15332 42242
rect 15108 42230 15332 42236
rect 15120 42214 15332 42230
rect 15396 41750 15424 44746
rect 15476 43784 15528 43790
rect 15476 43726 15528 43732
rect 15488 43246 15516 43726
rect 15476 43240 15528 43246
rect 15476 43182 15528 43188
rect 15488 42702 15516 43182
rect 15580 43110 15608 50118
rect 15672 49842 15700 51274
rect 15856 51066 15884 51342
rect 16028 51332 16080 51338
rect 16028 51274 16080 51280
rect 15844 51060 15896 51066
rect 15844 51002 15896 51008
rect 16040 50726 16068 51274
rect 16132 50862 16160 51410
rect 16120 50856 16172 50862
rect 16120 50798 16172 50804
rect 15844 50720 15896 50726
rect 15844 50662 15896 50668
rect 16028 50720 16080 50726
rect 16028 50662 16080 50668
rect 15660 49836 15712 49842
rect 15660 49778 15712 49784
rect 15660 49700 15712 49706
rect 15660 49642 15712 49648
rect 15568 43104 15620 43110
rect 15568 43046 15620 43052
rect 15476 42696 15528 42702
rect 15476 42638 15528 42644
rect 15568 42016 15620 42022
rect 15672 42004 15700 49642
rect 15856 49434 15884 50662
rect 16132 50522 16160 50798
rect 16120 50516 16172 50522
rect 16120 50458 16172 50464
rect 16212 50380 16264 50386
rect 16212 50322 16264 50328
rect 16028 49768 16080 49774
rect 16028 49710 16080 49716
rect 15844 49428 15896 49434
rect 15844 49370 15896 49376
rect 16040 47190 16068 49710
rect 16120 49088 16172 49094
rect 16120 49030 16172 49036
rect 16132 48754 16160 49030
rect 16120 48748 16172 48754
rect 16120 48690 16172 48696
rect 16224 48686 16252 50322
rect 16316 48890 16344 51750
rect 16396 49632 16448 49638
rect 16396 49574 16448 49580
rect 16408 49314 16436 49574
rect 16500 49434 16528 53994
rect 17052 52562 17080 56200
rect 17696 53038 17724 56200
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 17868 54188 17920 54194
rect 17868 54130 17920 54136
rect 17776 53100 17828 53106
rect 17776 53042 17828 53048
rect 17684 53032 17736 53038
rect 17684 52974 17736 52980
rect 17040 52556 17092 52562
rect 17040 52498 17092 52504
rect 16856 52488 16908 52494
rect 16856 52430 16908 52436
rect 16868 50454 16896 52430
rect 17788 52154 17816 53042
rect 17880 52154 17908 54130
rect 18340 53650 18368 56200
rect 18696 54528 18748 54534
rect 18696 54470 18748 54476
rect 18512 53984 18564 53990
rect 18512 53926 18564 53932
rect 18328 53644 18380 53650
rect 18328 53586 18380 53592
rect 18420 53440 18472 53446
rect 18420 53382 18472 53388
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17776 52148 17828 52154
rect 17776 52090 17828 52096
rect 17868 52148 17920 52154
rect 17868 52090 17920 52096
rect 17684 52012 17736 52018
rect 17684 51954 17736 51960
rect 17316 51536 17368 51542
rect 17316 51478 17368 51484
rect 17328 50998 17356 51478
rect 17408 51332 17460 51338
rect 17408 51274 17460 51280
rect 17420 51066 17448 51274
rect 17500 51264 17552 51270
rect 17500 51206 17552 51212
rect 17408 51060 17460 51066
rect 17408 51002 17460 51008
rect 17316 50992 17368 50998
rect 17316 50934 17368 50940
rect 17040 50924 17092 50930
rect 17040 50866 17092 50872
rect 16856 50448 16908 50454
rect 16856 50390 16908 50396
rect 17052 50318 17080 50866
rect 17408 50720 17460 50726
rect 17408 50662 17460 50668
rect 17420 50386 17448 50662
rect 17408 50380 17460 50386
rect 17408 50322 17460 50328
rect 17040 50312 17092 50318
rect 17040 50254 17092 50260
rect 16580 49972 16632 49978
rect 16580 49914 16632 49920
rect 16488 49428 16540 49434
rect 16488 49370 16540 49376
rect 16408 49298 16528 49314
rect 16408 49292 16540 49298
rect 16408 49286 16488 49292
rect 16304 48884 16356 48890
rect 16304 48826 16356 48832
rect 16212 48680 16264 48686
rect 16212 48622 16264 48628
rect 16408 48346 16436 49286
rect 16488 49234 16540 49240
rect 16396 48340 16448 48346
rect 16396 48282 16448 48288
rect 16212 48068 16264 48074
rect 16212 48010 16264 48016
rect 16224 47734 16252 48010
rect 16212 47728 16264 47734
rect 16212 47670 16264 47676
rect 16028 47184 16080 47190
rect 16080 47132 16160 47138
rect 16028 47126 16160 47132
rect 16040 47110 16160 47126
rect 16028 47048 16080 47054
rect 16028 46990 16080 46996
rect 16040 45558 16068 46990
rect 16132 46034 16160 47110
rect 16224 46986 16252 47670
rect 16304 47252 16356 47258
rect 16304 47194 16356 47200
rect 16212 46980 16264 46986
rect 16212 46922 16264 46928
rect 16224 46578 16252 46922
rect 16316 46714 16344 47194
rect 16396 47184 16448 47190
rect 16396 47126 16448 47132
rect 16304 46708 16356 46714
rect 16304 46650 16356 46656
rect 16212 46572 16264 46578
rect 16212 46514 16264 46520
rect 16120 46028 16172 46034
rect 16120 45970 16172 45976
rect 16028 45552 16080 45558
rect 15934 45520 15990 45529
rect 16028 45494 16080 45500
rect 15934 45455 15990 45464
rect 15948 45422 15976 45455
rect 16132 45422 16160 45970
rect 16224 45898 16252 46514
rect 16212 45892 16264 45898
rect 16212 45834 16264 45840
rect 15936 45416 15988 45422
rect 15936 45358 15988 45364
rect 16120 45416 16172 45422
rect 16120 45358 16172 45364
rect 16120 44736 16172 44742
rect 16120 44678 16172 44684
rect 16132 44402 16160 44678
rect 16120 44396 16172 44402
rect 16120 44338 16172 44344
rect 16224 43722 16252 45834
rect 16408 44946 16436 47126
rect 16592 46646 16620 49914
rect 17052 49910 17080 50254
rect 17040 49904 17092 49910
rect 17040 49846 17092 49852
rect 17052 49298 17080 49846
rect 17040 49292 17092 49298
rect 17040 49234 17092 49240
rect 16672 48612 16724 48618
rect 16672 48554 16724 48560
rect 16580 46640 16632 46646
rect 16580 46582 16632 46588
rect 16684 45558 16712 48554
rect 17052 48210 17080 49234
rect 17512 49094 17540 51206
rect 17592 50516 17644 50522
rect 17592 50458 17644 50464
rect 17604 49842 17632 50458
rect 17592 49836 17644 49842
rect 17592 49778 17644 49784
rect 17500 49088 17552 49094
rect 17500 49030 17552 49036
rect 17500 48612 17552 48618
rect 17500 48554 17552 48560
rect 17316 48544 17368 48550
rect 17316 48486 17368 48492
rect 17040 48204 17092 48210
rect 17040 48146 17092 48152
rect 16764 48000 16816 48006
rect 16764 47942 16816 47948
rect 16672 45552 16724 45558
rect 16672 45494 16724 45500
rect 16488 45484 16540 45490
rect 16488 45426 16540 45432
rect 16396 44940 16448 44946
rect 16396 44882 16448 44888
rect 15752 43716 15804 43722
rect 15752 43658 15804 43664
rect 16028 43716 16080 43722
rect 16028 43658 16080 43664
rect 16212 43716 16264 43722
rect 16212 43658 16264 43664
rect 15764 42362 15792 43658
rect 15844 43308 15896 43314
rect 15844 43250 15896 43256
rect 15752 42356 15804 42362
rect 15752 42298 15804 42304
rect 15620 41976 15700 42004
rect 15568 41958 15620 41964
rect 15384 41744 15436 41750
rect 15384 41686 15436 41692
rect 15752 41676 15804 41682
rect 15752 41618 15804 41624
rect 15764 41274 15792 41618
rect 15752 41268 15804 41274
rect 15752 41210 15804 41216
rect 14922 41032 14978 41041
rect 14922 40967 14978 40976
rect 15108 39840 15160 39846
rect 15108 39782 15160 39788
rect 14792 39528 14872 39556
rect 14740 39510 14792 39516
rect 15016 39092 15068 39098
rect 15016 39034 15068 39040
rect 14740 38888 14792 38894
rect 14740 38830 14792 38836
rect 14556 38412 14608 38418
rect 14556 38354 14608 38360
rect 14464 38208 14516 38214
rect 14464 38150 14516 38156
rect 14476 38010 14504 38150
rect 14464 38004 14516 38010
rect 14464 37946 14516 37952
rect 14476 37194 14504 37946
rect 14568 37874 14596 38354
rect 14556 37868 14608 37874
rect 14556 37810 14608 37816
rect 14556 37732 14608 37738
rect 14556 37674 14608 37680
rect 14464 37188 14516 37194
rect 14464 37130 14516 37136
rect 14464 35760 14516 35766
rect 14464 35702 14516 35708
rect 14372 34468 14424 34474
rect 14372 34410 14424 34416
rect 14280 33992 14332 33998
rect 14280 33934 14332 33940
rect 14292 33590 14320 33934
rect 14280 33584 14332 33590
rect 14476 33538 14504 35702
rect 14280 33526 14332 33532
rect 14292 32570 14320 33526
rect 14384 33510 14504 33538
rect 14280 32564 14332 32570
rect 14280 32506 14332 32512
rect 14384 29850 14412 33510
rect 14464 32564 14516 32570
rect 14464 32506 14516 32512
rect 14476 32434 14504 32506
rect 14464 32428 14516 32434
rect 14464 32370 14516 32376
rect 14568 31754 14596 37674
rect 14752 36378 14780 38830
rect 14832 38276 14884 38282
rect 14832 38218 14884 38224
rect 14844 37670 14872 38218
rect 14832 37664 14884 37670
rect 14832 37606 14884 37612
rect 14844 36718 14872 37606
rect 14832 36712 14884 36718
rect 14832 36654 14884 36660
rect 14740 36372 14792 36378
rect 14740 36314 14792 36320
rect 14648 35624 14700 35630
rect 14648 35566 14700 35572
rect 14660 35086 14688 35566
rect 14648 35080 14700 35086
rect 14648 35022 14700 35028
rect 14752 34082 14780 36314
rect 14924 35148 14976 35154
rect 14924 35090 14976 35096
rect 14832 34536 14884 34542
rect 14936 34524 14964 35090
rect 14884 34496 14964 34524
rect 14832 34478 14884 34484
rect 14660 34066 14780 34082
rect 14648 34060 14780 34066
rect 14700 34054 14780 34060
rect 14648 34002 14700 34008
rect 14646 33960 14702 33969
rect 14646 33895 14648 33904
rect 14700 33895 14702 33904
rect 14648 33866 14700 33872
rect 14660 32570 14688 33866
rect 14740 33516 14792 33522
rect 14740 33458 14792 33464
rect 14648 32564 14700 32570
rect 14648 32506 14700 32512
rect 14568 31726 14688 31754
rect 14556 31272 14608 31278
rect 14556 31214 14608 31220
rect 14568 30802 14596 31214
rect 14556 30796 14608 30802
rect 14556 30738 14608 30744
rect 14464 30728 14516 30734
rect 14464 30670 14516 30676
rect 14372 29844 14424 29850
rect 14372 29786 14424 29792
rect 14476 29646 14504 30670
rect 14660 30054 14688 31726
rect 14648 30048 14700 30054
rect 14648 29990 14700 29996
rect 14752 29646 14780 33458
rect 14844 32570 14872 34478
rect 14924 32768 14976 32774
rect 14924 32710 14976 32716
rect 14832 32564 14884 32570
rect 14832 32506 14884 32512
rect 14936 32366 14964 32710
rect 14924 32360 14976 32366
rect 14924 32302 14976 32308
rect 14924 32224 14976 32230
rect 14924 32166 14976 32172
rect 14936 32026 14964 32166
rect 14924 32020 14976 32026
rect 14924 31962 14976 31968
rect 14924 31408 14976 31414
rect 14924 31350 14976 31356
rect 14832 31272 14884 31278
rect 14832 31214 14884 31220
rect 14464 29640 14516 29646
rect 14464 29582 14516 29588
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 14740 29504 14792 29510
rect 14740 29446 14792 29452
rect 14752 28490 14780 29446
rect 14740 28484 14792 28490
rect 14740 28426 14792 28432
rect 14188 27464 14240 27470
rect 14188 27406 14240 27412
rect 13912 24404 13964 24410
rect 13912 24346 13964 24352
rect 14844 24274 14872 31214
rect 14936 30938 14964 31350
rect 14924 30932 14976 30938
rect 14924 30874 14976 30880
rect 15028 29306 15056 39034
rect 15120 38554 15148 39782
rect 15200 39500 15252 39506
rect 15200 39442 15252 39448
rect 15568 39500 15620 39506
rect 15568 39442 15620 39448
rect 15212 39302 15240 39442
rect 15200 39296 15252 39302
rect 15200 39238 15252 39244
rect 15292 39296 15344 39302
rect 15292 39238 15344 39244
rect 15108 38548 15160 38554
rect 15108 38490 15160 38496
rect 15200 37800 15252 37806
rect 15200 37742 15252 37748
rect 15108 36916 15160 36922
rect 15212 36904 15240 37742
rect 15160 36876 15240 36904
rect 15108 36858 15160 36864
rect 15200 36780 15252 36786
rect 15200 36722 15252 36728
rect 15212 34406 15240 36722
rect 15304 36650 15332 39238
rect 15476 38956 15528 38962
rect 15476 38898 15528 38904
rect 15382 38176 15438 38185
rect 15382 38111 15438 38120
rect 15396 37942 15424 38111
rect 15384 37936 15436 37942
rect 15384 37878 15436 37884
rect 15396 37194 15424 37878
rect 15384 37188 15436 37194
rect 15384 37130 15436 37136
rect 15292 36644 15344 36650
rect 15292 36586 15344 36592
rect 15396 36106 15424 37130
rect 15488 36922 15516 38898
rect 15580 38214 15608 39442
rect 15660 38752 15712 38758
rect 15660 38694 15712 38700
rect 15568 38208 15620 38214
rect 15568 38150 15620 38156
rect 15580 37330 15608 38150
rect 15568 37324 15620 37330
rect 15568 37266 15620 37272
rect 15476 36916 15528 36922
rect 15476 36858 15528 36864
rect 15384 36100 15436 36106
rect 15384 36042 15436 36048
rect 15396 34678 15424 36042
rect 15384 34672 15436 34678
rect 15384 34614 15436 34620
rect 15200 34400 15252 34406
rect 15200 34342 15252 34348
rect 15672 33658 15700 38694
rect 15856 35562 15884 43250
rect 16040 42634 16068 43658
rect 16028 42628 16080 42634
rect 15948 42588 16028 42616
rect 15948 42226 15976 42588
rect 16028 42570 16080 42576
rect 16396 42288 16448 42294
rect 16396 42230 16448 42236
rect 15936 42220 15988 42226
rect 15936 42162 15988 42168
rect 15948 41478 15976 42162
rect 16028 42084 16080 42090
rect 16028 42026 16080 42032
rect 15936 41472 15988 41478
rect 15936 41414 15988 41420
rect 15948 41138 15976 41414
rect 15936 41132 15988 41138
rect 15936 41074 15988 41080
rect 15948 40458 15976 41074
rect 15936 40452 15988 40458
rect 15936 40394 15988 40400
rect 15948 38185 15976 40394
rect 16040 38962 16068 42026
rect 16120 41472 16172 41478
rect 16120 41414 16172 41420
rect 16132 40390 16160 41414
rect 16304 41064 16356 41070
rect 16304 41006 16356 41012
rect 16120 40384 16172 40390
rect 16120 40326 16172 40332
rect 16028 38956 16080 38962
rect 16028 38898 16080 38904
rect 16120 38208 16172 38214
rect 15934 38176 15990 38185
rect 16120 38150 16172 38156
rect 15934 38111 15990 38120
rect 16132 37806 16160 38150
rect 16120 37800 16172 37806
rect 16120 37742 16172 37748
rect 16120 37324 16172 37330
rect 16120 37266 16172 37272
rect 15936 37120 15988 37126
rect 15988 37080 16068 37108
rect 15936 37062 15988 37068
rect 16040 36718 16068 37080
rect 16028 36712 16080 36718
rect 16028 36654 16080 36660
rect 16040 36242 16068 36654
rect 16028 36236 16080 36242
rect 16028 36178 16080 36184
rect 15844 35556 15896 35562
rect 15844 35498 15896 35504
rect 15936 34944 15988 34950
rect 15936 34886 15988 34892
rect 15948 34202 15976 34886
rect 16132 34746 16160 37266
rect 16212 36032 16264 36038
rect 16212 35974 16264 35980
rect 16224 35086 16252 35974
rect 16316 35290 16344 41006
rect 16408 36922 16436 42230
rect 16500 41274 16528 45426
rect 16776 45082 16804 47942
rect 17132 47592 17184 47598
rect 17132 47534 17184 47540
rect 17144 46578 17172 47534
rect 17328 47530 17356 48486
rect 17408 48204 17460 48210
rect 17408 48146 17460 48152
rect 17420 47734 17448 48146
rect 17408 47728 17460 47734
rect 17408 47670 17460 47676
rect 17316 47524 17368 47530
rect 17316 47466 17368 47472
rect 17408 47456 17460 47462
rect 17408 47398 17460 47404
rect 17420 47122 17448 47398
rect 17408 47116 17460 47122
rect 17408 47058 17460 47064
rect 17132 46572 17184 46578
rect 17132 46514 17184 46520
rect 17040 46368 17092 46374
rect 17040 46310 17092 46316
rect 16764 45076 16816 45082
rect 16764 45018 16816 45024
rect 16856 45008 16908 45014
rect 16856 44950 16908 44956
rect 16672 43648 16724 43654
rect 16672 43590 16724 43596
rect 16764 43648 16816 43654
rect 16764 43590 16816 43596
rect 16684 43110 16712 43590
rect 16672 43104 16724 43110
rect 16672 43046 16724 43052
rect 16776 42906 16804 43590
rect 16868 43194 16896 44950
rect 17052 44878 17080 46310
rect 17144 46034 17172 46514
rect 17408 46504 17460 46510
rect 17512 46492 17540 48554
rect 17460 46464 17540 46492
rect 17408 46446 17460 46452
rect 17420 46170 17448 46446
rect 17408 46164 17460 46170
rect 17408 46106 17460 46112
rect 17132 46028 17184 46034
rect 17132 45970 17184 45976
rect 17408 45484 17460 45490
rect 17408 45426 17460 45432
rect 17132 45008 17184 45014
rect 17132 44950 17184 44956
rect 17040 44872 17092 44878
rect 17040 44814 17092 44820
rect 17144 44538 17172 44950
rect 17132 44532 17184 44538
rect 17132 44474 17184 44480
rect 17224 43784 17276 43790
rect 17224 43726 17276 43732
rect 17040 43308 17092 43314
rect 17040 43250 17092 43256
rect 16868 43166 16988 43194
rect 16764 42900 16816 42906
rect 16764 42842 16816 42848
rect 16764 42220 16816 42226
rect 16764 42162 16816 42168
rect 16488 41268 16540 41274
rect 16488 41210 16540 41216
rect 16488 41132 16540 41138
rect 16488 41074 16540 41080
rect 16500 39642 16528 41074
rect 16488 39636 16540 39642
rect 16488 39578 16540 39584
rect 16488 38412 16540 38418
rect 16488 38354 16540 38360
rect 16500 37874 16528 38354
rect 16672 38276 16724 38282
rect 16672 38218 16724 38224
rect 16488 37868 16540 37874
rect 16488 37810 16540 37816
rect 16684 37670 16712 38218
rect 16672 37664 16724 37670
rect 16672 37606 16724 37612
rect 16396 36916 16448 36922
rect 16396 36858 16448 36864
rect 16580 36916 16632 36922
rect 16580 36858 16632 36864
rect 16592 35834 16620 36858
rect 16580 35828 16632 35834
rect 16580 35770 16632 35776
rect 16304 35284 16356 35290
rect 16304 35226 16356 35232
rect 16684 35154 16712 37606
rect 16672 35148 16724 35154
rect 16672 35090 16724 35096
rect 16212 35080 16264 35086
rect 16212 35022 16264 35028
rect 16212 34944 16264 34950
rect 16212 34886 16264 34892
rect 16120 34740 16172 34746
rect 16120 34682 16172 34688
rect 16224 34678 16252 34886
rect 16212 34672 16264 34678
rect 16212 34614 16264 34620
rect 16672 34536 16724 34542
rect 16672 34478 16724 34484
rect 16488 34400 16540 34406
rect 16488 34342 16540 34348
rect 15936 34196 15988 34202
rect 15936 34138 15988 34144
rect 16500 33930 16528 34342
rect 16684 33998 16712 34478
rect 16672 33992 16724 33998
rect 16672 33934 16724 33940
rect 16120 33924 16172 33930
rect 16120 33866 16172 33872
rect 16488 33924 16540 33930
rect 16488 33866 16540 33872
rect 15660 33652 15712 33658
rect 15660 33594 15712 33600
rect 15384 33516 15436 33522
rect 15384 33458 15436 33464
rect 15108 33448 15160 33454
rect 15108 33390 15160 33396
rect 15120 31482 15148 33390
rect 15292 31884 15344 31890
rect 15292 31826 15344 31832
rect 15108 31476 15160 31482
rect 15108 31418 15160 31424
rect 15120 30666 15148 31418
rect 15108 30660 15160 30666
rect 15108 30602 15160 30608
rect 15016 29300 15068 29306
rect 15016 29242 15068 29248
rect 15304 28558 15332 31826
rect 15396 30598 15424 33458
rect 15476 32768 15528 32774
rect 15476 32710 15528 32716
rect 16028 32768 16080 32774
rect 16028 32710 16080 32716
rect 15488 32609 15516 32710
rect 15474 32600 15530 32609
rect 15474 32535 15530 32544
rect 16040 31890 16068 32710
rect 16028 31884 16080 31890
rect 16028 31826 16080 31832
rect 15660 31748 15712 31754
rect 15660 31690 15712 31696
rect 15672 30938 15700 31690
rect 15660 30932 15712 30938
rect 15660 30874 15712 30880
rect 15672 30666 15700 30874
rect 15660 30660 15712 30666
rect 15660 30602 15712 30608
rect 15384 30592 15436 30598
rect 15384 30534 15436 30540
rect 16132 29714 16160 33866
rect 16684 33590 16712 33934
rect 16776 33658 16804 42162
rect 16960 39642 16988 43166
rect 17052 40118 17080 43250
rect 17236 42242 17264 43726
rect 17316 43648 17368 43654
rect 17316 43590 17368 43596
rect 17328 43382 17356 43590
rect 17316 43376 17368 43382
rect 17316 43318 17368 43324
rect 17316 43172 17368 43178
rect 17316 43114 17368 43120
rect 17328 42770 17356 43114
rect 17316 42764 17368 42770
rect 17316 42706 17368 42712
rect 17236 42214 17356 42242
rect 17224 42152 17276 42158
rect 17224 42094 17276 42100
rect 17236 41750 17264 42094
rect 17224 41744 17276 41750
rect 17224 41686 17276 41692
rect 17040 40112 17092 40118
rect 17040 40054 17092 40060
rect 16948 39636 17000 39642
rect 16948 39578 17000 39584
rect 17224 39296 17276 39302
rect 17224 39238 17276 39244
rect 16948 39092 17000 39098
rect 16948 39034 17000 39040
rect 16856 38956 16908 38962
rect 16856 38898 16908 38904
rect 16868 36786 16896 38898
rect 16960 38049 16988 39034
rect 17236 38434 17264 39238
rect 17144 38406 17264 38434
rect 16946 38040 17002 38049
rect 16946 37975 17002 37984
rect 16856 36780 16908 36786
rect 16856 36722 16908 36728
rect 16948 36780 17000 36786
rect 16948 36722 17000 36728
rect 16856 36236 16908 36242
rect 16856 36178 16908 36184
rect 16764 33652 16816 33658
rect 16764 33594 16816 33600
rect 16672 33584 16724 33590
rect 16672 33526 16724 33532
rect 16488 33516 16540 33522
rect 16488 33458 16540 33464
rect 16500 32910 16528 33458
rect 16488 32904 16540 32910
rect 16488 32846 16540 32852
rect 16868 32842 16896 36178
rect 16856 32836 16908 32842
rect 16856 32778 16908 32784
rect 16764 32020 16816 32026
rect 16764 31962 16816 31968
rect 16776 31346 16804 31962
rect 16764 31340 16816 31346
rect 16764 31282 16816 31288
rect 16776 30802 16804 31282
rect 16868 30938 16896 32778
rect 16960 32230 16988 36722
rect 17040 35556 17092 35562
rect 17040 35498 17092 35504
rect 17052 35222 17080 35498
rect 17040 35216 17092 35222
rect 17040 35158 17092 35164
rect 17144 33318 17172 38406
rect 17224 38276 17276 38282
rect 17224 38218 17276 38224
rect 17236 38185 17264 38218
rect 17222 38176 17278 38185
rect 17222 38111 17278 38120
rect 17236 37942 17264 38111
rect 17224 37936 17276 37942
rect 17224 37878 17276 37884
rect 17224 37188 17276 37194
rect 17224 37130 17276 37136
rect 17236 34678 17264 37130
rect 17328 35494 17356 42214
rect 17420 40186 17448 45426
rect 17696 43994 17724 51954
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 18432 51074 18460 53382
rect 18524 51406 18552 53926
rect 18604 51604 18656 51610
rect 18604 51546 18656 51552
rect 18512 51400 18564 51406
rect 18512 51342 18564 51348
rect 18616 51270 18644 51546
rect 18604 51264 18656 51270
rect 18604 51206 18656 51212
rect 18432 51046 18552 51074
rect 18420 50924 18472 50930
rect 18420 50866 18472 50872
rect 17776 50856 17828 50862
rect 17776 50798 17828 50804
rect 17788 50182 17816 50798
rect 18432 50250 18460 50866
rect 18420 50244 18472 50250
rect 18420 50186 18472 50192
rect 17776 50176 17828 50182
rect 17776 50118 17828 50124
rect 17788 49298 17816 50118
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 18328 49836 18380 49842
rect 18328 49778 18380 49784
rect 17776 49292 17828 49298
rect 17776 49234 17828 49240
rect 17776 49088 17828 49094
rect 17776 49030 17828 49036
rect 17788 44878 17816 49030
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 17866 48104 17922 48113
rect 17866 48039 17868 48048
rect 17920 48039 17922 48048
rect 17868 48010 17920 48016
rect 17880 47716 17908 48010
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 17960 47728 18012 47734
rect 17880 47688 17960 47716
rect 17960 47670 18012 47676
rect 17868 46980 17920 46986
rect 17868 46922 17920 46928
rect 17880 46646 17908 46922
rect 18340 46918 18368 49778
rect 18432 49162 18460 50186
rect 18524 49434 18552 51046
rect 18616 50386 18644 51206
rect 18604 50380 18656 50386
rect 18604 50322 18656 50328
rect 18708 49978 18736 54470
rect 18984 54262 19012 56200
rect 18972 54256 19024 54262
rect 18972 54198 19024 54204
rect 19628 53038 19656 56200
rect 19984 54324 20036 54330
rect 19984 54266 20036 54272
rect 19708 54188 19760 54194
rect 19708 54130 19760 54136
rect 19616 53032 19668 53038
rect 19616 52974 19668 52980
rect 18972 52012 19024 52018
rect 18972 51954 19024 51960
rect 18984 51074 19012 51954
rect 19524 51264 19576 51270
rect 19524 51206 19576 51212
rect 19616 51264 19668 51270
rect 19616 51206 19668 51212
rect 19536 51074 19564 51206
rect 18800 51046 19012 51074
rect 19352 51046 19564 51074
rect 18696 49972 18748 49978
rect 18696 49914 18748 49920
rect 18512 49428 18564 49434
rect 18512 49370 18564 49376
rect 18604 49360 18656 49366
rect 18604 49302 18656 49308
rect 18420 49156 18472 49162
rect 18420 49098 18472 49104
rect 18432 48113 18460 49098
rect 18616 48822 18644 49302
rect 18696 49156 18748 49162
rect 18696 49098 18748 49104
rect 18604 48816 18656 48822
rect 18604 48758 18656 48764
rect 18512 48748 18564 48754
rect 18512 48690 18564 48696
rect 18418 48104 18474 48113
rect 18418 48039 18474 48048
rect 18328 46912 18380 46918
rect 18328 46854 18380 46860
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 17868 46640 17920 46646
rect 17868 46582 17920 46588
rect 18420 46368 18472 46374
rect 18420 46310 18472 46316
rect 17868 45892 17920 45898
rect 17868 45834 17920 45840
rect 17776 44872 17828 44878
rect 17776 44814 17828 44820
rect 17776 44396 17828 44402
rect 17776 44338 17828 44344
rect 17684 43988 17736 43994
rect 17684 43930 17736 43936
rect 17684 43444 17736 43450
rect 17684 43386 17736 43392
rect 17592 43308 17644 43314
rect 17592 43250 17644 43256
rect 17500 42220 17552 42226
rect 17500 42162 17552 42168
rect 17512 41857 17540 42162
rect 17498 41848 17554 41857
rect 17498 41783 17554 41792
rect 17500 41744 17552 41750
rect 17500 41686 17552 41692
rect 17512 41478 17540 41686
rect 17500 41472 17552 41478
rect 17500 41414 17552 41420
rect 17500 40928 17552 40934
rect 17500 40870 17552 40876
rect 17408 40180 17460 40186
rect 17408 40122 17460 40128
rect 17512 40066 17540 40870
rect 17420 40038 17540 40066
rect 17420 37194 17448 40038
rect 17604 39658 17632 43250
rect 17696 42090 17724 43386
rect 17684 42084 17736 42090
rect 17684 42026 17736 42032
rect 17788 41414 17816 44338
rect 17880 43450 17908 45834
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 18328 45416 18380 45422
rect 18328 45358 18380 45364
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 17868 43444 17920 43450
rect 17868 43386 17920 43392
rect 18340 43382 18368 45358
rect 18432 44946 18460 46310
rect 18420 44940 18472 44946
rect 18420 44882 18472 44888
rect 18420 44328 18472 44334
rect 18420 44270 18472 44276
rect 18328 43376 18380 43382
rect 18328 43318 18380 43324
rect 17868 43104 17920 43110
rect 17868 43046 17920 43052
rect 17880 42158 17908 43046
rect 18328 42696 18380 42702
rect 18328 42638 18380 42644
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 18340 42362 18368 42638
rect 18328 42356 18380 42362
rect 18328 42298 18380 42304
rect 17868 42152 17920 42158
rect 17868 42094 17920 42100
rect 18144 42152 18196 42158
rect 18144 42094 18196 42100
rect 17960 42016 18012 42022
rect 17960 41958 18012 41964
rect 17972 41818 18000 41958
rect 17960 41812 18012 41818
rect 17960 41754 18012 41760
rect 18156 41750 18184 42094
rect 18144 41744 18196 41750
rect 18144 41686 18196 41692
rect 18236 41676 18288 41682
rect 18236 41618 18288 41624
rect 18248 41585 18276 41618
rect 18328 41608 18380 41614
rect 18234 41576 18290 41585
rect 18328 41550 18380 41556
rect 18234 41511 18290 41520
rect 17512 39630 17632 39658
rect 17696 41386 17816 41414
rect 17408 37188 17460 37194
rect 17408 37130 17460 37136
rect 17408 36712 17460 36718
rect 17408 36654 17460 36660
rect 17420 36378 17448 36654
rect 17408 36372 17460 36378
rect 17408 36314 17460 36320
rect 17408 35624 17460 35630
rect 17408 35566 17460 35572
rect 17316 35488 17368 35494
rect 17316 35430 17368 35436
rect 17420 35290 17448 35566
rect 17408 35284 17460 35290
rect 17408 35226 17460 35232
rect 17316 35012 17368 35018
rect 17316 34954 17368 34960
rect 17224 34672 17276 34678
rect 17224 34614 17276 34620
rect 17328 34474 17356 34954
rect 17420 34678 17448 35226
rect 17512 34950 17540 39630
rect 17592 39500 17644 39506
rect 17592 39442 17644 39448
rect 17604 37806 17632 39442
rect 17592 37800 17644 37806
rect 17592 37742 17644 37748
rect 17696 36582 17724 41386
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 17868 41064 17920 41070
rect 17868 41006 17920 41012
rect 17776 39568 17828 39574
rect 17776 39510 17828 39516
rect 17788 39098 17816 39510
rect 17776 39092 17828 39098
rect 17776 39034 17828 39040
rect 17880 38486 17908 41006
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 18340 40118 18368 41550
rect 18328 40112 18380 40118
rect 18328 40054 18380 40060
rect 18328 39976 18380 39982
rect 18328 39918 18380 39924
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 18234 38992 18290 39001
rect 18234 38927 18236 38936
rect 18288 38927 18290 38936
rect 18236 38898 18288 38904
rect 17868 38480 17920 38486
rect 17868 38422 17920 38428
rect 17774 38176 17830 38185
rect 17774 38111 17830 38120
rect 17788 37233 17816 38111
rect 17880 38010 17908 38422
rect 18340 38418 18368 39918
rect 18432 39642 18460 44270
rect 18524 42702 18552 48690
rect 18708 47954 18736 49098
rect 18616 47926 18736 47954
rect 18512 42696 18564 42702
rect 18512 42638 18564 42644
rect 18512 42560 18564 42566
rect 18512 42502 18564 42508
rect 18524 42362 18552 42502
rect 18512 42356 18564 42362
rect 18512 42298 18564 42304
rect 18616 42242 18644 47926
rect 18800 47784 18828 51046
rect 18972 50312 19024 50318
rect 18972 50254 19024 50260
rect 18880 49292 18932 49298
rect 18880 49234 18932 49240
rect 18892 48210 18920 49234
rect 18880 48204 18932 48210
rect 18880 48146 18932 48152
rect 18984 48006 19012 50254
rect 19352 49366 19380 51046
rect 19432 50924 19484 50930
rect 19432 50866 19484 50872
rect 19340 49360 19392 49366
rect 19340 49302 19392 49308
rect 19064 49224 19116 49230
rect 19064 49166 19116 49172
rect 18972 48000 19024 48006
rect 18972 47942 19024 47948
rect 18708 47756 18828 47784
rect 18708 44538 18736 47756
rect 18984 47598 19012 47942
rect 18972 47592 19024 47598
rect 18972 47534 19024 47540
rect 19076 47258 19104 49166
rect 19444 48770 19472 50866
rect 19524 50720 19576 50726
rect 19524 50662 19576 50668
rect 19168 48742 19472 48770
rect 19168 48686 19196 48742
rect 19156 48680 19208 48686
rect 19156 48622 19208 48628
rect 19432 48340 19484 48346
rect 19432 48282 19484 48288
rect 19248 47456 19300 47462
rect 19248 47398 19300 47404
rect 19064 47252 19116 47258
rect 19064 47194 19116 47200
rect 18788 46912 18840 46918
rect 18788 46854 18840 46860
rect 18800 45558 18828 46854
rect 19076 46510 19104 47194
rect 19260 47138 19288 47398
rect 19168 47110 19288 47138
rect 19064 46504 19116 46510
rect 19064 46446 19116 46452
rect 18788 45552 18840 45558
rect 18788 45494 18840 45500
rect 19168 45354 19196 47110
rect 19248 46980 19300 46986
rect 19248 46922 19300 46928
rect 19260 46374 19288 46922
rect 19248 46368 19300 46374
rect 19248 46310 19300 46316
rect 19340 45960 19392 45966
rect 19340 45902 19392 45908
rect 19156 45348 19208 45354
rect 19156 45290 19208 45296
rect 19248 45280 19300 45286
rect 19248 45222 19300 45228
rect 19260 44946 19288 45222
rect 19248 44940 19300 44946
rect 19248 44882 19300 44888
rect 19352 44878 19380 45902
rect 19444 45626 19472 48282
rect 19536 47802 19564 50662
rect 19628 50522 19656 51206
rect 19616 50516 19668 50522
rect 19616 50458 19668 50464
rect 19616 50176 19668 50182
rect 19616 50118 19668 50124
rect 19524 47796 19576 47802
rect 19524 47738 19576 47744
rect 19628 47138 19656 50118
rect 19720 49366 19748 54130
rect 19892 53100 19944 53106
rect 19892 53042 19944 53048
rect 19708 49360 19760 49366
rect 19708 49302 19760 49308
rect 19904 48890 19932 53042
rect 19996 51474 20024 54266
rect 20272 54126 20300 56200
rect 20536 54256 20588 54262
rect 20364 54204 20536 54210
rect 20364 54198 20588 54204
rect 20364 54194 20576 54198
rect 20352 54188 20576 54194
rect 20404 54182 20576 54188
rect 20352 54130 20404 54136
rect 20260 54120 20312 54126
rect 20260 54062 20312 54068
rect 20916 53650 20944 56200
rect 20904 53644 20956 53650
rect 20904 53586 20956 53592
rect 20812 53576 20864 53582
rect 20812 53518 20864 53524
rect 20996 53576 21048 53582
rect 20996 53518 21048 53524
rect 19984 51468 20036 51474
rect 19984 51410 20036 51416
rect 20444 51264 20496 51270
rect 20444 51206 20496 51212
rect 20168 50924 20220 50930
rect 20168 50866 20220 50872
rect 20180 50794 20208 50866
rect 20456 50862 20484 51206
rect 20824 51066 20852 53518
rect 21008 52698 21036 53518
rect 21560 53106 21588 56200
rect 22204 53582 22232 56200
rect 22560 54528 22612 54534
rect 22560 54470 22612 54476
rect 22572 54330 22600 54470
rect 22468 54324 22520 54330
rect 22468 54266 22520 54272
rect 22560 54324 22612 54330
rect 22560 54266 22612 54272
rect 22652 54324 22704 54330
rect 22652 54266 22704 54272
rect 22480 53990 22508 54266
rect 22664 54210 22692 54266
rect 22572 54182 22692 54210
rect 22848 54194 22876 56200
rect 23492 54194 23520 56200
rect 23572 54324 23624 54330
rect 23572 54266 23624 54272
rect 22836 54188 22888 54194
rect 22572 54126 22600 54182
rect 22836 54130 22888 54136
rect 23480 54188 23532 54194
rect 23480 54130 23532 54136
rect 22560 54120 22612 54126
rect 22560 54062 22612 54068
rect 22652 54120 22704 54126
rect 22652 54062 22704 54068
rect 22468 53984 22520 53990
rect 22468 53926 22520 53932
rect 22192 53576 22244 53582
rect 22192 53518 22244 53524
rect 21548 53100 21600 53106
rect 21548 53042 21600 53048
rect 21272 52896 21324 52902
rect 21272 52838 21324 52844
rect 20996 52692 21048 52698
rect 20996 52634 21048 52640
rect 21180 52488 21232 52494
rect 21180 52430 21232 52436
rect 20812 51060 20864 51066
rect 20812 51002 20864 51008
rect 20444 50856 20496 50862
rect 20444 50798 20496 50804
rect 20168 50788 20220 50794
rect 20168 50730 20220 50736
rect 20076 50516 20128 50522
rect 20076 50458 20128 50464
rect 20088 50386 20116 50458
rect 20076 50380 20128 50386
rect 20076 50322 20128 50328
rect 20088 50250 20116 50322
rect 20904 50312 20956 50318
rect 20956 50272 21036 50300
rect 20904 50254 20956 50260
rect 20076 50244 20128 50250
rect 20076 50186 20128 50192
rect 20260 50244 20312 50250
rect 20260 50186 20312 50192
rect 19892 48884 19944 48890
rect 19892 48826 19944 48832
rect 20272 48686 20300 50186
rect 21008 49978 21036 50272
rect 20996 49972 21048 49978
rect 20996 49914 21048 49920
rect 21008 49706 21036 49914
rect 20996 49700 21048 49706
rect 20996 49642 21048 49648
rect 21088 49632 21140 49638
rect 21088 49574 21140 49580
rect 21100 48890 21128 49574
rect 21088 48884 21140 48890
rect 21088 48826 21140 48832
rect 20260 48680 20312 48686
rect 20260 48622 20312 48628
rect 20720 48544 20772 48550
rect 20720 48486 20772 48492
rect 20996 48544 21048 48550
rect 20996 48486 21048 48492
rect 20536 48204 20588 48210
rect 20536 48146 20588 48152
rect 19536 47110 19656 47138
rect 19536 46186 19564 47110
rect 19616 47048 19668 47054
rect 19668 47008 19748 47036
rect 19616 46990 19668 46996
rect 19720 46714 19748 47008
rect 19708 46708 19760 46714
rect 19708 46650 19760 46656
rect 19720 46510 19748 46650
rect 19708 46504 19760 46510
rect 19708 46446 19760 46452
rect 19984 46504 20036 46510
rect 19984 46446 20036 46452
rect 19536 46158 19656 46186
rect 19524 46028 19576 46034
rect 19524 45970 19576 45976
rect 19432 45620 19484 45626
rect 19432 45562 19484 45568
rect 19340 44872 19392 44878
rect 19340 44814 19392 44820
rect 19536 44742 19564 45970
rect 19628 44810 19656 46158
rect 19720 46034 19748 46446
rect 19708 46028 19760 46034
rect 19708 45970 19760 45976
rect 19720 44946 19748 45970
rect 19996 45830 20024 46446
rect 20352 46028 20404 46034
rect 20352 45970 20404 45976
rect 19984 45824 20036 45830
rect 19984 45766 20036 45772
rect 19708 44940 19760 44946
rect 19708 44882 19760 44888
rect 19616 44804 19668 44810
rect 19616 44746 19668 44752
rect 19708 44804 19760 44810
rect 19708 44746 19760 44752
rect 19524 44736 19576 44742
rect 19524 44678 19576 44684
rect 18696 44532 18748 44538
rect 18696 44474 18748 44480
rect 19156 44396 19208 44402
rect 19156 44338 19208 44344
rect 19168 43994 19196 44338
rect 19720 44266 19748 44746
rect 19892 44464 19944 44470
rect 19892 44406 19944 44412
rect 19708 44260 19760 44266
rect 19708 44202 19760 44208
rect 19156 43988 19208 43994
rect 19156 43930 19208 43936
rect 19720 43450 19748 44202
rect 19904 43790 19932 44406
rect 19996 44334 20024 45766
rect 20364 45422 20392 45970
rect 20442 45520 20498 45529
rect 20442 45455 20498 45464
rect 20352 45416 20404 45422
rect 20352 45358 20404 45364
rect 20076 44736 20128 44742
rect 20076 44678 20128 44684
rect 19984 44328 20036 44334
rect 19984 44270 20036 44276
rect 20088 43858 20116 44678
rect 20456 44470 20484 45455
rect 20444 44464 20496 44470
rect 20444 44406 20496 44412
rect 20548 44266 20576 48146
rect 20732 47598 20760 48486
rect 21008 48142 21036 48486
rect 20996 48136 21048 48142
rect 20996 48078 21048 48084
rect 21192 48006 21220 52430
rect 21284 48822 21312 52838
rect 22664 50998 22692 54062
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 23480 53712 23532 53718
rect 23480 53654 23532 53660
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 23492 51066 23520 53654
rect 23480 51060 23532 51066
rect 23480 51002 23532 51008
rect 22652 50992 22704 50998
rect 22652 50934 22704 50940
rect 21456 50924 21508 50930
rect 21456 50866 21508 50872
rect 21548 50924 21600 50930
rect 21548 50866 21600 50872
rect 21468 50402 21496 50866
rect 21560 50522 21588 50866
rect 23296 50856 23348 50862
rect 23296 50798 23348 50804
rect 22468 50720 22520 50726
rect 22468 50662 22520 50668
rect 21548 50516 21600 50522
rect 21548 50458 21600 50464
rect 21732 50516 21784 50522
rect 21732 50458 21784 50464
rect 21376 50374 21496 50402
rect 21548 50380 21600 50386
rect 21272 48816 21324 48822
rect 21272 48758 21324 48764
rect 21272 48136 21324 48142
rect 21272 48078 21324 48084
rect 21180 48000 21232 48006
rect 21180 47942 21232 47948
rect 20996 47660 21048 47666
rect 20916 47620 20996 47648
rect 20628 47592 20680 47598
rect 20628 47534 20680 47540
rect 20720 47592 20772 47598
rect 20720 47534 20772 47540
rect 20640 47410 20668 47534
rect 20640 47382 20852 47410
rect 20824 46714 20852 47382
rect 20916 46986 20944 47620
rect 20996 47602 21048 47608
rect 20904 46980 20956 46986
rect 20904 46922 20956 46928
rect 20812 46708 20864 46714
rect 20812 46650 20864 46656
rect 20720 46640 20772 46646
rect 20720 46582 20772 46588
rect 20732 46492 20760 46582
rect 20916 46492 20944 46922
rect 20732 46464 20944 46492
rect 20824 45898 20852 46464
rect 20812 45892 20864 45898
rect 20812 45834 20864 45840
rect 20824 45286 20852 45834
rect 20812 45280 20864 45286
rect 20812 45222 20864 45228
rect 20824 44878 20852 45222
rect 20812 44872 20864 44878
rect 20812 44814 20864 44820
rect 20904 44396 20956 44402
rect 20904 44338 20956 44344
rect 20536 44260 20588 44266
rect 20536 44202 20588 44208
rect 20916 43994 20944 44338
rect 20904 43988 20956 43994
rect 20904 43930 20956 43936
rect 20076 43852 20128 43858
rect 20076 43794 20128 43800
rect 19892 43784 19944 43790
rect 19892 43726 19944 43732
rect 21284 43450 21312 48078
rect 21376 44198 21404 50374
rect 21548 50322 21600 50328
rect 21456 50244 21508 50250
rect 21456 50186 21508 50192
rect 21468 49774 21496 50186
rect 21560 49910 21588 50322
rect 21548 49904 21600 49910
rect 21548 49846 21600 49852
rect 21456 49768 21508 49774
rect 21456 49710 21508 49716
rect 21456 49632 21508 49638
rect 21456 49574 21508 49580
rect 21548 49632 21600 49638
rect 21548 49574 21600 49580
rect 21468 49298 21496 49574
rect 21560 49434 21588 49574
rect 21548 49428 21600 49434
rect 21548 49370 21600 49376
rect 21640 49428 21692 49434
rect 21640 49370 21692 49376
rect 21456 49292 21508 49298
rect 21456 49234 21508 49240
rect 21468 48822 21496 49234
rect 21456 48816 21508 48822
rect 21456 48758 21508 48764
rect 21456 48680 21508 48686
rect 21456 48622 21508 48628
rect 21468 47462 21496 48622
rect 21456 47456 21508 47462
rect 21456 47398 21508 47404
rect 21468 45354 21496 47398
rect 21652 47258 21680 49370
rect 21744 48074 21772 50458
rect 21824 49768 21876 49774
rect 21824 49710 21876 49716
rect 21732 48068 21784 48074
rect 21732 48010 21784 48016
rect 21640 47252 21692 47258
rect 21640 47194 21692 47200
rect 21652 46170 21680 47194
rect 21836 46714 21864 49710
rect 22192 49088 22244 49094
rect 22192 49030 22244 49036
rect 22204 48906 22232 49030
rect 22204 48878 22416 48906
rect 21916 48748 21968 48754
rect 21916 48690 21968 48696
rect 21928 48210 21956 48690
rect 22388 48686 22416 48878
rect 22376 48680 22428 48686
rect 22376 48622 22428 48628
rect 22480 48550 22508 50662
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22652 50380 22704 50386
rect 22652 50322 22704 50328
rect 22664 50182 22692 50322
rect 22652 50176 22704 50182
rect 22652 50118 22704 50124
rect 22664 49960 22692 50118
rect 22572 49932 22692 49960
rect 22744 49972 22796 49978
rect 22572 49298 22600 49932
rect 22744 49914 22796 49920
rect 22560 49292 22612 49298
rect 22560 49234 22612 49240
rect 22560 49088 22612 49094
rect 22560 49030 22612 49036
rect 22468 48544 22520 48550
rect 22468 48486 22520 48492
rect 22572 48210 22600 49030
rect 21916 48204 21968 48210
rect 21916 48146 21968 48152
rect 22560 48204 22612 48210
rect 22560 48146 22612 48152
rect 22284 48136 22336 48142
rect 22284 48078 22336 48084
rect 22296 47802 22324 48078
rect 22284 47796 22336 47802
rect 22284 47738 22336 47744
rect 22468 47456 22520 47462
rect 22468 47398 22520 47404
rect 22284 47048 22336 47054
rect 22284 46990 22336 46996
rect 21824 46708 21876 46714
rect 21824 46650 21876 46656
rect 22296 46510 22324 46990
rect 22284 46504 22336 46510
rect 22284 46446 22336 46452
rect 21640 46164 21692 46170
rect 21640 46106 21692 46112
rect 22296 45966 22324 46446
rect 22284 45960 22336 45966
rect 22284 45902 22336 45908
rect 22296 45422 22324 45902
rect 22284 45416 22336 45422
rect 22284 45358 22336 45364
rect 21456 45348 21508 45354
rect 21456 45290 21508 45296
rect 21640 44736 21692 44742
rect 21640 44678 21692 44684
rect 22008 44736 22060 44742
rect 22008 44678 22060 44684
rect 21364 44192 21416 44198
rect 21364 44134 21416 44140
rect 21652 43926 21680 44678
rect 22020 44402 22048 44678
rect 22008 44396 22060 44402
rect 22008 44338 22060 44344
rect 21640 43920 21692 43926
rect 21640 43862 21692 43868
rect 21824 43784 21876 43790
rect 21824 43726 21876 43732
rect 22284 43784 22336 43790
rect 22284 43726 22336 43732
rect 21836 43450 21864 43726
rect 19708 43444 19760 43450
rect 19708 43386 19760 43392
rect 21272 43444 21324 43450
rect 21272 43386 21324 43392
rect 21824 43444 21876 43450
rect 21824 43386 21876 43392
rect 20812 43308 20864 43314
rect 20812 43250 20864 43256
rect 20260 42900 20312 42906
rect 20260 42842 20312 42848
rect 19984 42764 20036 42770
rect 19984 42706 20036 42712
rect 18694 42664 18750 42673
rect 18694 42599 18696 42608
rect 18748 42599 18750 42608
rect 18696 42570 18748 42576
rect 18788 42560 18840 42566
rect 18788 42502 18840 42508
rect 18972 42560 19024 42566
rect 18972 42502 19024 42508
rect 19800 42560 19852 42566
rect 19800 42502 19852 42508
rect 18524 42214 18644 42242
rect 18524 42158 18552 42214
rect 18512 42152 18564 42158
rect 18512 42094 18564 42100
rect 18696 42152 18748 42158
rect 18696 42094 18748 42100
rect 18510 41576 18566 41585
rect 18510 41511 18566 41520
rect 18524 40497 18552 41511
rect 18510 40488 18566 40497
rect 18510 40423 18566 40432
rect 18512 40112 18564 40118
rect 18512 40054 18564 40060
rect 18420 39636 18472 39642
rect 18420 39578 18472 39584
rect 18420 39296 18472 39302
rect 18420 39238 18472 39244
rect 18432 38758 18460 39238
rect 18420 38752 18472 38758
rect 18420 38694 18472 38700
rect 18328 38412 18380 38418
rect 18328 38354 18380 38360
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 17868 38004 17920 38010
rect 17868 37946 17920 37952
rect 18418 37768 18474 37777
rect 18418 37703 18474 37712
rect 17774 37224 17830 37233
rect 17774 37159 17776 37168
rect 17828 37159 17830 37168
rect 17776 37130 17828 37136
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 18052 36848 18104 36854
rect 18052 36790 18104 36796
rect 18064 36582 18092 36790
rect 17684 36576 17736 36582
rect 17684 36518 17736 36524
rect 17776 36576 17828 36582
rect 17776 36518 17828 36524
rect 18052 36576 18104 36582
rect 18052 36518 18104 36524
rect 17788 35834 17816 36518
rect 18432 36174 18460 37703
rect 18420 36168 18472 36174
rect 18420 36110 18472 36116
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 17776 35828 17828 35834
rect 17776 35770 17828 35776
rect 17696 35686 17908 35714
rect 17500 34944 17552 34950
rect 17500 34886 17552 34892
rect 17500 34740 17552 34746
rect 17500 34682 17552 34688
rect 17408 34672 17460 34678
rect 17408 34614 17460 34620
rect 17316 34468 17368 34474
rect 17316 34410 17368 34416
rect 17132 33312 17184 33318
rect 17132 33254 17184 33260
rect 16948 32224 17000 32230
rect 16948 32166 17000 32172
rect 16856 30932 16908 30938
rect 16856 30874 16908 30880
rect 16764 30796 16816 30802
rect 16764 30738 16816 30744
rect 17328 30190 17356 34410
rect 17406 33960 17462 33969
rect 17406 33895 17408 33904
rect 17460 33895 17462 33904
rect 17408 33866 17460 33872
rect 17420 32502 17448 33866
rect 17408 32496 17460 32502
rect 17408 32438 17460 32444
rect 17512 32366 17540 34682
rect 17592 33516 17644 33522
rect 17592 33458 17644 33464
rect 17500 32360 17552 32366
rect 17420 32308 17500 32314
rect 17420 32302 17552 32308
rect 17420 32286 17540 32302
rect 17316 30184 17368 30190
rect 17316 30126 17368 30132
rect 16120 29708 16172 29714
rect 16120 29650 16172 29656
rect 15292 28552 15344 28558
rect 15292 28494 15344 28500
rect 15108 27872 15160 27878
rect 15108 27814 15160 27820
rect 14832 24268 14884 24274
rect 14832 24210 14884 24216
rect 12808 24200 12860 24206
rect 12808 24142 12860 24148
rect 13820 24200 13872 24206
rect 13820 24142 13872 24148
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12820 10470 12848 24142
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 15120 20942 15148 27814
rect 17132 27328 17184 27334
rect 17132 27270 17184 27276
rect 16212 26784 16264 26790
rect 16212 26726 16264 26732
rect 15108 20936 15160 20942
rect 15108 20878 15160 20884
rect 16224 20466 16252 26726
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 17144 17202 17172 27270
rect 17420 23662 17448 32286
rect 17500 32020 17552 32026
rect 17500 31962 17552 31968
rect 17512 31278 17540 31962
rect 17500 31272 17552 31278
rect 17500 31214 17552 31220
rect 17408 23656 17460 23662
rect 17408 23598 17460 23604
rect 17604 23322 17632 33458
rect 17696 32026 17724 35686
rect 17880 35630 17908 35686
rect 17776 35624 17828 35630
rect 17776 35566 17828 35572
rect 17868 35624 17920 35630
rect 17868 35566 17920 35572
rect 17788 33862 17816 35566
rect 18420 35488 18472 35494
rect 18420 35430 18472 35436
rect 17868 35012 17920 35018
rect 17868 34954 17920 34960
rect 17880 34660 17908 34954
rect 18328 34944 18380 34950
rect 18328 34886 18380 34892
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 17960 34672 18012 34678
rect 17880 34632 17960 34660
rect 17880 33969 17908 34632
rect 17960 34614 18012 34620
rect 17866 33960 17922 33969
rect 17866 33895 17922 33904
rect 17776 33856 17828 33862
rect 17776 33798 17828 33804
rect 17684 32020 17736 32026
rect 17684 31962 17736 31968
rect 17788 31890 17816 33798
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 18340 33658 18368 34886
rect 18328 33652 18380 33658
rect 18328 33594 18380 33600
rect 18432 33386 18460 35430
rect 18524 33658 18552 40054
rect 18708 39545 18736 42094
rect 18800 41993 18828 42502
rect 18786 41984 18842 41993
rect 18786 41919 18842 41928
rect 18788 41064 18840 41070
rect 18788 41006 18840 41012
rect 18800 40390 18828 41006
rect 18880 40452 18932 40458
rect 18880 40394 18932 40400
rect 18788 40384 18840 40390
rect 18788 40326 18840 40332
rect 18694 39536 18750 39545
rect 18694 39471 18750 39480
rect 18696 38888 18748 38894
rect 18696 38830 18748 38836
rect 18604 37936 18656 37942
rect 18604 37878 18656 37884
rect 18616 36786 18644 37878
rect 18708 37262 18736 38830
rect 18800 37942 18828 40326
rect 18892 40089 18920 40394
rect 18878 40080 18934 40089
rect 18878 40015 18934 40024
rect 18880 39976 18932 39982
rect 18880 39918 18932 39924
rect 18788 37936 18840 37942
rect 18788 37878 18840 37884
rect 18788 37800 18840 37806
rect 18788 37742 18840 37748
rect 18800 37466 18828 37742
rect 18788 37460 18840 37466
rect 18788 37402 18840 37408
rect 18892 37330 18920 39918
rect 18880 37324 18932 37330
rect 18880 37266 18932 37272
rect 18696 37256 18748 37262
rect 18696 37198 18748 37204
rect 18786 37224 18842 37233
rect 18708 37126 18736 37198
rect 18786 37159 18788 37168
rect 18840 37159 18842 37168
rect 18788 37130 18840 37136
rect 18696 37120 18748 37126
rect 18696 37062 18748 37068
rect 18708 36786 18736 37062
rect 18880 36848 18932 36854
rect 18880 36790 18932 36796
rect 18604 36780 18656 36786
rect 18604 36722 18656 36728
rect 18696 36780 18748 36786
rect 18696 36722 18748 36728
rect 18892 36718 18920 36790
rect 18788 36712 18840 36718
rect 18788 36654 18840 36660
rect 18880 36712 18932 36718
rect 18880 36654 18932 36660
rect 18800 34406 18828 36654
rect 18788 34400 18840 34406
rect 18788 34342 18840 34348
rect 18892 33844 18920 36654
rect 18984 36582 19012 42502
rect 19708 42288 19760 42294
rect 19708 42230 19760 42236
rect 19720 42022 19748 42230
rect 19812 42226 19840 42502
rect 19996 42276 20024 42706
rect 20076 42288 20128 42294
rect 19996 42248 20076 42276
rect 19800 42220 19852 42226
rect 19800 42162 19852 42168
rect 19248 42016 19300 42022
rect 19248 41958 19300 41964
rect 19708 42016 19760 42022
rect 19708 41958 19760 41964
rect 19260 41274 19288 41958
rect 19614 41440 19670 41449
rect 19614 41375 19670 41384
rect 19248 41268 19300 41274
rect 19248 41210 19300 41216
rect 19524 41200 19576 41206
rect 19524 41142 19576 41148
rect 19536 41002 19564 41142
rect 19628 41070 19656 41375
rect 19616 41064 19668 41070
rect 19616 41006 19668 41012
rect 19524 40996 19576 41002
rect 19524 40938 19576 40944
rect 19996 40730 20024 42248
rect 20076 42230 20128 42236
rect 20168 42220 20220 42226
rect 20168 42162 20220 42168
rect 19984 40724 20036 40730
rect 19984 40666 20036 40672
rect 19064 40656 19116 40662
rect 19064 40598 19116 40604
rect 19076 40118 19104 40598
rect 19708 40588 19760 40594
rect 19708 40530 19760 40536
rect 19156 40520 19208 40526
rect 19156 40462 19208 40468
rect 19168 40118 19196 40462
rect 19064 40112 19116 40118
rect 19064 40054 19116 40060
rect 19156 40112 19208 40118
rect 19156 40054 19208 40060
rect 19720 40050 19748 40530
rect 19800 40384 19852 40390
rect 19800 40326 19852 40332
rect 19708 40044 19760 40050
rect 19708 39986 19760 39992
rect 19720 39506 19748 39986
rect 19812 39574 19840 40326
rect 19984 40112 20036 40118
rect 19984 40054 20036 40060
rect 19800 39568 19852 39574
rect 19800 39510 19852 39516
rect 19708 39500 19760 39506
rect 19708 39442 19760 39448
rect 19996 39438 20024 40054
rect 19984 39432 20036 39438
rect 19984 39374 20036 39380
rect 19996 39098 20024 39374
rect 19984 39092 20036 39098
rect 19984 39034 20036 39040
rect 20180 38894 20208 42162
rect 20272 42158 20300 42842
rect 20718 42800 20774 42809
rect 20718 42735 20774 42744
rect 20352 42220 20404 42226
rect 20352 42162 20404 42168
rect 20260 42152 20312 42158
rect 20260 42094 20312 42100
rect 20364 41478 20392 42162
rect 20732 41614 20760 42735
rect 20824 41818 20852 43250
rect 21364 43240 21416 43246
rect 21364 43182 21416 43188
rect 21376 42362 21404 43182
rect 21456 42764 21508 42770
rect 21456 42706 21508 42712
rect 21732 42764 21784 42770
rect 21732 42706 21784 42712
rect 21088 42356 21140 42362
rect 21088 42298 21140 42304
rect 21364 42356 21416 42362
rect 21364 42298 21416 42304
rect 20904 42084 20956 42090
rect 20904 42026 20956 42032
rect 20812 41812 20864 41818
rect 20812 41754 20864 41760
rect 20720 41608 20772 41614
rect 20720 41550 20772 41556
rect 20916 41478 20944 42026
rect 21100 42022 21128 42298
rect 21364 42220 21416 42226
rect 21284 42180 21364 42208
rect 21088 42016 21140 42022
rect 21088 41958 21140 41964
rect 20996 41812 21048 41818
rect 20996 41754 21048 41760
rect 21008 41721 21036 41754
rect 20994 41712 21050 41721
rect 20994 41647 21050 41656
rect 20996 41608 21048 41614
rect 20996 41550 21048 41556
rect 20352 41472 20404 41478
rect 20352 41414 20404 41420
rect 20904 41472 20956 41478
rect 20904 41414 20956 41420
rect 20628 40724 20680 40730
rect 20628 40666 20680 40672
rect 20640 40390 20668 40666
rect 20916 40458 20944 41414
rect 20904 40452 20956 40458
rect 20904 40394 20956 40400
rect 20352 40384 20404 40390
rect 20352 40326 20404 40332
rect 20628 40384 20680 40390
rect 20628 40326 20680 40332
rect 20364 39370 20392 40326
rect 20720 40180 20772 40186
rect 20720 40122 20772 40128
rect 20352 39364 20404 39370
rect 20352 39306 20404 39312
rect 19248 38888 19300 38894
rect 19248 38830 19300 38836
rect 19892 38888 19944 38894
rect 19892 38830 19944 38836
rect 20168 38888 20220 38894
rect 20168 38830 20220 38836
rect 19260 38758 19288 38830
rect 19156 38752 19208 38758
rect 19156 38694 19208 38700
rect 19248 38752 19300 38758
rect 19248 38694 19300 38700
rect 19430 38720 19486 38729
rect 19064 38548 19116 38554
rect 19064 38490 19116 38496
rect 18972 36576 19024 36582
rect 18972 36518 19024 36524
rect 19076 36310 19104 38490
rect 19064 36304 19116 36310
rect 19064 36246 19116 36252
rect 19076 35034 19104 36246
rect 18708 33816 18920 33844
rect 18984 35006 19104 35034
rect 18512 33652 18564 33658
rect 18512 33594 18564 33600
rect 18420 33380 18472 33386
rect 18420 33322 18472 33328
rect 17868 32836 17920 32842
rect 17868 32778 17920 32784
rect 17880 32366 17908 32778
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 18420 32564 18472 32570
rect 18420 32506 18472 32512
rect 17868 32360 17920 32366
rect 17868 32302 17920 32308
rect 17880 32230 17908 32302
rect 17868 32224 17920 32230
rect 17868 32166 17920 32172
rect 17776 31884 17828 31890
rect 17776 31826 17828 31832
rect 17880 31414 17908 32166
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 18432 31414 18460 32506
rect 17868 31408 17920 31414
rect 17868 31350 17920 31356
rect 18420 31408 18472 31414
rect 18420 31350 18472 31356
rect 18328 31272 18380 31278
rect 18328 31214 18380 31220
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17592 23316 17644 23322
rect 17592 23258 17644 23264
rect 18340 23186 18368 31214
rect 18708 27402 18736 33816
rect 18788 33516 18840 33522
rect 18788 33458 18840 33464
rect 18696 27396 18748 27402
rect 18696 27338 18748 27344
rect 18800 23866 18828 33458
rect 18984 32774 19012 35006
rect 19064 34060 19116 34066
rect 19064 34002 19116 34008
rect 19076 33454 19104 34002
rect 19064 33448 19116 33454
rect 19064 33390 19116 33396
rect 18972 32768 19024 32774
rect 18972 32710 19024 32716
rect 19076 32570 19104 33390
rect 19168 33114 19196 38694
rect 19156 33108 19208 33114
rect 19156 33050 19208 33056
rect 19260 32978 19288 38694
rect 19430 38655 19486 38664
rect 19340 36848 19392 36854
rect 19340 36790 19392 36796
rect 19352 36310 19380 36790
rect 19340 36304 19392 36310
rect 19340 36246 19392 36252
rect 19444 35834 19472 38655
rect 19432 35828 19484 35834
rect 19432 35770 19484 35776
rect 19340 35556 19392 35562
rect 19340 35498 19392 35504
rect 19352 35222 19380 35498
rect 19708 35488 19760 35494
rect 19708 35430 19760 35436
rect 19340 35216 19392 35222
rect 19340 35158 19392 35164
rect 19720 35154 19748 35430
rect 19708 35148 19760 35154
rect 19708 35090 19760 35096
rect 19720 34610 19748 35090
rect 19708 34604 19760 34610
rect 19708 34546 19760 34552
rect 19720 33930 19748 34546
rect 19708 33924 19760 33930
rect 19708 33866 19760 33872
rect 19432 33516 19484 33522
rect 19432 33458 19484 33464
rect 19248 32972 19300 32978
rect 19248 32914 19300 32920
rect 19064 32564 19116 32570
rect 19064 32506 19116 32512
rect 19444 31482 19472 33458
rect 19524 32836 19576 32842
rect 19524 32778 19576 32784
rect 19432 31476 19484 31482
rect 19432 31418 19484 31424
rect 18788 23860 18840 23866
rect 18788 23802 18840 23808
rect 18328 23180 18380 23186
rect 18328 23122 18380 23128
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 19156 21072 19208 21078
rect 19156 21014 19208 21020
rect 18604 20800 18656 20806
rect 18604 20742 18656 20748
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 15856 7886 15884 17070
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 17236 6798 17264 13806
rect 17788 8974 17816 16934
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 17880 13870 17908 14962
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 18616 13938 18644 20742
rect 18696 20256 18748 20262
rect 18696 20198 18748 20204
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18708 12918 18736 20198
rect 18696 12912 18748 12918
rect 18696 12854 18748 12860
rect 19168 12850 19196 21014
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19156 12844 19208 12850
rect 19156 12786 19208 12792
rect 19352 12782 19380 13126
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 15292 6724 15344 6730
rect 15292 6666 15344 6672
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 15212 2514 15240 6054
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 10692 2304 10744 2310
rect 10692 2246 10744 2252
rect 12176 800 12204 2450
rect 15304 2378 15332 6666
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 19352 6390 19380 12718
rect 19432 8900 19484 8906
rect 19432 8842 19484 8848
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 18328 5568 18380 5574
rect 18328 5510 18380 5516
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15292 2372 15344 2378
rect 15292 2314 15344 2320
rect 15488 800 15516 2450
rect 18340 2446 18368 5510
rect 18788 2508 18840 2514
rect 18788 2450 18840 2456
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18800 800 18828 2450
rect 19444 2446 19472 8842
rect 19536 2854 19564 32778
rect 19708 32224 19760 32230
rect 19708 32166 19760 32172
rect 19720 13938 19748 32166
rect 19904 28422 19932 38830
rect 20536 38344 20588 38350
rect 20536 38286 20588 38292
rect 20548 37806 20576 38286
rect 20732 37942 20760 40122
rect 20720 37936 20772 37942
rect 20720 37878 20772 37884
rect 20168 37800 20220 37806
rect 20168 37742 20220 37748
rect 20536 37800 20588 37806
rect 20536 37742 20588 37748
rect 20180 37262 20208 37742
rect 20168 37256 20220 37262
rect 20168 37198 20220 37204
rect 20180 36242 20208 37198
rect 20812 37188 20864 37194
rect 20812 37130 20864 37136
rect 20720 37120 20772 37126
rect 20720 37062 20772 37068
rect 20732 36854 20760 37062
rect 20720 36848 20772 36854
rect 20720 36790 20772 36796
rect 20168 36236 20220 36242
rect 20168 36178 20220 36184
rect 20732 36106 20760 36790
rect 20824 36582 20852 37130
rect 20812 36576 20864 36582
rect 20812 36518 20864 36524
rect 20444 36100 20496 36106
rect 20444 36042 20496 36048
rect 20720 36100 20772 36106
rect 20720 36042 20772 36048
rect 20456 33522 20484 36042
rect 20732 35766 20760 36042
rect 20720 35760 20772 35766
rect 20720 35702 20772 35708
rect 20628 35148 20680 35154
rect 20628 35090 20680 35096
rect 20444 33516 20496 33522
rect 20444 33458 20496 33464
rect 20640 32570 20668 35090
rect 20732 34678 20760 35702
rect 20720 34672 20772 34678
rect 20720 34614 20772 34620
rect 20732 33912 20760 34614
rect 20812 33924 20864 33930
rect 20732 33884 20812 33912
rect 20628 32564 20680 32570
rect 20628 32506 20680 32512
rect 20640 31278 20668 32506
rect 20732 32434 20760 33884
rect 20812 33866 20864 33872
rect 20720 32428 20772 32434
rect 20720 32370 20772 32376
rect 20628 31272 20680 31278
rect 20628 31214 20680 31220
rect 19892 28416 19944 28422
rect 19892 28358 19944 28364
rect 20732 17270 20760 32370
rect 21008 28082 21036 41550
rect 21284 41478 21312 42180
rect 21364 42162 21416 42168
rect 21468 42158 21496 42706
rect 21744 42566 21772 42706
rect 21732 42560 21784 42566
rect 21732 42502 21784 42508
rect 21916 42560 21968 42566
rect 21916 42502 21968 42508
rect 21824 42356 21876 42362
rect 21824 42298 21876 42304
rect 21456 42152 21508 42158
rect 21456 42094 21508 42100
rect 21272 41472 21324 41478
rect 21272 41414 21324 41420
rect 21364 41472 21416 41478
rect 21364 41414 21416 41420
rect 21468 41414 21496 42094
rect 21640 41472 21692 41478
rect 21640 41414 21692 41420
rect 21272 40452 21324 40458
rect 21272 40394 21324 40400
rect 21284 40118 21312 40394
rect 21272 40112 21324 40118
rect 21272 40054 21324 40060
rect 21284 39370 21312 40054
rect 21272 39364 21324 39370
rect 21272 39306 21324 39312
rect 21284 39030 21312 39306
rect 21272 39024 21324 39030
rect 21272 38966 21324 38972
rect 21284 38282 21312 38966
rect 21376 38729 21404 41414
rect 21468 41386 21588 41414
rect 21560 40526 21588 41386
rect 21548 40520 21600 40526
rect 21548 40462 21600 40468
rect 21456 40112 21508 40118
rect 21456 40054 21508 40060
rect 21468 39846 21496 40054
rect 21560 39982 21588 40462
rect 21548 39976 21600 39982
rect 21548 39918 21600 39924
rect 21456 39840 21508 39846
rect 21456 39782 21508 39788
rect 21362 38720 21418 38729
rect 21362 38655 21418 38664
rect 21468 38418 21496 39782
rect 21652 39302 21680 41414
rect 21836 40594 21864 42298
rect 21928 42294 21956 42502
rect 21916 42288 21968 42294
rect 21916 42230 21968 42236
rect 22296 42226 22324 43726
rect 22480 43450 22508 47398
rect 22652 46504 22704 46510
rect 22652 46446 22704 46452
rect 22664 45830 22692 46446
rect 22652 45824 22704 45830
rect 22652 45766 22704 45772
rect 22664 44946 22692 45766
rect 22756 45082 22784 49914
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 23204 49156 23256 49162
rect 23204 49098 23256 49104
rect 23216 48634 23244 49098
rect 23308 48890 23336 50798
rect 23388 50312 23440 50318
rect 23388 50254 23440 50260
rect 23400 49230 23428 50254
rect 23584 50250 23612 54266
rect 24136 54194 24164 56200
rect 24780 54210 24808 56200
rect 24780 54194 24900 54210
rect 25424 54194 25452 56200
rect 26068 54210 26096 56200
rect 26068 54194 26280 54210
rect 26712 54194 26740 56200
rect 27356 55026 27384 56200
rect 27356 54998 27660 55026
rect 27632 54194 27660 54998
rect 27712 54664 27764 54670
rect 28000 54618 28028 56200
rect 27712 54606 27764 54612
rect 27724 54330 27752 54606
rect 27816 54590 28028 54618
rect 27712 54324 27764 54330
rect 27712 54266 27764 54272
rect 24124 54188 24176 54194
rect 24780 54188 24912 54194
rect 24780 54182 24860 54188
rect 24124 54130 24176 54136
rect 24860 54130 24912 54136
rect 25412 54188 25464 54194
rect 26068 54188 26292 54194
rect 26068 54182 26240 54188
rect 25412 54130 25464 54136
rect 26240 54130 26292 54136
rect 26700 54188 26752 54194
rect 26700 54130 26752 54136
rect 27620 54188 27672 54194
rect 27620 54130 27672 54136
rect 27160 53984 27212 53990
rect 27160 53926 27212 53932
rect 24860 53508 24912 53514
rect 24860 53450 24912 53456
rect 24768 50788 24820 50794
rect 24768 50730 24820 50736
rect 23572 50244 23624 50250
rect 23572 50186 23624 50192
rect 23664 50176 23716 50182
rect 23664 50118 23716 50124
rect 23388 49224 23440 49230
rect 23388 49166 23440 49172
rect 23296 48884 23348 48890
rect 23296 48826 23348 48832
rect 23400 48754 23428 49166
rect 23388 48748 23440 48754
rect 23388 48690 23440 48696
rect 23216 48606 23336 48634
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 22836 45416 22888 45422
rect 22836 45358 22888 45364
rect 22744 45076 22796 45082
rect 22744 45018 22796 45024
rect 22652 44940 22704 44946
rect 22652 44882 22704 44888
rect 22848 44402 22876 45358
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 23308 44538 23336 48606
rect 23400 48090 23428 48690
rect 23676 48686 23704 50118
rect 24780 49162 24808 50730
rect 24872 50318 24900 53450
rect 25044 53440 25096 53446
rect 25044 53382 25096 53388
rect 25056 53174 25084 53382
rect 25044 53168 25096 53174
rect 25044 53110 25096 53116
rect 26148 50924 26200 50930
rect 26148 50866 26200 50872
rect 24952 50720 25004 50726
rect 24952 50662 25004 50668
rect 24860 50312 24912 50318
rect 24860 50254 24912 50260
rect 24860 49836 24912 49842
rect 24964 49824 24992 50662
rect 24912 49796 24992 49824
rect 24860 49778 24912 49784
rect 24768 49156 24820 49162
rect 24768 49098 24820 49104
rect 24872 48754 24900 49778
rect 26056 49292 26108 49298
rect 26056 49234 26108 49240
rect 25504 49088 25556 49094
rect 25504 49030 25556 49036
rect 25872 49088 25924 49094
rect 25872 49030 25924 49036
rect 24860 48748 24912 48754
rect 24860 48690 24912 48696
rect 23664 48680 23716 48686
rect 23664 48622 23716 48628
rect 24768 48680 24820 48686
rect 24768 48622 24820 48628
rect 23400 48074 23612 48090
rect 23400 48068 23624 48074
rect 23400 48062 23572 48068
rect 23572 48010 23624 48016
rect 23584 47734 23612 48010
rect 23572 47728 23624 47734
rect 23572 47670 23624 47676
rect 23584 46986 23612 47670
rect 23572 46980 23624 46986
rect 23572 46922 23624 46928
rect 23584 46714 23612 46922
rect 23572 46708 23624 46714
rect 23572 46650 23624 46656
rect 23584 45898 23612 46650
rect 23676 46458 23704 48622
rect 24780 47598 24808 48622
rect 24952 48544 25004 48550
rect 24952 48486 25004 48492
rect 24860 48272 24912 48278
rect 24860 48214 24912 48220
rect 24032 47592 24084 47598
rect 24032 47534 24084 47540
rect 24768 47592 24820 47598
rect 24768 47534 24820 47540
rect 24044 47258 24072 47534
rect 24308 47524 24360 47530
rect 24308 47466 24360 47472
rect 24032 47252 24084 47258
rect 24032 47194 24084 47200
rect 24320 46714 24348 47466
rect 24308 46708 24360 46714
rect 24308 46650 24360 46656
rect 23676 46430 23796 46458
rect 23572 45892 23624 45898
rect 23572 45834 23624 45840
rect 23584 45558 23612 45834
rect 23768 45626 23796 46430
rect 24032 46436 24084 46442
rect 24032 46378 24084 46384
rect 23756 45620 23808 45626
rect 23756 45562 23808 45568
rect 23572 45552 23624 45558
rect 23768 45529 23796 45562
rect 23572 45494 23624 45500
rect 23754 45520 23810 45529
rect 23584 45286 23612 45494
rect 23754 45455 23810 45464
rect 23572 45280 23624 45286
rect 23572 45222 23624 45228
rect 23296 44532 23348 44538
rect 23296 44474 23348 44480
rect 23584 44470 23612 45222
rect 23664 44804 23716 44810
rect 23664 44746 23716 44752
rect 23572 44464 23624 44470
rect 23572 44406 23624 44412
rect 22836 44396 22888 44402
rect 22836 44338 22888 44344
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 23572 43852 23624 43858
rect 23572 43794 23624 43800
rect 22468 43444 22520 43450
rect 22468 43386 22520 43392
rect 23584 43246 23612 43794
rect 23572 43240 23624 43246
rect 23572 43182 23624 43188
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 22928 42764 22980 42770
rect 22928 42706 22980 42712
rect 22468 42628 22520 42634
rect 22468 42570 22520 42576
rect 22284 42220 22336 42226
rect 22284 42162 22336 42168
rect 22376 42084 22428 42090
rect 22376 42026 22428 42032
rect 22388 41818 22416 42026
rect 22376 41812 22428 41818
rect 22376 41754 22428 41760
rect 22100 41676 22152 41682
rect 22100 41618 22152 41624
rect 21824 40588 21876 40594
rect 21824 40530 21876 40536
rect 21916 39840 21968 39846
rect 21916 39782 21968 39788
rect 21732 39568 21784 39574
rect 21732 39510 21784 39516
rect 21640 39296 21692 39302
rect 21640 39238 21692 39244
rect 21640 38820 21692 38826
rect 21640 38762 21692 38768
rect 21456 38412 21508 38418
rect 21456 38354 21508 38360
rect 21272 38276 21324 38282
rect 21272 38218 21324 38224
rect 21284 37194 21312 38218
rect 21364 37664 21416 37670
rect 21364 37606 21416 37612
rect 21272 37188 21324 37194
rect 21272 37130 21324 37136
rect 21180 37120 21232 37126
rect 21180 37062 21232 37068
rect 21192 35086 21220 37062
rect 21180 35080 21232 35086
rect 21180 35022 21232 35028
rect 21376 35018 21404 37606
rect 21456 37324 21508 37330
rect 21456 37266 21508 37272
rect 21364 35012 21416 35018
rect 21364 34954 21416 34960
rect 21272 34944 21324 34950
rect 21272 34886 21324 34892
rect 21284 33658 21312 34886
rect 21468 34202 21496 37266
rect 21548 36644 21600 36650
rect 21548 36586 21600 36592
rect 21560 35494 21588 36586
rect 21548 35488 21600 35494
rect 21548 35430 21600 35436
rect 21560 34542 21588 35430
rect 21652 35086 21680 38762
rect 21744 35154 21772 39510
rect 21928 39506 21956 39782
rect 22112 39506 22140 41618
rect 22192 41540 22244 41546
rect 22192 41482 22244 41488
rect 22204 41206 22232 41482
rect 22480 41414 22508 42570
rect 22940 42294 22968 42706
rect 22928 42288 22980 42294
rect 22928 42230 22980 42236
rect 22652 42152 22704 42158
rect 22652 42094 22704 42100
rect 22664 41750 22692 42094
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 22652 41744 22704 41750
rect 22652 41686 22704 41692
rect 23572 41676 23624 41682
rect 23572 41618 23624 41624
rect 22296 41386 22508 41414
rect 22192 41200 22244 41206
rect 22192 41142 22244 41148
rect 21916 39500 21968 39506
rect 21916 39442 21968 39448
rect 22100 39500 22152 39506
rect 22100 39442 22152 39448
rect 21928 36310 21956 39442
rect 22112 38758 22140 39442
rect 22204 39386 22232 41142
rect 22296 40458 22324 41386
rect 23204 41200 23256 41206
rect 23204 41142 23256 41148
rect 23216 40934 23244 41142
rect 23388 41132 23440 41138
rect 23388 41074 23440 41080
rect 22652 40928 22704 40934
rect 22652 40870 22704 40876
rect 23204 40928 23256 40934
rect 23204 40870 23256 40876
rect 22284 40452 22336 40458
rect 22284 40394 22336 40400
rect 22204 39358 22324 39386
rect 22192 39296 22244 39302
rect 22192 39238 22244 39244
rect 22100 38752 22152 38758
rect 22100 38694 22152 38700
rect 22008 37936 22060 37942
rect 22008 37878 22060 37884
rect 21916 36304 21968 36310
rect 21916 36246 21968 36252
rect 22020 35766 22048 37878
rect 22204 36378 22232 39238
rect 22296 38214 22324 39358
rect 22560 38888 22612 38894
rect 22560 38830 22612 38836
rect 22284 38208 22336 38214
rect 22284 38150 22336 38156
rect 22376 38208 22428 38214
rect 22376 38150 22428 38156
rect 22296 38010 22324 38150
rect 22284 38004 22336 38010
rect 22284 37946 22336 37952
rect 22284 37460 22336 37466
rect 22284 37402 22336 37408
rect 22192 36372 22244 36378
rect 22192 36314 22244 36320
rect 22296 35834 22324 37402
rect 22388 36922 22416 38150
rect 22376 36916 22428 36922
rect 22376 36858 22428 36864
rect 22284 35828 22336 35834
rect 22284 35770 22336 35776
rect 22008 35760 22060 35766
rect 22008 35702 22060 35708
rect 21732 35148 21784 35154
rect 21732 35090 21784 35096
rect 21824 35148 21876 35154
rect 21824 35090 21876 35096
rect 21640 35080 21692 35086
rect 21640 35022 21692 35028
rect 21836 34746 21864 35090
rect 21824 34740 21876 34746
rect 21824 34682 21876 34688
rect 21548 34536 21600 34542
rect 21548 34478 21600 34484
rect 21456 34196 21508 34202
rect 21456 34138 21508 34144
rect 21272 33652 21324 33658
rect 21272 33594 21324 33600
rect 21468 32366 21496 34138
rect 22020 33114 22048 35702
rect 22572 34474 22600 38830
rect 22664 36922 22692 40870
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 22836 40384 22888 40390
rect 22836 40326 22888 40332
rect 23296 40384 23348 40390
rect 23296 40326 23348 40332
rect 22744 39500 22796 39506
rect 22744 39442 22796 39448
rect 22756 38554 22784 39442
rect 22744 38548 22796 38554
rect 22744 38490 22796 38496
rect 22848 38350 22876 40326
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 23308 39506 23336 40326
rect 23296 39500 23348 39506
rect 23296 39442 23348 39448
rect 23308 38894 23336 39442
rect 23296 38888 23348 38894
rect 23296 38830 23348 38836
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 22836 38344 22888 38350
rect 22836 38286 22888 38292
rect 22848 37262 22876 38286
rect 23400 38010 23428 41074
rect 23480 40996 23532 41002
rect 23480 40938 23532 40944
rect 23492 40458 23520 40938
rect 23480 40452 23532 40458
rect 23480 40394 23532 40400
rect 23480 40044 23532 40050
rect 23480 39986 23532 39992
rect 23492 38962 23520 39986
rect 23584 39846 23612 41618
rect 23676 41614 23704 44746
rect 23848 44464 23900 44470
rect 23848 44406 23900 44412
rect 23860 43722 23888 44406
rect 24044 43994 24072 46378
rect 24320 45422 24348 46650
rect 24780 46034 24808 47534
rect 24872 47122 24900 48214
rect 24860 47116 24912 47122
rect 24860 47058 24912 47064
rect 24768 46028 24820 46034
rect 24768 45970 24820 45976
rect 24308 45416 24360 45422
rect 24308 45358 24360 45364
rect 24584 45280 24636 45286
rect 24584 45222 24636 45228
rect 24032 43988 24084 43994
rect 24032 43930 24084 43936
rect 23848 43716 23900 43722
rect 23848 43658 23900 43664
rect 23860 42634 23888 43658
rect 24044 42906 24072 43930
rect 24596 43858 24624 45222
rect 24964 44878 24992 48486
rect 25516 48346 25544 49030
rect 25504 48340 25556 48346
rect 25504 48282 25556 48288
rect 25884 48142 25912 49030
rect 26068 48278 26096 49234
rect 26056 48272 26108 48278
rect 26056 48214 26108 48220
rect 25872 48136 25924 48142
rect 25872 48078 25924 48084
rect 25780 48000 25832 48006
rect 25780 47942 25832 47948
rect 25412 46572 25464 46578
rect 25412 46514 25464 46520
rect 25136 46368 25188 46374
rect 25136 46310 25188 46316
rect 24952 44872 25004 44878
rect 24952 44814 25004 44820
rect 24952 43988 25004 43994
rect 24952 43930 25004 43936
rect 24860 43920 24912 43926
rect 24860 43862 24912 43868
rect 24584 43852 24636 43858
rect 24584 43794 24636 43800
rect 24584 43648 24636 43654
rect 24584 43590 24636 43596
rect 24596 43382 24624 43590
rect 24584 43376 24636 43382
rect 24584 43318 24636 43324
rect 24032 42900 24084 42906
rect 24032 42842 24084 42848
rect 23848 42628 23900 42634
rect 23848 42570 23900 42576
rect 23860 42242 23888 42570
rect 23768 42226 23888 42242
rect 23756 42220 23888 42226
rect 23808 42214 23888 42220
rect 23756 42162 23808 42168
rect 24676 42084 24728 42090
rect 24676 42026 24728 42032
rect 23848 41676 23900 41682
rect 23848 41618 23900 41624
rect 23664 41608 23716 41614
rect 23664 41550 23716 41556
rect 23676 40730 23704 41550
rect 23756 41472 23808 41478
rect 23754 41440 23756 41449
rect 23808 41440 23810 41449
rect 23754 41375 23810 41384
rect 23860 41070 23888 41618
rect 24492 41540 24544 41546
rect 24492 41482 24544 41488
rect 24504 41274 24532 41482
rect 24400 41268 24452 41274
rect 24400 41210 24452 41216
rect 24492 41268 24544 41274
rect 24492 41210 24544 41216
rect 23940 41132 23992 41138
rect 23940 41074 23992 41080
rect 23848 41064 23900 41070
rect 23848 41006 23900 41012
rect 23664 40724 23716 40730
rect 23664 40666 23716 40672
rect 23756 40520 23808 40526
rect 23756 40462 23808 40468
rect 23664 40452 23716 40458
rect 23664 40394 23716 40400
rect 23572 39840 23624 39846
rect 23572 39782 23624 39788
rect 23572 39296 23624 39302
rect 23676 39284 23704 40394
rect 23768 39302 23796 40462
rect 23848 39976 23900 39982
rect 23848 39918 23900 39924
rect 23860 39846 23888 39918
rect 23848 39840 23900 39846
rect 23848 39782 23900 39788
rect 23624 39256 23704 39284
rect 23756 39296 23808 39302
rect 23572 39238 23624 39244
rect 23756 39238 23808 39244
rect 23480 38956 23532 38962
rect 23480 38898 23532 38904
rect 23388 38004 23440 38010
rect 23388 37946 23440 37952
rect 23296 37800 23348 37806
rect 23296 37742 23348 37748
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 23308 37330 23336 37742
rect 23296 37324 23348 37330
rect 23296 37266 23348 37272
rect 22836 37256 22888 37262
rect 22836 37198 22888 37204
rect 22652 36916 22704 36922
rect 22652 36858 22704 36864
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 23400 36106 23428 37946
rect 23492 37913 23520 38898
rect 23572 38344 23624 38350
rect 23572 38286 23624 38292
rect 23478 37904 23534 37913
rect 23478 37839 23534 37848
rect 23584 37262 23612 38286
rect 23572 37256 23624 37262
rect 23572 37198 23624 37204
rect 23584 36786 23612 37198
rect 23572 36780 23624 36786
rect 23572 36722 23624 36728
rect 23388 36100 23440 36106
rect 23388 36042 23440 36048
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 23768 35222 23796 39238
rect 23860 39098 23888 39782
rect 23848 39092 23900 39098
rect 23848 39034 23900 39040
rect 23952 38418 23980 41074
rect 24412 40730 24440 41210
rect 24400 40724 24452 40730
rect 24400 40666 24452 40672
rect 24308 39840 24360 39846
rect 24308 39782 24360 39788
rect 24320 39438 24348 39782
rect 24308 39432 24360 39438
rect 24308 39374 24360 39380
rect 23940 38412 23992 38418
rect 23940 38354 23992 38360
rect 23952 37466 23980 38354
rect 24412 38350 24440 40666
rect 24584 40384 24636 40390
rect 24584 40326 24636 40332
rect 24596 39370 24624 40326
rect 24688 40050 24716 42026
rect 24872 41750 24900 43862
rect 24964 41818 24992 43930
rect 25148 42702 25176 46310
rect 25424 45626 25452 46514
rect 25412 45620 25464 45626
rect 25412 45562 25464 45568
rect 25228 44192 25280 44198
rect 25228 44134 25280 44140
rect 25240 43858 25268 44134
rect 25228 43852 25280 43858
rect 25228 43794 25280 43800
rect 25136 42696 25188 42702
rect 25136 42638 25188 42644
rect 25240 42158 25268 43794
rect 25228 42152 25280 42158
rect 25228 42094 25280 42100
rect 24952 41812 25004 41818
rect 24952 41754 25004 41760
rect 24860 41744 24912 41750
rect 24860 41686 24912 41692
rect 24872 41274 24900 41686
rect 24964 41274 24992 41754
rect 24860 41268 24912 41274
rect 24860 41210 24912 41216
rect 24952 41268 25004 41274
rect 24952 41210 25004 41216
rect 24768 40588 24820 40594
rect 24768 40530 24820 40536
rect 24780 40118 24808 40530
rect 24768 40112 24820 40118
rect 24768 40054 24820 40060
rect 24676 40044 24728 40050
rect 24676 39986 24728 39992
rect 24584 39364 24636 39370
rect 24584 39306 24636 39312
rect 24400 38344 24452 38350
rect 24400 38286 24452 38292
rect 23940 37460 23992 37466
rect 23940 37402 23992 37408
rect 24124 35624 24176 35630
rect 24124 35566 24176 35572
rect 23756 35216 23808 35222
rect 23756 35158 23808 35164
rect 22560 34468 22612 34474
rect 22560 34410 22612 34416
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 22008 33108 22060 33114
rect 22008 33050 22060 33056
rect 21456 32360 21508 32366
rect 21456 32302 21508 32308
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 20996 28076 21048 28082
rect 20996 28018 21048 28024
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 24136 24750 24164 35566
rect 24124 24744 24176 24750
rect 24124 24686 24176 24692
rect 24676 24744 24728 24750
rect 24676 24686 24728 24692
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23572 20256 23624 20262
rect 23572 20198 23624 20204
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20732 14006 20760 17206
rect 23584 17202 23612 20198
rect 24492 17536 24544 17542
rect 24492 17478 24544 17484
rect 23572 17196 23624 17202
rect 23572 17138 23624 17144
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 23584 16590 23612 17138
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 24504 15162 24532 17478
rect 24688 17202 24716 24686
rect 25424 17746 25452 45562
rect 25792 43654 25820 47942
rect 26160 47666 26188 50866
rect 27172 49638 27200 53926
rect 27816 53582 27844 54590
rect 27950 54428 28258 54437
rect 27950 54426 27956 54428
rect 28012 54426 28036 54428
rect 28092 54426 28116 54428
rect 28172 54426 28196 54428
rect 28252 54426 28258 54428
rect 28012 54374 28014 54426
rect 28194 54374 28196 54426
rect 27950 54372 27956 54374
rect 28012 54372 28036 54374
rect 28092 54372 28116 54374
rect 28172 54372 28196 54374
rect 28252 54372 28258 54374
rect 27950 54363 28258 54372
rect 28644 54262 28672 56200
rect 28908 54732 28960 54738
rect 28908 54674 28960 54680
rect 28920 54330 28948 54674
rect 28908 54324 28960 54330
rect 28908 54266 28960 54272
rect 29288 54262 29316 56200
rect 29932 56114 29960 56200
rect 30024 56114 30052 56222
rect 29932 56086 30052 56114
rect 28632 54256 28684 54262
rect 28632 54198 28684 54204
rect 29276 54256 29328 54262
rect 29276 54198 29328 54204
rect 30300 54210 30328 56222
rect 30562 56200 30618 57000
rect 31206 56200 31262 57000
rect 31850 56200 31906 57000
rect 32494 56200 32550 57000
rect 33138 56200 33194 57000
rect 33782 56200 33838 57000
rect 34426 56200 34482 57000
rect 35070 56200 35126 57000
rect 35714 56200 35770 57000
rect 36358 56200 36414 57000
rect 37002 56200 37058 57000
rect 37646 56200 37702 57000
rect 38290 56200 38346 57000
rect 38934 56200 38990 57000
rect 39578 56200 39634 57000
rect 40222 56200 40278 57000
rect 42154 56200 42210 57000
rect 42798 56200 42854 57000
rect 43442 56200 43498 57000
rect 44086 56200 44142 57000
rect 44730 56200 44786 57000
rect 45374 56200 45430 57000
rect 46018 56200 46074 57000
rect 46662 56200 46718 57000
rect 47306 56200 47362 57000
rect 47950 56200 48006 57000
rect 48594 56200 48650 57000
rect 49238 56200 49294 57000
rect 30576 54262 30604 56200
rect 30564 54256 30616 54262
rect 30300 54194 30420 54210
rect 30564 54198 30616 54204
rect 30300 54188 30432 54194
rect 30300 54182 30380 54188
rect 30380 54130 30432 54136
rect 28908 54120 28960 54126
rect 28908 54062 28960 54068
rect 27804 53576 27856 53582
rect 27804 53518 27856 53524
rect 27950 53340 28258 53349
rect 27950 53338 27956 53340
rect 28012 53338 28036 53340
rect 28092 53338 28116 53340
rect 28172 53338 28196 53340
rect 28252 53338 28258 53340
rect 28012 53286 28014 53338
rect 28194 53286 28196 53338
rect 27950 53284 27956 53286
rect 28012 53284 28036 53286
rect 28092 53284 28116 53286
rect 28172 53284 28196 53286
rect 28252 53284 28258 53286
rect 27950 53275 28258 53284
rect 27950 52252 28258 52261
rect 27950 52250 27956 52252
rect 28012 52250 28036 52252
rect 28092 52250 28116 52252
rect 28172 52250 28196 52252
rect 28252 52250 28258 52252
rect 28012 52198 28014 52250
rect 28194 52198 28196 52250
rect 27950 52196 27956 52198
rect 28012 52196 28036 52198
rect 28092 52196 28116 52198
rect 28172 52196 28196 52198
rect 28252 52196 28258 52198
rect 27950 52187 28258 52196
rect 27950 51164 28258 51173
rect 27950 51162 27956 51164
rect 28012 51162 28036 51164
rect 28092 51162 28116 51164
rect 28172 51162 28196 51164
rect 28252 51162 28258 51164
rect 28012 51110 28014 51162
rect 28194 51110 28196 51162
rect 27950 51108 27956 51110
rect 28012 51108 28036 51110
rect 28092 51108 28116 51110
rect 28172 51108 28196 51110
rect 28252 51108 28258 51110
rect 27950 51099 28258 51108
rect 27620 50720 27672 50726
rect 27620 50662 27672 50668
rect 27160 49632 27212 49638
rect 27160 49574 27212 49580
rect 26148 47660 26200 47666
rect 26148 47602 26200 47608
rect 25780 43648 25832 43654
rect 25780 43590 25832 43596
rect 25872 20460 25924 20466
rect 25872 20402 25924 20408
rect 25412 17740 25464 17746
rect 25412 17682 25464 17688
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 24676 17196 24728 17202
rect 24676 17138 24728 17144
rect 24676 17060 24728 17066
rect 24676 17002 24728 17008
rect 24492 15156 24544 15162
rect 24492 15098 24544 15104
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 24688 14074 24716 17002
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 24676 14068 24728 14074
rect 24676 14010 24728 14016
rect 20720 14000 20772 14006
rect 20720 13942 20772 13948
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 20628 13728 20680 13734
rect 20628 13670 20680 13676
rect 20640 11354 20668 13670
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20640 7818 20668 11290
rect 20732 7954 20760 13942
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20628 7812 20680 7818
rect 20628 7754 20680 7760
rect 20916 6798 20944 14010
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 24688 13530 24716 14010
rect 24676 13524 24728 13530
rect 24676 13466 24728 13472
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 21364 12776 21416 12782
rect 21364 12718 21416 12724
rect 21376 12442 21404 12718
rect 22652 12708 22704 12714
rect 22652 12650 22704 12656
rect 21364 12436 21416 12442
rect 21364 12378 21416 12384
rect 21376 11218 21404 12378
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 21376 5710 21404 11154
rect 22664 6798 22692 12650
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23400 11150 23428 13262
rect 24124 12640 24176 12646
rect 24124 12582 24176 12588
rect 23388 11144 23440 11150
rect 23388 11086 23440 11092
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 22192 6724 22244 6730
rect 22192 6666 22244 6672
rect 23480 6724 23532 6730
rect 23480 6666 23532 6672
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 19524 2848 19576 2854
rect 19524 2790 19576 2796
rect 22100 2508 22152 2514
rect 22100 2450 22152 2456
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 22112 800 22140 2450
rect 22204 2446 22232 6666
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 23492 2446 23520 6666
rect 24136 6390 24164 12582
rect 24124 6384 24176 6390
rect 24124 6326 24176 6332
rect 24964 2582 24992 17614
rect 25136 17604 25188 17610
rect 25136 17546 25188 17552
rect 25148 16590 25176 17546
rect 25136 16584 25188 16590
rect 25136 16526 25188 16532
rect 25884 15502 25912 20402
rect 26160 17746 26188 47602
rect 27632 44946 27660 50662
rect 27950 50076 28258 50085
rect 27950 50074 27956 50076
rect 28012 50074 28036 50076
rect 28092 50074 28116 50076
rect 28172 50074 28196 50076
rect 28252 50074 28258 50076
rect 28012 50022 28014 50074
rect 28194 50022 28196 50074
rect 27950 50020 27956 50022
rect 28012 50020 28036 50022
rect 28092 50020 28116 50022
rect 28172 50020 28196 50022
rect 28252 50020 28258 50022
rect 27950 50011 28258 50020
rect 27950 48988 28258 48997
rect 27950 48986 27956 48988
rect 28012 48986 28036 48988
rect 28092 48986 28116 48988
rect 28172 48986 28196 48988
rect 28252 48986 28258 48988
rect 28012 48934 28014 48986
rect 28194 48934 28196 48986
rect 27950 48932 27956 48934
rect 28012 48932 28036 48934
rect 28092 48932 28116 48934
rect 28172 48932 28196 48934
rect 28252 48932 28258 48934
rect 27950 48923 28258 48932
rect 28920 48890 28948 54062
rect 29828 53984 29880 53990
rect 29828 53926 29880 53932
rect 30472 53984 30524 53990
rect 30472 53926 30524 53932
rect 31116 53984 31168 53990
rect 31116 53926 31168 53932
rect 28908 48884 28960 48890
rect 28908 48826 28960 48832
rect 27950 47900 28258 47909
rect 27950 47898 27956 47900
rect 28012 47898 28036 47900
rect 28092 47898 28116 47900
rect 28172 47898 28196 47900
rect 28252 47898 28258 47900
rect 28012 47846 28014 47898
rect 28194 47846 28196 47898
rect 27950 47844 27956 47846
rect 28012 47844 28036 47846
rect 28092 47844 28116 47846
rect 28172 47844 28196 47846
rect 28252 47844 28258 47846
rect 27950 47835 28258 47844
rect 27950 46812 28258 46821
rect 27950 46810 27956 46812
rect 28012 46810 28036 46812
rect 28092 46810 28116 46812
rect 28172 46810 28196 46812
rect 28252 46810 28258 46812
rect 28012 46758 28014 46810
rect 28194 46758 28196 46810
rect 27950 46756 27956 46758
rect 28012 46756 28036 46758
rect 28092 46756 28116 46758
rect 28172 46756 28196 46758
rect 28252 46756 28258 46758
rect 27950 46747 28258 46756
rect 27950 45724 28258 45733
rect 27950 45722 27956 45724
rect 28012 45722 28036 45724
rect 28092 45722 28116 45724
rect 28172 45722 28196 45724
rect 28252 45722 28258 45724
rect 28012 45670 28014 45722
rect 28194 45670 28196 45722
rect 27950 45668 27956 45670
rect 28012 45668 28036 45670
rect 28092 45668 28116 45670
rect 28172 45668 28196 45670
rect 28252 45668 28258 45670
rect 27950 45659 28258 45668
rect 27620 44940 27672 44946
rect 27620 44882 27672 44888
rect 26792 44736 26844 44742
rect 26792 44678 26844 44684
rect 27252 44736 27304 44742
rect 27252 44678 27304 44684
rect 26804 43790 26832 44678
rect 26792 43784 26844 43790
rect 26792 43726 26844 43732
rect 27264 41478 27292 44678
rect 27632 44334 27660 44882
rect 27950 44636 28258 44645
rect 27950 44634 27956 44636
rect 28012 44634 28036 44636
rect 28092 44634 28116 44636
rect 28172 44634 28196 44636
rect 28252 44634 28258 44636
rect 28012 44582 28014 44634
rect 28194 44582 28196 44634
rect 27950 44580 27956 44582
rect 28012 44580 28036 44582
rect 28092 44580 28116 44582
rect 28172 44580 28196 44582
rect 28252 44580 28258 44582
rect 27950 44571 28258 44580
rect 27620 44328 27672 44334
rect 27620 44270 27672 44276
rect 27632 43858 27660 44270
rect 27620 43852 27672 43858
rect 27620 43794 27672 43800
rect 27950 43548 28258 43557
rect 27950 43546 27956 43548
rect 28012 43546 28036 43548
rect 28092 43546 28116 43548
rect 28172 43546 28196 43548
rect 28252 43546 28258 43548
rect 28012 43494 28014 43546
rect 28194 43494 28196 43546
rect 27950 43492 27956 43494
rect 28012 43492 28036 43494
rect 28092 43492 28116 43494
rect 28172 43492 28196 43494
rect 28252 43492 28258 43494
rect 27950 43483 28258 43492
rect 29840 43353 29868 53926
rect 30380 53780 30432 53786
rect 30380 53722 30432 53728
rect 30392 47802 30420 53722
rect 30484 49230 30512 53926
rect 31128 49978 31156 53926
rect 31220 53582 31248 56200
rect 31864 53582 31892 56200
rect 32508 54262 32536 56200
rect 32772 54596 32824 54602
rect 32772 54538 32824 54544
rect 32784 54330 32812 54538
rect 32772 54324 32824 54330
rect 32772 54266 32824 54272
rect 33152 54262 33180 56200
rect 33796 54262 33824 56200
rect 34440 54262 34468 56200
rect 32496 54256 32548 54262
rect 32496 54198 32548 54204
rect 33140 54256 33192 54262
rect 33140 54198 33192 54204
rect 33784 54256 33836 54262
rect 33784 54198 33836 54204
rect 34428 54256 34480 54262
rect 34428 54198 34480 54204
rect 35084 54194 35112 56200
rect 35072 54188 35124 54194
rect 35728 54176 35756 56200
rect 35900 54188 35952 54194
rect 35728 54148 35900 54176
rect 35072 54130 35124 54136
rect 35900 54130 35952 54136
rect 35070 54088 35126 54097
rect 33784 54052 33836 54058
rect 35070 54023 35126 54032
rect 33784 53994 33836 54000
rect 32950 53884 33258 53893
rect 32950 53882 32956 53884
rect 33012 53882 33036 53884
rect 33092 53882 33116 53884
rect 33172 53882 33196 53884
rect 33252 53882 33258 53884
rect 33012 53830 33014 53882
rect 33194 53830 33196 53882
rect 32950 53828 32956 53830
rect 33012 53828 33036 53830
rect 33092 53828 33116 53830
rect 33172 53828 33196 53830
rect 33252 53828 33258 53830
rect 32950 53819 33258 53828
rect 33508 53712 33560 53718
rect 33508 53654 33560 53660
rect 31208 53576 31260 53582
rect 31208 53518 31260 53524
rect 31852 53576 31904 53582
rect 31852 53518 31904 53524
rect 32950 52796 33258 52805
rect 32950 52794 32956 52796
rect 33012 52794 33036 52796
rect 33092 52794 33116 52796
rect 33172 52794 33196 52796
rect 33252 52794 33258 52796
rect 33012 52742 33014 52794
rect 33194 52742 33196 52794
rect 32950 52740 32956 52742
rect 33012 52740 33036 52742
rect 33092 52740 33116 52742
rect 33172 52740 33196 52742
rect 33252 52740 33258 52742
rect 32950 52731 33258 52740
rect 32950 51708 33258 51717
rect 32950 51706 32956 51708
rect 33012 51706 33036 51708
rect 33092 51706 33116 51708
rect 33172 51706 33196 51708
rect 33252 51706 33258 51708
rect 33012 51654 33014 51706
rect 33194 51654 33196 51706
rect 32950 51652 32956 51654
rect 33012 51652 33036 51654
rect 33092 51652 33116 51654
rect 33172 51652 33196 51654
rect 33252 51652 33258 51654
rect 32950 51643 33258 51652
rect 33416 51060 33468 51066
rect 33416 51002 33468 51008
rect 32950 50620 33258 50629
rect 32950 50618 32956 50620
rect 33012 50618 33036 50620
rect 33092 50618 33116 50620
rect 33172 50618 33196 50620
rect 33252 50618 33258 50620
rect 33012 50566 33014 50618
rect 33194 50566 33196 50618
rect 32950 50564 32956 50566
rect 33012 50564 33036 50566
rect 33092 50564 33116 50566
rect 33172 50564 33196 50566
rect 33252 50564 33258 50566
rect 32950 50555 33258 50564
rect 31208 50244 31260 50250
rect 31208 50186 31260 50192
rect 31220 49978 31248 50186
rect 33428 49978 33456 51002
rect 31116 49972 31168 49978
rect 31116 49914 31168 49920
rect 31208 49972 31260 49978
rect 31208 49914 31260 49920
rect 33416 49972 33468 49978
rect 33416 49914 33468 49920
rect 32950 49532 33258 49541
rect 32950 49530 32956 49532
rect 33012 49530 33036 49532
rect 33092 49530 33116 49532
rect 33172 49530 33196 49532
rect 33252 49530 33258 49532
rect 33012 49478 33014 49530
rect 33194 49478 33196 49530
rect 32950 49476 32956 49478
rect 33012 49476 33036 49478
rect 33092 49476 33116 49478
rect 33172 49476 33196 49478
rect 33252 49476 33258 49478
rect 32950 49467 33258 49476
rect 30472 49224 30524 49230
rect 30472 49166 30524 49172
rect 30748 48748 30800 48754
rect 30748 48690 30800 48696
rect 30380 47796 30432 47802
rect 30380 47738 30432 47744
rect 29826 43344 29882 43353
rect 29826 43279 29882 43288
rect 27950 42460 28258 42469
rect 27950 42458 27956 42460
rect 28012 42458 28036 42460
rect 28092 42458 28116 42460
rect 28172 42458 28196 42460
rect 28252 42458 28258 42460
rect 28012 42406 28014 42458
rect 28194 42406 28196 42458
rect 27950 42404 27956 42406
rect 28012 42404 28036 42406
rect 28092 42404 28116 42406
rect 28172 42404 28196 42406
rect 28252 42404 28258 42406
rect 27950 42395 28258 42404
rect 27252 41472 27304 41478
rect 27252 41414 27304 41420
rect 27950 41372 28258 41381
rect 27950 41370 27956 41372
rect 28012 41370 28036 41372
rect 28092 41370 28116 41372
rect 28172 41370 28196 41372
rect 28252 41370 28258 41372
rect 28012 41318 28014 41370
rect 28194 41318 28196 41370
rect 27950 41316 27956 41318
rect 28012 41316 28036 41318
rect 28092 41316 28116 41318
rect 28172 41316 28196 41318
rect 28252 41316 28258 41318
rect 27950 41307 28258 41316
rect 27950 40284 28258 40293
rect 27950 40282 27956 40284
rect 28012 40282 28036 40284
rect 28092 40282 28116 40284
rect 28172 40282 28196 40284
rect 28252 40282 28258 40284
rect 28012 40230 28014 40282
rect 28194 40230 28196 40282
rect 27950 40228 27956 40230
rect 28012 40228 28036 40230
rect 28092 40228 28116 40230
rect 28172 40228 28196 40230
rect 28252 40228 28258 40230
rect 27950 40219 28258 40228
rect 27950 39196 28258 39205
rect 27950 39194 27956 39196
rect 28012 39194 28036 39196
rect 28092 39194 28116 39196
rect 28172 39194 28196 39196
rect 28252 39194 28258 39196
rect 28012 39142 28014 39194
rect 28194 39142 28196 39194
rect 27950 39140 27956 39142
rect 28012 39140 28036 39142
rect 28092 39140 28116 39142
rect 28172 39140 28196 39142
rect 28252 39140 28258 39142
rect 27950 39131 28258 39140
rect 27950 38108 28258 38117
rect 27950 38106 27956 38108
rect 28012 38106 28036 38108
rect 28092 38106 28116 38108
rect 28172 38106 28196 38108
rect 28252 38106 28258 38108
rect 28012 38054 28014 38106
rect 28194 38054 28196 38106
rect 27950 38052 27956 38054
rect 28012 38052 28036 38054
rect 28092 38052 28116 38054
rect 28172 38052 28196 38054
rect 28252 38052 28258 38054
rect 27950 38043 28258 38052
rect 27950 37020 28258 37029
rect 27950 37018 27956 37020
rect 28012 37018 28036 37020
rect 28092 37018 28116 37020
rect 28172 37018 28196 37020
rect 28252 37018 28258 37020
rect 28012 36966 28014 37018
rect 28194 36966 28196 37018
rect 27950 36964 27956 36966
rect 28012 36964 28036 36966
rect 28092 36964 28116 36966
rect 28172 36964 28196 36966
rect 28252 36964 28258 36966
rect 27950 36955 28258 36964
rect 27950 35932 28258 35941
rect 27950 35930 27956 35932
rect 28012 35930 28036 35932
rect 28092 35930 28116 35932
rect 28172 35930 28196 35932
rect 28252 35930 28258 35932
rect 28012 35878 28014 35930
rect 28194 35878 28196 35930
rect 27950 35876 27956 35878
rect 28012 35876 28036 35878
rect 28092 35876 28116 35878
rect 28172 35876 28196 35878
rect 28252 35876 28258 35878
rect 27950 35867 28258 35876
rect 27950 34844 28258 34853
rect 27950 34842 27956 34844
rect 28012 34842 28036 34844
rect 28092 34842 28116 34844
rect 28172 34842 28196 34844
rect 28252 34842 28258 34844
rect 28012 34790 28014 34842
rect 28194 34790 28196 34842
rect 27950 34788 27956 34790
rect 28012 34788 28036 34790
rect 28092 34788 28116 34790
rect 28172 34788 28196 34790
rect 28252 34788 28258 34790
rect 27950 34779 28258 34788
rect 27950 33756 28258 33765
rect 27950 33754 27956 33756
rect 28012 33754 28036 33756
rect 28092 33754 28116 33756
rect 28172 33754 28196 33756
rect 28252 33754 28258 33756
rect 28012 33702 28014 33754
rect 28194 33702 28196 33754
rect 27950 33700 27956 33702
rect 28012 33700 28036 33702
rect 28092 33700 28116 33702
rect 28172 33700 28196 33702
rect 28252 33700 28258 33702
rect 27950 33691 28258 33700
rect 27950 32668 28258 32677
rect 27950 32666 27956 32668
rect 28012 32666 28036 32668
rect 28092 32666 28116 32668
rect 28172 32666 28196 32668
rect 28252 32666 28258 32668
rect 28012 32614 28014 32666
rect 28194 32614 28196 32666
rect 27950 32612 27956 32614
rect 28012 32612 28036 32614
rect 28092 32612 28116 32614
rect 28172 32612 28196 32614
rect 28252 32612 28258 32614
rect 27950 32603 28258 32612
rect 27950 31580 28258 31589
rect 27950 31578 27956 31580
rect 28012 31578 28036 31580
rect 28092 31578 28116 31580
rect 28172 31578 28196 31580
rect 28252 31578 28258 31580
rect 28012 31526 28014 31578
rect 28194 31526 28196 31578
rect 27950 31524 27956 31526
rect 28012 31524 28036 31526
rect 28092 31524 28116 31526
rect 28172 31524 28196 31526
rect 28252 31524 28258 31526
rect 27950 31515 28258 31524
rect 27950 30492 28258 30501
rect 27950 30490 27956 30492
rect 28012 30490 28036 30492
rect 28092 30490 28116 30492
rect 28172 30490 28196 30492
rect 28252 30490 28258 30492
rect 28012 30438 28014 30490
rect 28194 30438 28196 30490
rect 27950 30436 27956 30438
rect 28012 30436 28036 30438
rect 28092 30436 28116 30438
rect 28172 30436 28196 30438
rect 28252 30436 28258 30438
rect 27950 30427 28258 30436
rect 27950 29404 28258 29413
rect 27950 29402 27956 29404
rect 28012 29402 28036 29404
rect 28092 29402 28116 29404
rect 28172 29402 28196 29404
rect 28252 29402 28258 29404
rect 28012 29350 28014 29402
rect 28194 29350 28196 29402
rect 27950 29348 27956 29350
rect 28012 29348 28036 29350
rect 28092 29348 28116 29350
rect 28172 29348 28196 29350
rect 28252 29348 28258 29350
rect 27950 29339 28258 29348
rect 27950 28316 28258 28325
rect 27950 28314 27956 28316
rect 28012 28314 28036 28316
rect 28092 28314 28116 28316
rect 28172 28314 28196 28316
rect 28252 28314 28258 28316
rect 28012 28262 28014 28314
rect 28194 28262 28196 28314
rect 27950 28260 27956 28262
rect 28012 28260 28036 28262
rect 28092 28260 28116 28262
rect 28172 28260 28196 28262
rect 28252 28260 28258 28262
rect 27950 28251 28258 28260
rect 27950 27228 28258 27237
rect 27950 27226 27956 27228
rect 28012 27226 28036 27228
rect 28092 27226 28116 27228
rect 28172 27226 28196 27228
rect 28252 27226 28258 27228
rect 28012 27174 28014 27226
rect 28194 27174 28196 27226
rect 27950 27172 27956 27174
rect 28012 27172 28036 27174
rect 28092 27172 28116 27174
rect 28172 27172 28196 27174
rect 28252 27172 28258 27174
rect 27950 27163 28258 27172
rect 27950 26140 28258 26149
rect 27950 26138 27956 26140
rect 28012 26138 28036 26140
rect 28092 26138 28116 26140
rect 28172 26138 28196 26140
rect 28252 26138 28258 26140
rect 28012 26086 28014 26138
rect 28194 26086 28196 26138
rect 27950 26084 27956 26086
rect 28012 26084 28036 26086
rect 28092 26084 28116 26086
rect 28172 26084 28196 26086
rect 28252 26084 28258 26086
rect 27950 26075 28258 26084
rect 27950 25052 28258 25061
rect 27950 25050 27956 25052
rect 28012 25050 28036 25052
rect 28092 25050 28116 25052
rect 28172 25050 28196 25052
rect 28252 25050 28258 25052
rect 28012 24998 28014 25050
rect 28194 24998 28196 25050
rect 27950 24996 27956 24998
rect 28012 24996 28036 24998
rect 28092 24996 28116 24998
rect 28172 24996 28196 24998
rect 28252 24996 28258 24998
rect 27950 24987 28258 24996
rect 26424 24676 26476 24682
rect 26424 24618 26476 24624
rect 26148 17740 26200 17746
rect 26148 17682 26200 17688
rect 26436 17338 26464 24618
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 27252 17672 27304 17678
rect 27252 17614 27304 17620
rect 26424 17332 26476 17338
rect 26424 17274 26476 17280
rect 26436 15706 26464 17274
rect 26424 15700 26476 15706
rect 26424 15642 26476 15648
rect 25872 15496 25924 15502
rect 25872 15438 25924 15444
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 25056 13190 25084 14350
rect 25884 13326 25912 15438
rect 25964 15360 26016 15366
rect 25964 15302 26016 15308
rect 25976 15026 26004 15302
rect 25964 15020 26016 15026
rect 25964 14962 26016 14968
rect 26700 13932 26752 13938
rect 26700 13874 26752 13880
rect 25872 13320 25924 13326
rect 25872 13262 25924 13268
rect 25044 13184 25096 13190
rect 25044 13126 25096 13132
rect 26712 12442 26740 13874
rect 26700 12436 26752 12442
rect 26700 12378 26752 12384
rect 24952 2576 25004 2582
rect 24952 2518 25004 2524
rect 25412 2508 25464 2514
rect 25412 2450 25464 2456
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 25424 800 25452 2450
rect 27264 2378 27292 17614
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 30760 17270 30788 48690
rect 32950 48444 33258 48453
rect 32950 48442 32956 48444
rect 33012 48442 33036 48444
rect 33092 48442 33116 48444
rect 33172 48442 33196 48444
rect 33252 48442 33258 48444
rect 33012 48390 33014 48442
rect 33194 48390 33196 48442
rect 32950 48388 32956 48390
rect 33012 48388 33036 48390
rect 33092 48388 33116 48390
rect 33172 48388 33196 48390
rect 33252 48388 33258 48390
rect 32950 48379 33258 48388
rect 32864 48136 32916 48142
rect 32864 48078 32916 48084
rect 30748 17264 30800 17270
rect 30748 17206 30800 17212
rect 28908 17128 28960 17134
rect 28908 17070 28960 17076
rect 29092 17128 29144 17134
rect 29092 17070 29144 17076
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 28816 6180 28868 6186
rect 28816 6122 28868 6128
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 28828 3058 28856 6122
rect 28816 3052 28868 3058
rect 28816 2994 28868 3000
rect 28724 2984 28776 2990
rect 28724 2926 28776 2932
rect 27252 2372 27304 2378
rect 27252 2314 27304 2320
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 28736 800 28764 2926
rect 28920 2582 28948 17070
rect 29104 14278 29132 17070
rect 31024 16652 31076 16658
rect 31024 16594 31076 16600
rect 29092 14272 29144 14278
rect 29092 14214 29144 14220
rect 31036 2650 31064 16594
rect 32876 16590 32904 48078
rect 32950 47356 33258 47365
rect 32950 47354 32956 47356
rect 33012 47354 33036 47356
rect 33092 47354 33116 47356
rect 33172 47354 33196 47356
rect 33252 47354 33258 47356
rect 33012 47302 33014 47354
rect 33194 47302 33196 47354
rect 32950 47300 32956 47302
rect 33012 47300 33036 47302
rect 33092 47300 33116 47302
rect 33172 47300 33196 47302
rect 33252 47300 33258 47302
rect 32950 47291 33258 47300
rect 33520 46578 33548 53654
rect 33692 49972 33744 49978
rect 33692 49914 33744 49920
rect 33508 46572 33560 46578
rect 33508 46514 33560 46520
rect 32950 46268 33258 46277
rect 32950 46266 32956 46268
rect 33012 46266 33036 46268
rect 33092 46266 33116 46268
rect 33172 46266 33196 46268
rect 33252 46266 33258 46268
rect 33012 46214 33014 46266
rect 33194 46214 33196 46266
rect 32950 46212 32956 46214
rect 33012 46212 33036 46214
rect 33092 46212 33116 46214
rect 33172 46212 33196 46214
rect 33252 46212 33258 46214
rect 32950 46203 33258 46212
rect 32950 45180 33258 45189
rect 32950 45178 32956 45180
rect 33012 45178 33036 45180
rect 33092 45178 33116 45180
rect 33172 45178 33196 45180
rect 33252 45178 33258 45180
rect 33012 45126 33014 45178
rect 33194 45126 33196 45178
rect 32950 45124 32956 45126
rect 33012 45124 33036 45126
rect 33092 45124 33116 45126
rect 33172 45124 33196 45126
rect 33252 45124 33258 45126
rect 32950 45115 33258 45124
rect 32950 44092 33258 44101
rect 32950 44090 32956 44092
rect 33012 44090 33036 44092
rect 33092 44090 33116 44092
rect 33172 44090 33196 44092
rect 33252 44090 33258 44092
rect 33012 44038 33014 44090
rect 33194 44038 33196 44090
rect 32950 44036 32956 44038
rect 33012 44036 33036 44038
rect 33092 44036 33116 44038
rect 33172 44036 33196 44038
rect 33252 44036 33258 44038
rect 32950 44027 33258 44036
rect 32950 43004 33258 43013
rect 32950 43002 32956 43004
rect 33012 43002 33036 43004
rect 33092 43002 33116 43004
rect 33172 43002 33196 43004
rect 33252 43002 33258 43004
rect 33012 42950 33014 43002
rect 33194 42950 33196 43002
rect 32950 42948 32956 42950
rect 33012 42948 33036 42950
rect 33092 42948 33116 42950
rect 33172 42948 33196 42950
rect 33252 42948 33258 42950
rect 32950 42939 33258 42948
rect 32950 41916 33258 41925
rect 32950 41914 32956 41916
rect 33012 41914 33036 41916
rect 33092 41914 33116 41916
rect 33172 41914 33196 41916
rect 33252 41914 33258 41916
rect 33012 41862 33014 41914
rect 33194 41862 33196 41914
rect 32950 41860 32956 41862
rect 33012 41860 33036 41862
rect 33092 41860 33116 41862
rect 33172 41860 33196 41862
rect 33252 41860 33258 41862
rect 32950 41851 33258 41860
rect 32950 40828 33258 40837
rect 32950 40826 32956 40828
rect 33012 40826 33036 40828
rect 33092 40826 33116 40828
rect 33172 40826 33196 40828
rect 33252 40826 33258 40828
rect 33012 40774 33014 40826
rect 33194 40774 33196 40826
rect 32950 40772 32956 40774
rect 33012 40772 33036 40774
rect 33092 40772 33116 40774
rect 33172 40772 33196 40774
rect 33252 40772 33258 40774
rect 32950 40763 33258 40772
rect 32950 39740 33258 39749
rect 32950 39738 32956 39740
rect 33012 39738 33036 39740
rect 33092 39738 33116 39740
rect 33172 39738 33196 39740
rect 33252 39738 33258 39740
rect 33012 39686 33014 39738
rect 33194 39686 33196 39738
rect 32950 39684 32956 39686
rect 33012 39684 33036 39686
rect 33092 39684 33116 39686
rect 33172 39684 33196 39686
rect 33252 39684 33258 39686
rect 32950 39675 33258 39684
rect 32950 38652 33258 38661
rect 32950 38650 32956 38652
rect 33012 38650 33036 38652
rect 33092 38650 33116 38652
rect 33172 38650 33196 38652
rect 33252 38650 33258 38652
rect 33012 38598 33014 38650
rect 33194 38598 33196 38650
rect 32950 38596 32956 38598
rect 33012 38596 33036 38598
rect 33092 38596 33116 38598
rect 33172 38596 33196 38598
rect 33252 38596 33258 38598
rect 32950 38587 33258 38596
rect 32950 37564 33258 37573
rect 32950 37562 32956 37564
rect 33012 37562 33036 37564
rect 33092 37562 33116 37564
rect 33172 37562 33196 37564
rect 33252 37562 33258 37564
rect 33012 37510 33014 37562
rect 33194 37510 33196 37562
rect 32950 37508 32956 37510
rect 33012 37508 33036 37510
rect 33092 37508 33116 37510
rect 33172 37508 33196 37510
rect 33252 37508 33258 37510
rect 32950 37499 33258 37508
rect 32950 36476 33258 36485
rect 32950 36474 32956 36476
rect 33012 36474 33036 36476
rect 33092 36474 33116 36476
rect 33172 36474 33196 36476
rect 33252 36474 33258 36476
rect 33012 36422 33014 36474
rect 33194 36422 33196 36474
rect 32950 36420 32956 36422
rect 33012 36420 33036 36422
rect 33092 36420 33116 36422
rect 33172 36420 33196 36422
rect 33252 36420 33258 36422
rect 32950 36411 33258 36420
rect 32950 35388 33258 35397
rect 32950 35386 32956 35388
rect 33012 35386 33036 35388
rect 33092 35386 33116 35388
rect 33172 35386 33196 35388
rect 33252 35386 33258 35388
rect 33012 35334 33014 35386
rect 33194 35334 33196 35386
rect 32950 35332 32956 35334
rect 33012 35332 33036 35334
rect 33092 35332 33116 35334
rect 33172 35332 33196 35334
rect 33252 35332 33258 35334
rect 32950 35323 33258 35332
rect 32950 34300 33258 34309
rect 32950 34298 32956 34300
rect 33012 34298 33036 34300
rect 33092 34298 33116 34300
rect 33172 34298 33196 34300
rect 33252 34298 33258 34300
rect 33012 34246 33014 34298
rect 33194 34246 33196 34298
rect 32950 34244 32956 34246
rect 33012 34244 33036 34246
rect 33092 34244 33116 34246
rect 33172 34244 33196 34246
rect 33252 34244 33258 34246
rect 32950 34235 33258 34244
rect 32950 33212 33258 33221
rect 32950 33210 32956 33212
rect 33012 33210 33036 33212
rect 33092 33210 33116 33212
rect 33172 33210 33196 33212
rect 33252 33210 33258 33212
rect 33012 33158 33014 33210
rect 33194 33158 33196 33210
rect 32950 33156 32956 33158
rect 33012 33156 33036 33158
rect 33092 33156 33116 33158
rect 33172 33156 33196 33158
rect 33252 33156 33258 33158
rect 32950 33147 33258 33156
rect 32950 32124 33258 32133
rect 32950 32122 32956 32124
rect 33012 32122 33036 32124
rect 33092 32122 33116 32124
rect 33172 32122 33196 32124
rect 33252 32122 33258 32124
rect 33012 32070 33014 32122
rect 33194 32070 33196 32122
rect 32950 32068 32956 32070
rect 33012 32068 33036 32070
rect 33092 32068 33116 32070
rect 33172 32068 33196 32070
rect 33252 32068 33258 32070
rect 32950 32059 33258 32068
rect 32950 31036 33258 31045
rect 32950 31034 32956 31036
rect 33012 31034 33036 31036
rect 33092 31034 33116 31036
rect 33172 31034 33196 31036
rect 33252 31034 33258 31036
rect 33012 30982 33014 31034
rect 33194 30982 33196 31034
rect 32950 30980 32956 30982
rect 33012 30980 33036 30982
rect 33092 30980 33116 30982
rect 33172 30980 33196 30982
rect 33252 30980 33258 30982
rect 32950 30971 33258 30980
rect 32950 29948 33258 29957
rect 32950 29946 32956 29948
rect 33012 29946 33036 29948
rect 33092 29946 33116 29948
rect 33172 29946 33196 29948
rect 33252 29946 33258 29948
rect 33012 29894 33014 29946
rect 33194 29894 33196 29946
rect 32950 29892 32956 29894
rect 33012 29892 33036 29894
rect 33092 29892 33116 29894
rect 33172 29892 33196 29894
rect 33252 29892 33258 29894
rect 32950 29883 33258 29892
rect 32950 28860 33258 28869
rect 32950 28858 32956 28860
rect 33012 28858 33036 28860
rect 33092 28858 33116 28860
rect 33172 28858 33196 28860
rect 33252 28858 33258 28860
rect 33012 28806 33014 28858
rect 33194 28806 33196 28858
rect 32950 28804 32956 28806
rect 33012 28804 33036 28806
rect 33092 28804 33116 28806
rect 33172 28804 33196 28806
rect 33252 28804 33258 28806
rect 32950 28795 33258 28804
rect 32950 27772 33258 27781
rect 32950 27770 32956 27772
rect 33012 27770 33036 27772
rect 33092 27770 33116 27772
rect 33172 27770 33196 27772
rect 33252 27770 33258 27772
rect 33012 27718 33014 27770
rect 33194 27718 33196 27770
rect 32950 27716 32956 27718
rect 33012 27716 33036 27718
rect 33092 27716 33116 27718
rect 33172 27716 33196 27718
rect 33252 27716 33258 27718
rect 32950 27707 33258 27716
rect 32950 26684 33258 26693
rect 32950 26682 32956 26684
rect 33012 26682 33036 26684
rect 33092 26682 33116 26684
rect 33172 26682 33196 26684
rect 33252 26682 33258 26684
rect 33012 26630 33014 26682
rect 33194 26630 33196 26682
rect 32950 26628 32956 26630
rect 33012 26628 33036 26630
rect 33092 26628 33116 26630
rect 33172 26628 33196 26630
rect 33252 26628 33258 26630
rect 32950 26619 33258 26628
rect 32950 25596 33258 25605
rect 32950 25594 32956 25596
rect 33012 25594 33036 25596
rect 33092 25594 33116 25596
rect 33172 25594 33196 25596
rect 33252 25594 33258 25596
rect 33012 25542 33014 25594
rect 33194 25542 33196 25594
rect 32950 25540 32956 25542
rect 33012 25540 33036 25542
rect 33092 25540 33116 25542
rect 33172 25540 33196 25542
rect 33252 25540 33258 25542
rect 32950 25531 33258 25540
rect 33704 24818 33732 49914
rect 33796 49094 33824 53994
rect 35084 53990 35112 54023
rect 34244 53984 34296 53990
rect 34244 53926 34296 53932
rect 35072 53984 35124 53990
rect 35072 53926 35124 53932
rect 33784 49088 33836 49094
rect 33784 49030 33836 49036
rect 34256 41177 34284 53926
rect 36372 53582 36400 56200
rect 37016 53582 37044 56200
rect 37660 54262 37688 56200
rect 37950 54428 38258 54437
rect 37950 54426 37956 54428
rect 38012 54426 38036 54428
rect 38092 54426 38116 54428
rect 38172 54426 38196 54428
rect 38252 54426 38258 54428
rect 38012 54374 38014 54426
rect 38194 54374 38196 54426
rect 37950 54372 37956 54374
rect 38012 54372 38036 54374
rect 38092 54372 38116 54374
rect 38172 54372 38196 54374
rect 38252 54372 38258 54374
rect 37950 54363 38258 54372
rect 37648 54256 37700 54262
rect 37648 54198 37700 54204
rect 37832 53984 37884 53990
rect 37832 53926 37884 53932
rect 36360 53576 36412 53582
rect 36360 53518 36412 53524
rect 37004 53576 37056 53582
rect 37004 53518 37056 53524
rect 37556 50856 37608 50862
rect 37556 50798 37608 50804
rect 37568 49774 37596 50798
rect 37556 49768 37608 49774
rect 37556 49710 37608 49716
rect 34242 41168 34298 41177
rect 34242 41103 34298 41112
rect 37844 39642 37872 53926
rect 38304 53582 38332 56200
rect 38948 54262 38976 56200
rect 38936 54256 38988 54262
rect 38936 54198 38988 54204
rect 39592 54194 39620 56200
rect 39580 54188 39632 54194
rect 39580 54130 39632 54136
rect 38844 54120 38896 54126
rect 38844 54062 38896 54068
rect 38292 53576 38344 53582
rect 38292 53518 38344 53524
rect 38660 53508 38712 53514
rect 38660 53450 38712 53456
rect 37950 53340 38258 53349
rect 37950 53338 37956 53340
rect 38012 53338 38036 53340
rect 38092 53338 38116 53340
rect 38172 53338 38196 53340
rect 38252 53338 38258 53340
rect 38012 53286 38014 53338
rect 38194 53286 38196 53338
rect 37950 53284 37956 53286
rect 38012 53284 38036 53286
rect 38092 53284 38116 53286
rect 38172 53284 38196 53286
rect 38252 53284 38258 53286
rect 37950 53275 38258 53284
rect 37950 52252 38258 52261
rect 37950 52250 37956 52252
rect 38012 52250 38036 52252
rect 38092 52250 38116 52252
rect 38172 52250 38196 52252
rect 38252 52250 38258 52252
rect 38012 52198 38014 52250
rect 38194 52198 38196 52250
rect 37950 52196 37956 52198
rect 38012 52196 38036 52198
rect 38092 52196 38116 52198
rect 38172 52196 38196 52198
rect 38252 52196 38258 52198
rect 37950 52187 38258 52196
rect 37950 51164 38258 51173
rect 37950 51162 37956 51164
rect 38012 51162 38036 51164
rect 38092 51162 38116 51164
rect 38172 51162 38196 51164
rect 38252 51162 38258 51164
rect 38012 51110 38014 51162
rect 38194 51110 38196 51162
rect 37950 51108 37956 51110
rect 38012 51108 38036 51110
rect 38092 51108 38116 51110
rect 38172 51108 38196 51110
rect 38252 51108 38258 51110
rect 37950 51099 38258 51108
rect 37950 50076 38258 50085
rect 37950 50074 37956 50076
rect 38012 50074 38036 50076
rect 38092 50074 38116 50076
rect 38172 50074 38196 50076
rect 38252 50074 38258 50076
rect 38012 50022 38014 50074
rect 38194 50022 38196 50074
rect 37950 50020 37956 50022
rect 38012 50020 38036 50022
rect 38092 50020 38116 50022
rect 38172 50020 38196 50022
rect 38252 50020 38258 50022
rect 37950 50011 38258 50020
rect 37950 48988 38258 48997
rect 37950 48986 37956 48988
rect 38012 48986 38036 48988
rect 38092 48986 38116 48988
rect 38172 48986 38196 48988
rect 38252 48986 38258 48988
rect 38012 48934 38014 48986
rect 38194 48934 38196 48986
rect 37950 48932 37956 48934
rect 38012 48932 38036 48934
rect 38092 48932 38116 48934
rect 38172 48932 38196 48934
rect 38252 48932 38258 48934
rect 37950 48923 38258 48932
rect 37950 47900 38258 47909
rect 37950 47898 37956 47900
rect 38012 47898 38036 47900
rect 38092 47898 38116 47900
rect 38172 47898 38196 47900
rect 38252 47898 38258 47900
rect 38012 47846 38014 47898
rect 38194 47846 38196 47898
rect 37950 47844 37956 47846
rect 38012 47844 38036 47846
rect 38092 47844 38116 47846
rect 38172 47844 38196 47846
rect 38252 47844 38258 47846
rect 37950 47835 38258 47844
rect 37950 46812 38258 46821
rect 37950 46810 37956 46812
rect 38012 46810 38036 46812
rect 38092 46810 38116 46812
rect 38172 46810 38196 46812
rect 38252 46810 38258 46812
rect 38012 46758 38014 46810
rect 38194 46758 38196 46810
rect 37950 46756 37956 46758
rect 38012 46756 38036 46758
rect 38092 46756 38116 46758
rect 38172 46756 38196 46758
rect 38252 46756 38258 46758
rect 37950 46747 38258 46756
rect 37950 45724 38258 45733
rect 37950 45722 37956 45724
rect 38012 45722 38036 45724
rect 38092 45722 38116 45724
rect 38172 45722 38196 45724
rect 38252 45722 38258 45724
rect 38012 45670 38014 45722
rect 38194 45670 38196 45722
rect 37950 45668 37956 45670
rect 38012 45668 38036 45670
rect 38092 45668 38116 45670
rect 38172 45668 38196 45670
rect 38252 45668 38258 45670
rect 37950 45659 38258 45668
rect 37950 44636 38258 44645
rect 37950 44634 37956 44636
rect 38012 44634 38036 44636
rect 38092 44634 38116 44636
rect 38172 44634 38196 44636
rect 38252 44634 38258 44636
rect 38012 44582 38014 44634
rect 38194 44582 38196 44634
rect 37950 44580 37956 44582
rect 38012 44580 38036 44582
rect 38092 44580 38116 44582
rect 38172 44580 38196 44582
rect 38252 44580 38258 44582
rect 37950 44571 38258 44580
rect 37950 43548 38258 43557
rect 37950 43546 37956 43548
rect 38012 43546 38036 43548
rect 38092 43546 38116 43548
rect 38172 43546 38196 43548
rect 38252 43546 38258 43548
rect 38012 43494 38014 43546
rect 38194 43494 38196 43546
rect 37950 43492 37956 43494
rect 38012 43492 38036 43494
rect 38092 43492 38116 43494
rect 38172 43492 38196 43494
rect 38252 43492 38258 43494
rect 37950 43483 38258 43492
rect 37950 42460 38258 42469
rect 37950 42458 37956 42460
rect 38012 42458 38036 42460
rect 38092 42458 38116 42460
rect 38172 42458 38196 42460
rect 38252 42458 38258 42460
rect 38012 42406 38014 42458
rect 38194 42406 38196 42458
rect 37950 42404 37956 42406
rect 38012 42404 38036 42406
rect 38092 42404 38116 42406
rect 38172 42404 38196 42406
rect 38252 42404 38258 42406
rect 37950 42395 38258 42404
rect 37950 41372 38258 41381
rect 37950 41370 37956 41372
rect 38012 41370 38036 41372
rect 38092 41370 38116 41372
rect 38172 41370 38196 41372
rect 38252 41370 38258 41372
rect 38012 41318 38014 41370
rect 38194 41318 38196 41370
rect 37950 41316 37956 41318
rect 38012 41316 38036 41318
rect 38092 41316 38116 41318
rect 38172 41316 38196 41318
rect 38252 41316 38258 41318
rect 37950 41307 38258 41316
rect 37950 40284 38258 40293
rect 37950 40282 37956 40284
rect 38012 40282 38036 40284
rect 38092 40282 38116 40284
rect 38172 40282 38196 40284
rect 38252 40282 38258 40284
rect 38012 40230 38014 40282
rect 38194 40230 38196 40282
rect 37950 40228 37956 40230
rect 38012 40228 38036 40230
rect 38092 40228 38116 40230
rect 38172 40228 38196 40230
rect 38252 40228 38258 40230
rect 37950 40219 38258 40228
rect 38672 39846 38700 53450
rect 38856 45554 38884 54062
rect 40236 53582 40264 56200
rect 42168 54262 42196 56200
rect 42156 54256 42208 54262
rect 42156 54198 42208 54204
rect 40316 54120 40368 54126
rect 40316 54062 40368 54068
rect 40224 53576 40276 53582
rect 40224 53518 40276 53524
rect 40040 53440 40092 53446
rect 40040 53382 40092 53388
rect 40052 48006 40080 53382
rect 40040 48000 40092 48006
rect 40040 47942 40092 47948
rect 40328 45554 40356 54062
rect 43904 53984 43956 53990
rect 43904 53926 43956 53932
rect 42950 53884 43258 53893
rect 42950 53882 42956 53884
rect 43012 53882 43036 53884
rect 43092 53882 43116 53884
rect 43172 53882 43196 53884
rect 43252 53882 43258 53884
rect 43012 53830 43014 53882
rect 43194 53830 43196 53882
rect 42950 53828 42956 53830
rect 43012 53828 43036 53830
rect 43092 53828 43116 53830
rect 43172 53828 43196 53830
rect 43252 53828 43258 53830
rect 42950 53819 43258 53828
rect 42950 52796 43258 52805
rect 42950 52794 42956 52796
rect 43012 52794 43036 52796
rect 43092 52794 43116 52796
rect 43172 52794 43196 52796
rect 43252 52794 43258 52796
rect 43012 52742 43014 52794
rect 43194 52742 43196 52794
rect 42950 52740 42956 52742
rect 43012 52740 43036 52742
rect 43092 52740 43116 52742
rect 43172 52740 43196 52742
rect 43252 52740 43258 52742
rect 42950 52731 43258 52740
rect 42950 51708 43258 51717
rect 42950 51706 42956 51708
rect 43012 51706 43036 51708
rect 43092 51706 43116 51708
rect 43172 51706 43196 51708
rect 43252 51706 43258 51708
rect 43012 51654 43014 51706
rect 43194 51654 43196 51706
rect 42950 51652 42956 51654
rect 43012 51652 43036 51654
rect 43092 51652 43116 51654
rect 43172 51652 43196 51654
rect 43252 51652 43258 51654
rect 42950 51643 43258 51652
rect 43916 50998 43944 53926
rect 44100 53582 44128 56200
rect 44744 54194 44772 56200
rect 45388 54618 45416 56200
rect 45388 54590 45600 54618
rect 45572 54194 45600 54590
rect 46032 54194 46060 56200
rect 44732 54188 44784 54194
rect 44732 54130 44784 54136
rect 45560 54188 45612 54194
rect 45560 54130 45612 54136
rect 46020 54188 46072 54194
rect 46020 54130 46072 54136
rect 45284 53984 45336 53990
rect 45284 53926 45336 53932
rect 46112 53984 46164 53990
rect 46112 53926 46164 53932
rect 44088 53576 44140 53582
rect 44088 53518 44140 53524
rect 44364 53440 44416 53446
rect 44364 53382 44416 53388
rect 43904 50992 43956 50998
rect 43904 50934 43956 50940
rect 42950 50620 43258 50629
rect 42950 50618 42956 50620
rect 43012 50618 43036 50620
rect 43092 50618 43116 50620
rect 43172 50618 43196 50620
rect 43252 50618 43258 50620
rect 43012 50566 43014 50618
rect 43194 50566 43196 50618
rect 42950 50564 42956 50566
rect 43012 50564 43036 50566
rect 43092 50564 43116 50566
rect 43172 50564 43196 50566
rect 43252 50564 43258 50566
rect 42950 50555 43258 50564
rect 42950 49532 43258 49541
rect 42950 49530 42956 49532
rect 43012 49530 43036 49532
rect 43092 49530 43116 49532
rect 43172 49530 43196 49532
rect 43252 49530 43258 49532
rect 43012 49478 43014 49530
rect 43194 49478 43196 49530
rect 42950 49476 42956 49478
rect 43012 49476 43036 49478
rect 43092 49476 43116 49478
rect 43172 49476 43196 49478
rect 43252 49476 43258 49478
rect 42950 49467 43258 49476
rect 42950 48444 43258 48453
rect 42950 48442 42956 48444
rect 43012 48442 43036 48444
rect 43092 48442 43116 48444
rect 43172 48442 43196 48444
rect 43252 48442 43258 48444
rect 43012 48390 43014 48442
rect 43194 48390 43196 48442
rect 42950 48388 42956 48390
rect 43012 48388 43036 48390
rect 43092 48388 43116 48390
rect 43172 48388 43196 48390
rect 43252 48388 43258 48390
rect 42950 48379 43258 48388
rect 42950 47356 43258 47365
rect 42950 47354 42956 47356
rect 43012 47354 43036 47356
rect 43092 47354 43116 47356
rect 43172 47354 43196 47356
rect 43252 47354 43258 47356
rect 43012 47302 43014 47354
rect 43194 47302 43196 47354
rect 42950 47300 42956 47302
rect 43012 47300 43036 47302
rect 43092 47300 43116 47302
rect 43172 47300 43196 47302
rect 43252 47300 43258 47302
rect 42950 47291 43258 47300
rect 42950 46268 43258 46277
rect 42950 46266 42956 46268
rect 43012 46266 43036 46268
rect 43092 46266 43116 46268
rect 43172 46266 43196 46268
rect 43252 46266 43258 46268
rect 43012 46214 43014 46266
rect 43194 46214 43196 46266
rect 42950 46212 42956 46214
rect 43012 46212 43036 46214
rect 43092 46212 43116 46214
rect 43172 46212 43196 46214
rect 43252 46212 43258 46214
rect 42950 46203 43258 46212
rect 38856 45526 38976 45554
rect 38948 42673 38976 45526
rect 40236 45526 40356 45554
rect 40236 42809 40264 45526
rect 42950 45180 43258 45189
rect 42950 45178 42956 45180
rect 43012 45178 43036 45180
rect 43092 45178 43116 45180
rect 43172 45178 43196 45180
rect 43252 45178 43258 45180
rect 43012 45126 43014 45178
rect 43194 45126 43196 45178
rect 42950 45124 42956 45126
rect 43012 45124 43036 45126
rect 43092 45124 43116 45126
rect 43172 45124 43196 45126
rect 43252 45124 43258 45126
rect 42950 45115 43258 45124
rect 44376 44810 44404 53382
rect 44364 44804 44416 44810
rect 44364 44746 44416 44752
rect 42950 44092 43258 44101
rect 42950 44090 42956 44092
rect 43012 44090 43036 44092
rect 43092 44090 43116 44092
rect 43172 44090 43196 44092
rect 43252 44090 43258 44092
rect 43012 44038 43014 44090
rect 43194 44038 43196 44090
rect 42950 44036 42956 44038
rect 43012 44036 43036 44038
rect 43092 44036 43116 44038
rect 43172 44036 43196 44038
rect 43252 44036 43258 44038
rect 42950 44027 43258 44036
rect 42950 43004 43258 43013
rect 42950 43002 42956 43004
rect 43012 43002 43036 43004
rect 43092 43002 43116 43004
rect 43172 43002 43196 43004
rect 43252 43002 43258 43004
rect 43012 42950 43014 43002
rect 43194 42950 43196 43002
rect 42950 42948 42956 42950
rect 43012 42948 43036 42950
rect 43092 42948 43116 42950
rect 43172 42948 43196 42950
rect 43252 42948 43258 42950
rect 42950 42939 43258 42948
rect 40222 42800 40278 42809
rect 40222 42735 40278 42744
rect 38934 42664 38990 42673
rect 38934 42599 38990 42608
rect 42950 41916 43258 41925
rect 42950 41914 42956 41916
rect 43012 41914 43036 41916
rect 43092 41914 43116 41916
rect 43172 41914 43196 41916
rect 43252 41914 43258 41916
rect 43012 41862 43014 41914
rect 43194 41862 43196 41914
rect 42950 41860 42956 41862
rect 43012 41860 43036 41862
rect 43092 41860 43116 41862
rect 43172 41860 43196 41862
rect 43252 41860 43258 41862
rect 42950 41851 43258 41860
rect 42950 40828 43258 40837
rect 42950 40826 42956 40828
rect 43012 40826 43036 40828
rect 43092 40826 43116 40828
rect 43172 40826 43196 40828
rect 43252 40826 43258 40828
rect 43012 40774 43014 40826
rect 43194 40774 43196 40826
rect 42950 40772 42956 40774
rect 43012 40772 43036 40774
rect 43092 40772 43116 40774
rect 43172 40772 43196 40774
rect 43252 40772 43258 40774
rect 42950 40763 43258 40772
rect 45296 40458 45324 53926
rect 46124 41274 46152 53926
rect 46676 53582 46704 56200
rect 47320 54194 47348 56200
rect 47964 55214 47992 56200
rect 47872 55186 47992 55214
rect 47872 54194 47900 55186
rect 47950 54428 48258 54437
rect 47950 54426 47956 54428
rect 48012 54426 48036 54428
rect 48092 54426 48116 54428
rect 48172 54426 48196 54428
rect 48252 54426 48258 54428
rect 48012 54374 48014 54426
rect 48194 54374 48196 54426
rect 47950 54372 47956 54374
rect 48012 54372 48036 54374
rect 48092 54372 48116 54374
rect 48172 54372 48196 54374
rect 48252 54372 48258 54374
rect 47950 54363 48258 54372
rect 47308 54188 47360 54194
rect 47308 54130 47360 54136
rect 47860 54188 47912 54194
rect 47860 54130 47912 54136
rect 46848 53984 46900 53990
rect 46848 53926 46900 53932
rect 47768 53984 47820 53990
rect 47768 53926 47820 53932
rect 46664 53576 46716 53582
rect 46664 53518 46716 53524
rect 46860 44878 46888 53926
rect 46940 53440 46992 53446
rect 46940 53382 46992 53388
rect 47032 53440 47084 53446
rect 47032 53382 47084 53388
rect 46848 44872 46900 44878
rect 46848 44814 46900 44820
rect 46112 41268 46164 41274
rect 46112 41210 46164 41216
rect 45284 40452 45336 40458
rect 45284 40394 45336 40400
rect 46952 40390 46980 53382
rect 47044 50862 47072 53382
rect 47032 50856 47084 50862
rect 47032 50798 47084 50804
rect 47780 41138 47808 53926
rect 48608 53582 48636 56200
rect 49054 54632 49110 54641
rect 49054 54567 49110 54576
rect 48688 53984 48740 53990
rect 48688 53926 48740 53932
rect 48596 53576 48648 53582
rect 48596 53518 48648 53524
rect 47950 53340 48258 53349
rect 47950 53338 47956 53340
rect 48012 53338 48036 53340
rect 48092 53338 48116 53340
rect 48172 53338 48196 53340
rect 48252 53338 48258 53340
rect 48012 53286 48014 53338
rect 48194 53286 48196 53338
rect 47950 53284 47956 53286
rect 48012 53284 48036 53286
rect 48092 53284 48116 53286
rect 48172 53284 48196 53286
rect 48252 53284 48258 53286
rect 47950 53275 48258 53284
rect 47950 52252 48258 52261
rect 47950 52250 47956 52252
rect 48012 52250 48036 52252
rect 48092 52250 48116 52252
rect 48172 52250 48196 52252
rect 48252 52250 48258 52252
rect 48012 52198 48014 52250
rect 48194 52198 48196 52250
rect 47950 52196 47956 52198
rect 48012 52196 48036 52198
rect 48092 52196 48116 52198
rect 48172 52196 48196 52198
rect 48252 52196 48258 52198
rect 47950 52187 48258 52196
rect 47950 51164 48258 51173
rect 47950 51162 47956 51164
rect 48012 51162 48036 51164
rect 48092 51162 48116 51164
rect 48172 51162 48196 51164
rect 48252 51162 48258 51164
rect 48012 51110 48014 51162
rect 48194 51110 48196 51162
rect 47950 51108 47956 51110
rect 48012 51108 48036 51110
rect 48092 51108 48116 51110
rect 48172 51108 48196 51110
rect 48252 51108 48258 51110
rect 47950 51099 48258 51108
rect 47950 50076 48258 50085
rect 47950 50074 47956 50076
rect 48012 50074 48036 50076
rect 48092 50074 48116 50076
rect 48172 50074 48196 50076
rect 48252 50074 48258 50076
rect 48012 50022 48014 50074
rect 48194 50022 48196 50074
rect 47950 50020 47956 50022
rect 48012 50020 48036 50022
rect 48092 50020 48116 50022
rect 48172 50020 48196 50022
rect 48252 50020 48258 50022
rect 47950 50011 48258 50020
rect 47950 48988 48258 48997
rect 47950 48986 47956 48988
rect 48012 48986 48036 48988
rect 48092 48986 48116 48988
rect 48172 48986 48196 48988
rect 48252 48986 48258 48988
rect 48012 48934 48014 48986
rect 48194 48934 48196 48986
rect 47950 48932 47956 48934
rect 48012 48932 48036 48934
rect 48092 48932 48116 48934
rect 48172 48932 48196 48934
rect 48252 48932 48258 48934
rect 47950 48923 48258 48932
rect 47950 47900 48258 47909
rect 47950 47898 47956 47900
rect 48012 47898 48036 47900
rect 48092 47898 48116 47900
rect 48172 47898 48196 47900
rect 48252 47898 48258 47900
rect 48012 47846 48014 47898
rect 48194 47846 48196 47898
rect 47950 47844 47956 47846
rect 48012 47844 48036 47846
rect 48092 47844 48116 47846
rect 48172 47844 48196 47846
rect 48252 47844 48258 47846
rect 47950 47835 48258 47844
rect 47950 46812 48258 46821
rect 47950 46810 47956 46812
rect 48012 46810 48036 46812
rect 48092 46810 48116 46812
rect 48172 46810 48196 46812
rect 48252 46810 48258 46812
rect 48012 46758 48014 46810
rect 48194 46758 48196 46810
rect 47950 46756 47956 46758
rect 48012 46756 48036 46758
rect 48092 46756 48116 46758
rect 48172 46756 48196 46758
rect 48252 46756 48258 46758
rect 47950 46747 48258 46756
rect 47860 45960 47912 45966
rect 47860 45902 47912 45908
rect 47768 41132 47820 41138
rect 47768 41074 47820 41080
rect 46940 40384 46992 40390
rect 46940 40326 46992 40332
rect 38660 39840 38712 39846
rect 38660 39782 38712 39788
rect 42950 39740 43258 39749
rect 42950 39738 42956 39740
rect 43012 39738 43036 39740
rect 43092 39738 43116 39740
rect 43172 39738 43196 39740
rect 43252 39738 43258 39740
rect 43012 39686 43014 39738
rect 43194 39686 43196 39738
rect 42950 39684 42956 39686
rect 43012 39684 43036 39686
rect 43092 39684 43116 39686
rect 43172 39684 43196 39686
rect 43252 39684 43258 39686
rect 42950 39675 43258 39684
rect 37832 39636 37884 39642
rect 37832 39578 37884 39584
rect 37950 39196 38258 39205
rect 37950 39194 37956 39196
rect 38012 39194 38036 39196
rect 38092 39194 38116 39196
rect 38172 39194 38196 39196
rect 38252 39194 38258 39196
rect 38012 39142 38014 39194
rect 38194 39142 38196 39194
rect 37950 39140 37956 39142
rect 38012 39140 38036 39142
rect 38092 39140 38116 39142
rect 38172 39140 38196 39142
rect 38252 39140 38258 39142
rect 37950 39131 38258 39140
rect 42950 38652 43258 38661
rect 42950 38650 42956 38652
rect 43012 38650 43036 38652
rect 43092 38650 43116 38652
rect 43172 38650 43196 38652
rect 43252 38650 43258 38652
rect 43012 38598 43014 38650
rect 43194 38598 43196 38650
rect 42950 38596 42956 38598
rect 43012 38596 43036 38598
rect 43092 38596 43116 38598
rect 43172 38596 43196 38598
rect 43252 38596 43258 38598
rect 42950 38587 43258 38596
rect 37950 38108 38258 38117
rect 37950 38106 37956 38108
rect 38012 38106 38036 38108
rect 38092 38106 38116 38108
rect 38172 38106 38196 38108
rect 38252 38106 38258 38108
rect 38012 38054 38014 38106
rect 38194 38054 38196 38106
rect 37950 38052 37956 38054
rect 38012 38052 38036 38054
rect 38092 38052 38116 38054
rect 38172 38052 38196 38054
rect 38252 38052 38258 38054
rect 37950 38043 38258 38052
rect 42950 37564 43258 37573
rect 42950 37562 42956 37564
rect 43012 37562 43036 37564
rect 43092 37562 43116 37564
rect 43172 37562 43196 37564
rect 43252 37562 43258 37564
rect 43012 37510 43014 37562
rect 43194 37510 43196 37562
rect 42950 37508 42956 37510
rect 43012 37508 43036 37510
rect 43092 37508 43116 37510
rect 43172 37508 43196 37510
rect 43252 37508 43258 37510
rect 42950 37499 43258 37508
rect 37950 37020 38258 37029
rect 37950 37018 37956 37020
rect 38012 37018 38036 37020
rect 38092 37018 38116 37020
rect 38172 37018 38196 37020
rect 38252 37018 38258 37020
rect 38012 36966 38014 37018
rect 38194 36966 38196 37018
rect 37950 36964 37956 36966
rect 38012 36964 38036 36966
rect 38092 36964 38116 36966
rect 38172 36964 38196 36966
rect 38252 36964 38258 36966
rect 37950 36955 38258 36964
rect 42950 36476 43258 36485
rect 42950 36474 42956 36476
rect 43012 36474 43036 36476
rect 43092 36474 43116 36476
rect 43172 36474 43196 36476
rect 43252 36474 43258 36476
rect 43012 36422 43014 36474
rect 43194 36422 43196 36474
rect 42950 36420 42956 36422
rect 43012 36420 43036 36422
rect 43092 36420 43116 36422
rect 43172 36420 43196 36422
rect 43252 36420 43258 36422
rect 42950 36411 43258 36420
rect 37950 35932 38258 35941
rect 37950 35930 37956 35932
rect 38012 35930 38036 35932
rect 38092 35930 38116 35932
rect 38172 35930 38196 35932
rect 38252 35930 38258 35932
rect 38012 35878 38014 35930
rect 38194 35878 38196 35930
rect 37950 35876 37956 35878
rect 38012 35876 38036 35878
rect 38092 35876 38116 35878
rect 38172 35876 38196 35878
rect 38252 35876 38258 35878
rect 37950 35867 38258 35876
rect 42950 35388 43258 35397
rect 42950 35386 42956 35388
rect 43012 35386 43036 35388
rect 43092 35386 43116 35388
rect 43172 35386 43196 35388
rect 43252 35386 43258 35388
rect 43012 35334 43014 35386
rect 43194 35334 43196 35386
rect 42950 35332 42956 35334
rect 43012 35332 43036 35334
rect 43092 35332 43116 35334
rect 43172 35332 43196 35334
rect 43252 35332 43258 35334
rect 42950 35323 43258 35332
rect 37950 34844 38258 34853
rect 37950 34842 37956 34844
rect 38012 34842 38036 34844
rect 38092 34842 38116 34844
rect 38172 34842 38196 34844
rect 38252 34842 38258 34844
rect 38012 34790 38014 34842
rect 38194 34790 38196 34842
rect 37950 34788 37956 34790
rect 38012 34788 38036 34790
rect 38092 34788 38116 34790
rect 38172 34788 38196 34790
rect 38252 34788 38258 34790
rect 37950 34779 38258 34788
rect 42950 34300 43258 34309
rect 42950 34298 42956 34300
rect 43012 34298 43036 34300
rect 43092 34298 43116 34300
rect 43172 34298 43196 34300
rect 43252 34298 43258 34300
rect 43012 34246 43014 34298
rect 43194 34246 43196 34298
rect 42950 34244 42956 34246
rect 43012 34244 43036 34246
rect 43092 34244 43116 34246
rect 43172 34244 43196 34246
rect 43252 34244 43258 34246
rect 42950 34235 43258 34244
rect 37950 33756 38258 33765
rect 37950 33754 37956 33756
rect 38012 33754 38036 33756
rect 38092 33754 38116 33756
rect 38172 33754 38196 33756
rect 38252 33754 38258 33756
rect 38012 33702 38014 33754
rect 38194 33702 38196 33754
rect 37950 33700 37956 33702
rect 38012 33700 38036 33702
rect 38092 33700 38116 33702
rect 38172 33700 38196 33702
rect 38252 33700 38258 33702
rect 37950 33691 38258 33700
rect 42950 33212 43258 33221
rect 42950 33210 42956 33212
rect 43012 33210 43036 33212
rect 43092 33210 43116 33212
rect 43172 33210 43196 33212
rect 43252 33210 43258 33212
rect 43012 33158 43014 33210
rect 43194 33158 43196 33210
rect 42950 33156 42956 33158
rect 43012 33156 43036 33158
rect 43092 33156 43116 33158
rect 43172 33156 43196 33158
rect 43252 33156 43258 33158
rect 42950 33147 43258 33156
rect 37950 32668 38258 32677
rect 37950 32666 37956 32668
rect 38012 32666 38036 32668
rect 38092 32666 38116 32668
rect 38172 32666 38196 32668
rect 38252 32666 38258 32668
rect 38012 32614 38014 32666
rect 38194 32614 38196 32666
rect 37950 32612 37956 32614
rect 38012 32612 38036 32614
rect 38092 32612 38116 32614
rect 38172 32612 38196 32614
rect 38252 32612 38258 32614
rect 37950 32603 38258 32612
rect 42950 32124 43258 32133
rect 42950 32122 42956 32124
rect 43012 32122 43036 32124
rect 43092 32122 43116 32124
rect 43172 32122 43196 32124
rect 43252 32122 43258 32124
rect 43012 32070 43014 32122
rect 43194 32070 43196 32122
rect 42950 32068 42956 32070
rect 43012 32068 43036 32070
rect 43092 32068 43116 32070
rect 43172 32068 43196 32070
rect 43252 32068 43258 32070
rect 42950 32059 43258 32068
rect 37950 31580 38258 31589
rect 37950 31578 37956 31580
rect 38012 31578 38036 31580
rect 38092 31578 38116 31580
rect 38172 31578 38196 31580
rect 38252 31578 38258 31580
rect 38012 31526 38014 31578
rect 38194 31526 38196 31578
rect 37950 31524 37956 31526
rect 38012 31524 38036 31526
rect 38092 31524 38116 31526
rect 38172 31524 38196 31526
rect 38252 31524 38258 31526
rect 37950 31515 38258 31524
rect 42950 31036 43258 31045
rect 42950 31034 42956 31036
rect 43012 31034 43036 31036
rect 43092 31034 43116 31036
rect 43172 31034 43196 31036
rect 43252 31034 43258 31036
rect 43012 30982 43014 31034
rect 43194 30982 43196 31034
rect 42950 30980 42956 30982
rect 43012 30980 43036 30982
rect 43092 30980 43116 30982
rect 43172 30980 43196 30982
rect 43252 30980 43258 30982
rect 42950 30971 43258 30980
rect 37950 30492 38258 30501
rect 37950 30490 37956 30492
rect 38012 30490 38036 30492
rect 38092 30490 38116 30492
rect 38172 30490 38196 30492
rect 38252 30490 38258 30492
rect 38012 30438 38014 30490
rect 38194 30438 38196 30490
rect 37950 30436 37956 30438
rect 38012 30436 38036 30438
rect 38092 30436 38116 30438
rect 38172 30436 38196 30438
rect 38252 30436 38258 30438
rect 37950 30427 38258 30436
rect 42950 29948 43258 29957
rect 42950 29946 42956 29948
rect 43012 29946 43036 29948
rect 43092 29946 43116 29948
rect 43172 29946 43196 29948
rect 43252 29946 43258 29948
rect 43012 29894 43014 29946
rect 43194 29894 43196 29946
rect 42950 29892 42956 29894
rect 43012 29892 43036 29894
rect 43092 29892 43116 29894
rect 43172 29892 43196 29894
rect 43252 29892 43258 29894
rect 42950 29883 43258 29892
rect 37950 29404 38258 29413
rect 37950 29402 37956 29404
rect 38012 29402 38036 29404
rect 38092 29402 38116 29404
rect 38172 29402 38196 29404
rect 38252 29402 38258 29404
rect 38012 29350 38014 29402
rect 38194 29350 38196 29402
rect 37950 29348 37956 29350
rect 38012 29348 38036 29350
rect 38092 29348 38116 29350
rect 38172 29348 38196 29350
rect 38252 29348 38258 29350
rect 37950 29339 38258 29348
rect 42950 28860 43258 28869
rect 42950 28858 42956 28860
rect 43012 28858 43036 28860
rect 43092 28858 43116 28860
rect 43172 28858 43196 28860
rect 43252 28858 43258 28860
rect 43012 28806 43014 28858
rect 43194 28806 43196 28858
rect 42950 28804 42956 28806
rect 43012 28804 43036 28806
rect 43092 28804 43116 28806
rect 43172 28804 43196 28806
rect 43252 28804 43258 28806
rect 42950 28795 43258 28804
rect 37950 28316 38258 28325
rect 37950 28314 37956 28316
rect 38012 28314 38036 28316
rect 38092 28314 38116 28316
rect 38172 28314 38196 28316
rect 38252 28314 38258 28316
rect 38012 28262 38014 28314
rect 38194 28262 38196 28314
rect 37950 28260 37956 28262
rect 38012 28260 38036 28262
rect 38092 28260 38116 28262
rect 38172 28260 38196 28262
rect 38252 28260 38258 28262
rect 37950 28251 38258 28260
rect 42950 27772 43258 27781
rect 42950 27770 42956 27772
rect 43012 27770 43036 27772
rect 43092 27770 43116 27772
rect 43172 27770 43196 27772
rect 43252 27770 43258 27772
rect 43012 27718 43014 27770
rect 43194 27718 43196 27770
rect 42950 27716 42956 27718
rect 43012 27716 43036 27718
rect 43092 27716 43116 27718
rect 43172 27716 43196 27718
rect 43252 27716 43258 27718
rect 42950 27707 43258 27716
rect 37950 27228 38258 27237
rect 37950 27226 37956 27228
rect 38012 27226 38036 27228
rect 38092 27226 38116 27228
rect 38172 27226 38196 27228
rect 38252 27226 38258 27228
rect 38012 27174 38014 27226
rect 38194 27174 38196 27226
rect 37950 27172 37956 27174
rect 38012 27172 38036 27174
rect 38092 27172 38116 27174
rect 38172 27172 38196 27174
rect 38252 27172 38258 27174
rect 37950 27163 38258 27172
rect 42950 26684 43258 26693
rect 42950 26682 42956 26684
rect 43012 26682 43036 26684
rect 43092 26682 43116 26684
rect 43172 26682 43196 26684
rect 43252 26682 43258 26684
rect 43012 26630 43014 26682
rect 43194 26630 43196 26682
rect 42950 26628 42956 26630
rect 43012 26628 43036 26630
rect 43092 26628 43116 26630
rect 43172 26628 43196 26630
rect 43252 26628 43258 26630
rect 42950 26619 43258 26628
rect 37950 26140 38258 26149
rect 37950 26138 37956 26140
rect 38012 26138 38036 26140
rect 38092 26138 38116 26140
rect 38172 26138 38196 26140
rect 38252 26138 38258 26140
rect 38012 26086 38014 26138
rect 38194 26086 38196 26138
rect 37950 26084 37956 26086
rect 38012 26084 38036 26086
rect 38092 26084 38116 26086
rect 38172 26084 38196 26086
rect 38252 26084 38258 26086
rect 37950 26075 38258 26084
rect 42950 25596 43258 25605
rect 42950 25594 42956 25596
rect 43012 25594 43036 25596
rect 43092 25594 43116 25596
rect 43172 25594 43196 25596
rect 43252 25594 43258 25596
rect 43012 25542 43014 25594
rect 43194 25542 43196 25594
rect 42950 25540 42956 25542
rect 43012 25540 43036 25542
rect 43092 25540 43116 25542
rect 43172 25540 43196 25542
rect 43252 25540 43258 25542
rect 42950 25531 43258 25540
rect 37950 25052 38258 25061
rect 37950 25050 37956 25052
rect 38012 25050 38036 25052
rect 38092 25050 38116 25052
rect 38172 25050 38196 25052
rect 38252 25050 38258 25052
rect 38012 24998 38014 25050
rect 38194 24998 38196 25050
rect 37950 24996 37956 24998
rect 38012 24996 38036 24998
rect 38092 24996 38116 24998
rect 38172 24996 38196 24998
rect 38252 24996 38258 24998
rect 37950 24987 38258 24996
rect 33692 24812 33744 24818
rect 33692 24754 33744 24760
rect 47872 24750 47900 45902
rect 47950 45724 48258 45733
rect 47950 45722 47956 45724
rect 48012 45722 48036 45724
rect 48092 45722 48116 45724
rect 48172 45722 48196 45724
rect 48252 45722 48258 45724
rect 48012 45670 48014 45722
rect 48194 45670 48196 45722
rect 47950 45668 47956 45670
rect 48012 45668 48036 45670
rect 48092 45668 48116 45670
rect 48172 45668 48196 45670
rect 48252 45668 48258 45670
rect 47950 45659 48258 45668
rect 48700 45554 48728 53926
rect 48872 53440 48924 53446
rect 48872 53382 48924 53388
rect 48780 52896 48832 52902
rect 48780 52838 48832 52844
rect 48608 45526 48728 45554
rect 47950 44636 48258 44645
rect 47950 44634 47956 44636
rect 48012 44634 48036 44636
rect 48092 44634 48116 44636
rect 48172 44634 48196 44636
rect 48252 44634 48258 44636
rect 48012 44582 48014 44634
rect 48194 44582 48196 44634
rect 47950 44580 47956 44582
rect 48012 44580 48036 44582
rect 48092 44580 48116 44582
rect 48172 44580 48196 44582
rect 48252 44580 48258 44582
rect 47950 44571 48258 44580
rect 48608 43722 48636 45526
rect 48596 43716 48648 43722
rect 48596 43658 48648 43664
rect 47950 43548 48258 43557
rect 47950 43546 47956 43548
rect 48012 43546 48036 43548
rect 48092 43546 48116 43548
rect 48172 43546 48196 43548
rect 48252 43546 48258 43548
rect 48012 43494 48014 43546
rect 48194 43494 48196 43546
rect 47950 43492 47956 43494
rect 48012 43492 48036 43494
rect 48092 43492 48116 43494
rect 48172 43492 48196 43494
rect 48252 43492 48258 43494
rect 47950 43483 48258 43492
rect 48792 42770 48820 52838
rect 48780 42764 48832 42770
rect 48780 42706 48832 42712
rect 47950 42460 48258 42469
rect 47950 42458 47956 42460
rect 48012 42458 48036 42460
rect 48092 42458 48116 42460
rect 48172 42458 48196 42460
rect 48252 42458 48258 42460
rect 48012 42406 48014 42458
rect 48194 42406 48196 42458
rect 47950 42404 47956 42406
rect 48012 42404 48036 42406
rect 48092 42404 48116 42406
rect 48172 42404 48196 42406
rect 48252 42404 48258 42406
rect 47950 42395 48258 42404
rect 47950 41372 48258 41381
rect 47950 41370 47956 41372
rect 48012 41370 48036 41372
rect 48092 41370 48116 41372
rect 48172 41370 48196 41372
rect 48252 41370 48258 41372
rect 48012 41318 48014 41370
rect 48194 41318 48196 41370
rect 47950 41316 47956 41318
rect 48012 41316 48036 41318
rect 48092 41316 48116 41318
rect 48172 41316 48196 41318
rect 48252 41316 48258 41318
rect 47950 41307 48258 41316
rect 47950 40284 48258 40293
rect 47950 40282 47956 40284
rect 48012 40282 48036 40284
rect 48092 40282 48116 40284
rect 48172 40282 48196 40284
rect 48252 40282 48258 40284
rect 48012 40230 48014 40282
rect 48194 40230 48196 40282
rect 47950 40228 47956 40230
rect 48012 40228 48036 40230
rect 48092 40228 48116 40230
rect 48172 40228 48196 40230
rect 48252 40228 48258 40230
rect 47950 40219 48258 40228
rect 47950 39196 48258 39205
rect 47950 39194 47956 39196
rect 48012 39194 48036 39196
rect 48092 39194 48116 39196
rect 48172 39194 48196 39196
rect 48252 39194 48258 39196
rect 48012 39142 48014 39194
rect 48194 39142 48196 39194
rect 47950 39140 47956 39142
rect 48012 39140 48036 39142
rect 48092 39140 48116 39142
rect 48172 39140 48196 39142
rect 48252 39140 48258 39142
rect 47950 39131 48258 39140
rect 48884 38894 48912 53382
rect 49068 53106 49096 54567
rect 49252 53650 49280 56200
rect 49240 53644 49292 53650
rect 49240 53586 49292 53592
rect 49056 53100 49108 53106
rect 49056 53042 49108 53048
rect 49148 52624 49200 52630
rect 49148 52566 49200 52572
rect 49056 52488 49108 52494
rect 49054 52456 49056 52465
rect 49108 52456 49110 52465
rect 49054 52391 49110 52400
rect 49056 50312 49108 50318
rect 49054 50280 49056 50289
rect 49108 50280 49110 50289
rect 49054 50215 49110 50224
rect 48962 48104 49018 48113
rect 48962 48039 48964 48048
rect 49016 48039 49018 48048
rect 48964 48010 49016 48016
rect 49056 48000 49108 48006
rect 49056 47942 49108 47948
rect 48964 47796 49016 47802
rect 48964 47738 49016 47744
rect 48976 42090 49004 47738
rect 48964 42084 49016 42090
rect 48964 42026 49016 42032
rect 49068 40730 49096 47942
rect 49160 47802 49188 52566
rect 49240 50176 49292 50182
rect 49240 50118 49292 50124
rect 49148 47796 49200 47802
rect 49148 47738 49200 47744
rect 49148 45960 49200 45966
rect 49146 45928 49148 45937
rect 49200 45928 49202 45937
rect 49146 45863 49202 45872
rect 49252 43654 49280 50118
rect 49240 43648 49292 43654
rect 49240 43590 49292 43596
rect 49056 40724 49108 40730
rect 49056 40666 49108 40672
rect 48872 38888 48924 38894
rect 48872 38830 48924 38836
rect 47950 38108 48258 38117
rect 47950 38106 47956 38108
rect 48012 38106 48036 38108
rect 48092 38106 48116 38108
rect 48172 38106 48196 38108
rect 48252 38106 48258 38108
rect 48012 38054 48014 38106
rect 48194 38054 48196 38106
rect 47950 38052 47956 38054
rect 48012 38052 48036 38054
rect 48092 38052 48116 38054
rect 48172 38052 48196 38054
rect 48252 38052 48258 38054
rect 47950 38043 48258 38052
rect 47950 37020 48258 37029
rect 47950 37018 47956 37020
rect 48012 37018 48036 37020
rect 48092 37018 48116 37020
rect 48172 37018 48196 37020
rect 48252 37018 48258 37020
rect 48012 36966 48014 37018
rect 48194 36966 48196 37018
rect 47950 36964 47956 36966
rect 48012 36964 48036 36966
rect 48092 36964 48116 36966
rect 48172 36964 48196 36966
rect 48252 36964 48258 36966
rect 47950 36955 48258 36964
rect 47950 35932 48258 35941
rect 47950 35930 47956 35932
rect 48012 35930 48036 35932
rect 48092 35930 48116 35932
rect 48172 35930 48196 35932
rect 48252 35930 48258 35932
rect 48012 35878 48014 35930
rect 48194 35878 48196 35930
rect 47950 35876 47956 35878
rect 48012 35876 48036 35878
rect 48092 35876 48116 35878
rect 48172 35876 48196 35878
rect 48252 35876 48258 35878
rect 47950 35867 48258 35876
rect 47950 34844 48258 34853
rect 47950 34842 47956 34844
rect 48012 34842 48036 34844
rect 48092 34842 48116 34844
rect 48172 34842 48196 34844
rect 48252 34842 48258 34844
rect 48012 34790 48014 34842
rect 48194 34790 48196 34842
rect 47950 34788 47956 34790
rect 48012 34788 48036 34790
rect 48092 34788 48116 34790
rect 48172 34788 48196 34790
rect 48252 34788 48258 34790
rect 47950 34779 48258 34788
rect 47950 33756 48258 33765
rect 47950 33754 47956 33756
rect 48012 33754 48036 33756
rect 48092 33754 48116 33756
rect 48172 33754 48196 33756
rect 48252 33754 48258 33756
rect 48012 33702 48014 33754
rect 48194 33702 48196 33754
rect 47950 33700 47956 33702
rect 48012 33700 48036 33702
rect 48092 33700 48116 33702
rect 48172 33700 48196 33702
rect 48252 33700 48258 33702
rect 47950 33691 48258 33700
rect 47950 32668 48258 32677
rect 47950 32666 47956 32668
rect 48012 32666 48036 32668
rect 48092 32666 48116 32668
rect 48172 32666 48196 32668
rect 48252 32666 48258 32668
rect 48012 32614 48014 32666
rect 48194 32614 48196 32666
rect 47950 32612 47956 32614
rect 48012 32612 48036 32614
rect 48092 32612 48116 32614
rect 48172 32612 48196 32614
rect 48252 32612 48258 32614
rect 47950 32603 48258 32612
rect 47950 31580 48258 31589
rect 47950 31578 47956 31580
rect 48012 31578 48036 31580
rect 48092 31578 48116 31580
rect 48172 31578 48196 31580
rect 48252 31578 48258 31580
rect 48012 31526 48014 31578
rect 48194 31526 48196 31578
rect 47950 31524 47956 31526
rect 48012 31524 48036 31526
rect 48092 31524 48116 31526
rect 48172 31524 48196 31526
rect 48252 31524 48258 31526
rect 47950 31515 48258 31524
rect 47950 30492 48258 30501
rect 47950 30490 47956 30492
rect 48012 30490 48036 30492
rect 48092 30490 48116 30492
rect 48172 30490 48196 30492
rect 48252 30490 48258 30492
rect 48012 30438 48014 30490
rect 48194 30438 48196 30490
rect 47950 30436 47956 30438
rect 48012 30436 48036 30438
rect 48092 30436 48116 30438
rect 48172 30436 48196 30438
rect 48252 30436 48258 30438
rect 47950 30427 48258 30436
rect 47950 29404 48258 29413
rect 47950 29402 47956 29404
rect 48012 29402 48036 29404
rect 48092 29402 48116 29404
rect 48172 29402 48196 29404
rect 48252 29402 48258 29404
rect 48012 29350 48014 29402
rect 48194 29350 48196 29402
rect 47950 29348 47956 29350
rect 48012 29348 48036 29350
rect 48092 29348 48116 29350
rect 48172 29348 48196 29350
rect 48252 29348 48258 29350
rect 47950 29339 48258 29348
rect 47950 28316 48258 28325
rect 47950 28314 47956 28316
rect 48012 28314 48036 28316
rect 48092 28314 48116 28316
rect 48172 28314 48196 28316
rect 48252 28314 48258 28316
rect 48012 28262 48014 28314
rect 48194 28262 48196 28314
rect 47950 28260 47956 28262
rect 48012 28260 48036 28262
rect 48092 28260 48116 28262
rect 48172 28260 48196 28262
rect 48252 28260 48258 28262
rect 47950 28251 48258 28260
rect 47950 27228 48258 27237
rect 47950 27226 47956 27228
rect 48012 27226 48036 27228
rect 48092 27226 48116 27228
rect 48172 27226 48196 27228
rect 48252 27226 48258 27228
rect 48012 27174 48014 27226
rect 48194 27174 48196 27226
rect 47950 27172 47956 27174
rect 48012 27172 48036 27174
rect 48092 27172 48116 27174
rect 48172 27172 48196 27174
rect 48252 27172 48258 27174
rect 47950 27163 48258 27172
rect 47950 26140 48258 26149
rect 47950 26138 47956 26140
rect 48012 26138 48036 26140
rect 48092 26138 48116 26140
rect 48172 26138 48196 26140
rect 48252 26138 48258 26140
rect 48012 26086 48014 26138
rect 48194 26086 48196 26138
rect 47950 26084 47956 26086
rect 48012 26084 48036 26086
rect 48092 26084 48116 26086
rect 48172 26084 48196 26086
rect 48252 26084 48258 26086
rect 47950 26075 48258 26084
rect 47950 25052 48258 25061
rect 47950 25050 47956 25052
rect 48012 25050 48036 25052
rect 48092 25050 48116 25052
rect 48172 25050 48196 25052
rect 48252 25050 48258 25052
rect 48012 24998 48014 25050
rect 48194 24998 48196 25050
rect 47950 24996 47956 24998
rect 48012 24996 48036 24998
rect 48092 24996 48116 24998
rect 48172 24996 48196 24998
rect 48252 24996 48258 24998
rect 47950 24987 48258 24996
rect 34336 24744 34388 24750
rect 34336 24686 34388 24692
rect 47860 24744 47912 24750
rect 47860 24686 47912 24692
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 34348 20262 34376 24686
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 34336 20256 34388 20262
rect 34336 20198 34388 20204
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 32864 16584 32916 16590
rect 32864 16526 32916 16532
rect 31208 16516 31260 16522
rect 31208 16458 31260 16464
rect 31220 14074 31248 16458
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 47950 15260 48258 15269
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 31208 14068 31260 14074
rect 31208 14010 31260 14016
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 45560 13184 45612 13190
rect 45560 13126 45612 13132
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 45572 2650 45600 13126
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 47950 11996 48258 12005
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 48596 3052 48648 3058
rect 48596 2994 48648 3000
rect 31024 2644 31076 2650
rect 31024 2586 31076 2592
rect 45560 2644 45612 2650
rect 45560 2586 45612 2592
rect 28908 2576 28960 2582
rect 28908 2518 28960 2524
rect 32036 2440 32088 2446
rect 32036 2382 32088 2388
rect 35348 2440 35400 2446
rect 35348 2382 35400 2388
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 41972 2440 42024 2446
rect 41972 2382 42024 2388
rect 32048 800 32076 2382
rect 35360 800 35388 2382
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 38672 800 38700 2382
rect 41984 800 42012 2382
rect 45284 2372 45336 2378
rect 45284 2314 45336 2320
rect 45296 800 45324 2314
rect 47950 2204 48258 2213
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 48608 800 48636 2994
rect 2226 0 2282 800
rect 5538 0 5594 800
rect 8850 0 8906 800
rect 12162 0 12218 800
rect 15474 0 15530 800
rect 18786 0 18842 800
rect 22098 0 22154 800
rect 25410 0 25466 800
rect 28722 0 28778 800
rect 32034 0 32090 800
rect 35346 0 35402 800
rect 38658 0 38714 800
rect 41970 0 42026 800
rect 45282 0 45338 800
rect 48594 0 48650 800
<< via2 >>
rect 1306 51312 1362 51368
rect 1306 50496 1362 50552
rect 1306 49716 1308 49736
rect 1308 49716 1360 49736
rect 1360 49716 1362 49736
rect 1306 49680 1362 49716
rect 1306 48864 1362 48920
rect 1306 48048 1362 48104
rect 1306 47232 1362 47288
rect 1306 46452 1308 46472
rect 1308 46452 1360 46472
rect 1360 46452 1362 46472
rect 1306 46416 1362 46452
rect 1306 45600 1362 45656
rect 1306 44784 1362 44840
rect 1306 43188 1308 43208
rect 1308 43188 1360 43208
rect 1360 43188 1362 43208
rect 1306 43152 1362 43188
rect 2778 53760 2834 53816
rect 3422 54576 3478 54632
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 3330 52128 3386 52184
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 3606 52944 3662 53000
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 2042 43968 2098 44024
rect 1306 42336 1362 42392
rect 1306 41520 1362 41576
rect 1306 40704 1362 40760
rect 1306 39072 1362 39128
rect 1306 38256 1362 38312
rect 1306 37440 1362 37496
rect 2042 39924 2044 39944
rect 2044 39924 2096 39944
rect 2096 39924 2098 39944
rect 2042 39888 2098 39924
rect 1306 36660 1308 36680
rect 1308 36660 1360 36680
rect 1360 36660 1362 36680
rect 1306 36624 1362 36660
rect 1306 34992 1362 35048
rect 1306 33396 1308 33416
rect 1308 33396 1360 33416
rect 1360 33396 1362 33416
rect 1306 33360 1362 33396
rect 1306 32544 1362 32600
rect 1306 31728 1362 31784
rect 1306 30912 1362 30968
rect 1306 30132 1308 30152
rect 1308 30132 1360 30152
rect 1360 30132 1362 30152
rect 1306 30096 1362 30132
rect 1306 29280 1362 29336
rect 1766 28600 1822 28656
rect 1306 28464 1362 28520
rect 1306 27648 1362 27704
rect 938 26832 994 26888
rect 1582 26016 1638 26072
rect 938 25236 940 25256
rect 940 25236 992 25256
rect 992 25236 994 25256
rect 938 25200 994 25236
rect 938 24384 994 24440
rect 938 23604 940 23624
rect 940 23604 992 23624
rect 992 23604 994 23624
rect 938 23568 994 23604
rect 938 22752 994 22808
rect 938 21972 940 21992
rect 940 21972 992 21992
rect 992 21972 994 21992
rect 938 21936 994 21972
rect 938 21120 994 21176
rect 938 20340 940 20360
rect 940 20340 992 20360
rect 992 20340 994 20360
rect 938 20304 994 20340
rect 938 19488 994 19544
rect 938 18708 940 18728
rect 940 18708 992 18728
rect 992 18708 994 18728
rect 938 18672 994 18708
rect 938 17040 994 17096
rect 938 16224 994 16280
rect 938 15428 994 15464
rect 938 15408 940 15428
rect 940 15408 992 15428
rect 992 15408 994 15428
rect 938 14592 994 14648
rect 938 13776 994 13832
rect 938 12960 994 13016
rect 938 12164 994 12200
rect 938 12144 940 12164
rect 940 12144 992 12164
rect 992 12144 994 12164
rect 938 11328 994 11384
rect 938 10512 994 10568
rect 938 9696 994 9752
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 3514 45464 3570 45520
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 2778 35808 2834 35864
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 2042 34176 2098 34232
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 6274 37304 6330 37360
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 7102 36660 7104 36680
rect 7104 36660 7156 36680
rect 7156 36660 7158 36680
rect 7102 36624 7158 36660
rect 7378 37440 7434 37496
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7470 36760 7526 36816
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 8206 36624 8262 36680
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 8114 35012 8170 35048
rect 8114 34992 8116 35012
rect 8116 34992 8168 35012
rect 8168 34992 8170 35012
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 1858 20304 1914 20360
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 1766 17856 1822 17912
rect 1950 17720 2006 17776
rect 1858 17076 1860 17096
rect 1860 17076 1912 17096
rect 1912 17076 1914 17096
rect 1858 17040 1914 17076
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 938 8916 940 8936
rect 940 8916 992 8936
rect 992 8916 994 8936
rect 938 8880 994 8916
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 1766 8064 1822 8120
rect 938 7248 994 7304
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 938 6432 994 6488
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 938 5636 994 5672
rect 938 5616 940 5636
rect 940 5616 992 5636
rect 992 5616 994 5636
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 938 4800 994 4856
rect 938 4020 940 4040
rect 940 4020 992 4040
rect 992 4020 994 4040
rect 938 3984 994 4020
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 938 3168 994 3224
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 9218 43152 9274 43208
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 9126 38664 9182 38720
rect 9034 37304 9090 37360
rect 9310 37440 9366 37496
rect 9862 40432 9918 40488
rect 9678 37440 9734 37496
rect 9218 32564 9274 32600
rect 9218 32544 9220 32564
rect 9220 32544 9272 32564
rect 9272 32544 9274 32564
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 9586 36916 9642 36952
rect 9586 36896 9588 36916
rect 9588 36896 9640 36916
rect 9640 36896 9642 36916
rect 9586 36660 9588 36680
rect 9588 36660 9640 36680
rect 9640 36660 9642 36680
rect 9586 36624 9642 36660
rect 10506 39480 10562 39536
rect 10782 40976 10838 41032
rect 10690 40876 10692 40896
rect 10692 40876 10744 40896
rect 10744 40876 10746 40896
rect 10690 40840 10746 40876
rect 10966 40024 11022 40080
rect 10874 38156 10876 38176
rect 10876 38156 10928 38176
rect 10928 38156 10930 38176
rect 10874 38120 10930 38156
rect 11058 37204 11060 37224
rect 11060 37204 11112 37224
rect 11112 37204 11114 37224
rect 11058 37168 11114 37204
rect 10690 33088 10746 33144
rect 10874 28736 10930 28792
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 12070 41112 12126 41168
rect 12254 40568 12310 40624
rect 12622 41112 12678 41168
rect 12162 40160 12218 40216
rect 12346 40180 12402 40216
rect 12346 40160 12348 40180
rect 12348 40160 12400 40180
rect 12400 40160 12402 40180
rect 11886 38836 11888 38856
rect 11888 38836 11940 38856
rect 11940 38836 11942 38856
rect 11886 38800 11942 38836
rect 12070 38936 12126 38992
rect 12254 39888 12310 39944
rect 11242 29008 11298 29064
rect 12254 36760 12310 36816
rect 12438 39924 12440 39944
rect 12440 39924 12492 39944
rect 12492 39924 12494 39944
rect 12438 39888 12494 39924
rect 12530 39208 12586 39264
rect 12530 38664 12586 38720
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 12990 40588 13046 40624
rect 12990 40568 12992 40588
rect 12992 40568 13044 40588
rect 13044 40568 13046 40588
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12898 39480 12954 39536
rect 13082 39480 13138 39536
rect 12990 39072 13046 39128
rect 14370 41792 14426 41848
rect 13542 39208 13598 39264
rect 13634 39072 13690 39128
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 12990 37748 12992 37768
rect 12992 37748 13044 37768
rect 13044 37748 13046 37768
rect 12990 37712 13046 37748
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 13818 37984 13874 38040
rect 12622 33904 12678 33960
rect 13358 35028 13360 35048
rect 13360 35028 13412 35048
rect 13412 35028 13414 35048
rect 13358 34992 13414 35028
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12622 29008 12678 29064
rect 14186 38800 14242 38856
rect 13266 28952 13322 29008
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 13910 29144 13966 29200
rect 13818 28952 13874 29008
rect 13818 28736 13874 28792
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 14002 28908 14004 28928
rect 14004 28908 14056 28928
rect 14056 28908 14058 28928
rect 14002 28872 14058 28908
rect 14738 41676 14794 41712
rect 14738 41656 14740 41676
rect 14740 41656 14792 41676
rect 14792 41656 14794 41676
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 15934 45464 15990 45520
rect 14922 40976 14978 41032
rect 14646 33924 14702 33960
rect 14646 33904 14648 33924
rect 14648 33904 14700 33924
rect 14700 33904 14702 33924
rect 15382 38120 15438 38176
rect 15934 38120 15990 38176
rect 15474 32544 15530 32600
rect 16946 37984 17002 38040
rect 17222 38120 17278 38176
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 17866 48068 17922 48104
rect 17866 48048 17868 48068
rect 17868 48048 17920 48068
rect 17920 48048 17922 48068
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 18418 48048 18474 48104
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17498 41792 17554 41848
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 18234 41520 18290 41576
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 18234 38956 18290 38992
rect 18234 38936 18236 38956
rect 18236 38936 18288 38956
rect 18288 38936 18290 38956
rect 17774 38120 17830 38176
rect 20442 45464 20498 45520
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 18694 42628 18750 42664
rect 18694 42608 18696 42628
rect 18696 42608 18748 42628
rect 18748 42608 18750 42628
rect 18510 41520 18566 41576
rect 18510 40432 18566 40488
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 18418 37712 18474 37768
rect 17774 37188 17830 37224
rect 17774 37168 17776 37188
rect 17776 37168 17828 37188
rect 17828 37168 17830 37188
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 17406 33924 17462 33960
rect 17406 33904 17408 33924
rect 17408 33904 17460 33924
rect 17460 33904 17462 33924
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 17866 33904 17922 33960
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 18786 41928 18842 41984
rect 18694 39480 18750 39536
rect 18878 40024 18934 40080
rect 18786 37188 18842 37224
rect 18786 37168 18788 37188
rect 18788 37168 18840 37188
rect 18840 37168 18842 37188
rect 19614 41384 19670 41440
rect 20718 42744 20774 42800
rect 20994 41656 21050 41712
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 19430 38664 19486 38720
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 21362 38664 21418 38720
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 23754 45464 23810 45520
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 23754 41420 23756 41440
rect 23756 41420 23808 41440
rect 23808 41420 23810 41440
rect 23754 41384 23810 41420
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 23478 37848 23534 37904
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 27956 54426 28012 54428
rect 28036 54426 28092 54428
rect 28116 54426 28172 54428
rect 28196 54426 28252 54428
rect 27956 54374 28002 54426
rect 28002 54374 28012 54426
rect 28036 54374 28066 54426
rect 28066 54374 28078 54426
rect 28078 54374 28092 54426
rect 28116 54374 28130 54426
rect 28130 54374 28142 54426
rect 28142 54374 28172 54426
rect 28196 54374 28206 54426
rect 28206 54374 28252 54426
rect 27956 54372 28012 54374
rect 28036 54372 28092 54374
rect 28116 54372 28172 54374
rect 28196 54372 28252 54374
rect 27956 53338 28012 53340
rect 28036 53338 28092 53340
rect 28116 53338 28172 53340
rect 28196 53338 28252 53340
rect 27956 53286 28002 53338
rect 28002 53286 28012 53338
rect 28036 53286 28066 53338
rect 28066 53286 28078 53338
rect 28078 53286 28092 53338
rect 28116 53286 28130 53338
rect 28130 53286 28142 53338
rect 28142 53286 28172 53338
rect 28196 53286 28206 53338
rect 28206 53286 28252 53338
rect 27956 53284 28012 53286
rect 28036 53284 28092 53286
rect 28116 53284 28172 53286
rect 28196 53284 28252 53286
rect 27956 52250 28012 52252
rect 28036 52250 28092 52252
rect 28116 52250 28172 52252
rect 28196 52250 28252 52252
rect 27956 52198 28002 52250
rect 28002 52198 28012 52250
rect 28036 52198 28066 52250
rect 28066 52198 28078 52250
rect 28078 52198 28092 52250
rect 28116 52198 28130 52250
rect 28130 52198 28142 52250
rect 28142 52198 28172 52250
rect 28196 52198 28206 52250
rect 28206 52198 28252 52250
rect 27956 52196 28012 52198
rect 28036 52196 28092 52198
rect 28116 52196 28172 52198
rect 28196 52196 28252 52198
rect 27956 51162 28012 51164
rect 28036 51162 28092 51164
rect 28116 51162 28172 51164
rect 28196 51162 28252 51164
rect 27956 51110 28002 51162
rect 28002 51110 28012 51162
rect 28036 51110 28066 51162
rect 28066 51110 28078 51162
rect 28078 51110 28092 51162
rect 28116 51110 28130 51162
rect 28130 51110 28142 51162
rect 28142 51110 28172 51162
rect 28196 51110 28206 51162
rect 28206 51110 28252 51162
rect 27956 51108 28012 51110
rect 28036 51108 28092 51110
rect 28116 51108 28172 51110
rect 28196 51108 28252 51110
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 27956 50074 28012 50076
rect 28036 50074 28092 50076
rect 28116 50074 28172 50076
rect 28196 50074 28252 50076
rect 27956 50022 28002 50074
rect 28002 50022 28012 50074
rect 28036 50022 28066 50074
rect 28066 50022 28078 50074
rect 28078 50022 28092 50074
rect 28116 50022 28130 50074
rect 28130 50022 28142 50074
rect 28142 50022 28172 50074
rect 28196 50022 28206 50074
rect 28206 50022 28252 50074
rect 27956 50020 28012 50022
rect 28036 50020 28092 50022
rect 28116 50020 28172 50022
rect 28196 50020 28252 50022
rect 27956 48986 28012 48988
rect 28036 48986 28092 48988
rect 28116 48986 28172 48988
rect 28196 48986 28252 48988
rect 27956 48934 28002 48986
rect 28002 48934 28012 48986
rect 28036 48934 28066 48986
rect 28066 48934 28078 48986
rect 28078 48934 28092 48986
rect 28116 48934 28130 48986
rect 28130 48934 28142 48986
rect 28142 48934 28172 48986
rect 28196 48934 28206 48986
rect 28206 48934 28252 48986
rect 27956 48932 28012 48934
rect 28036 48932 28092 48934
rect 28116 48932 28172 48934
rect 28196 48932 28252 48934
rect 27956 47898 28012 47900
rect 28036 47898 28092 47900
rect 28116 47898 28172 47900
rect 28196 47898 28252 47900
rect 27956 47846 28002 47898
rect 28002 47846 28012 47898
rect 28036 47846 28066 47898
rect 28066 47846 28078 47898
rect 28078 47846 28092 47898
rect 28116 47846 28130 47898
rect 28130 47846 28142 47898
rect 28142 47846 28172 47898
rect 28196 47846 28206 47898
rect 28206 47846 28252 47898
rect 27956 47844 28012 47846
rect 28036 47844 28092 47846
rect 28116 47844 28172 47846
rect 28196 47844 28252 47846
rect 27956 46810 28012 46812
rect 28036 46810 28092 46812
rect 28116 46810 28172 46812
rect 28196 46810 28252 46812
rect 27956 46758 28002 46810
rect 28002 46758 28012 46810
rect 28036 46758 28066 46810
rect 28066 46758 28078 46810
rect 28078 46758 28092 46810
rect 28116 46758 28130 46810
rect 28130 46758 28142 46810
rect 28142 46758 28172 46810
rect 28196 46758 28206 46810
rect 28206 46758 28252 46810
rect 27956 46756 28012 46758
rect 28036 46756 28092 46758
rect 28116 46756 28172 46758
rect 28196 46756 28252 46758
rect 27956 45722 28012 45724
rect 28036 45722 28092 45724
rect 28116 45722 28172 45724
rect 28196 45722 28252 45724
rect 27956 45670 28002 45722
rect 28002 45670 28012 45722
rect 28036 45670 28066 45722
rect 28066 45670 28078 45722
rect 28078 45670 28092 45722
rect 28116 45670 28130 45722
rect 28130 45670 28142 45722
rect 28142 45670 28172 45722
rect 28196 45670 28206 45722
rect 28206 45670 28252 45722
rect 27956 45668 28012 45670
rect 28036 45668 28092 45670
rect 28116 45668 28172 45670
rect 28196 45668 28252 45670
rect 27956 44634 28012 44636
rect 28036 44634 28092 44636
rect 28116 44634 28172 44636
rect 28196 44634 28252 44636
rect 27956 44582 28002 44634
rect 28002 44582 28012 44634
rect 28036 44582 28066 44634
rect 28066 44582 28078 44634
rect 28078 44582 28092 44634
rect 28116 44582 28130 44634
rect 28130 44582 28142 44634
rect 28142 44582 28172 44634
rect 28196 44582 28206 44634
rect 28206 44582 28252 44634
rect 27956 44580 28012 44582
rect 28036 44580 28092 44582
rect 28116 44580 28172 44582
rect 28196 44580 28252 44582
rect 27956 43546 28012 43548
rect 28036 43546 28092 43548
rect 28116 43546 28172 43548
rect 28196 43546 28252 43548
rect 27956 43494 28002 43546
rect 28002 43494 28012 43546
rect 28036 43494 28066 43546
rect 28066 43494 28078 43546
rect 28078 43494 28092 43546
rect 28116 43494 28130 43546
rect 28130 43494 28142 43546
rect 28142 43494 28172 43546
rect 28196 43494 28206 43546
rect 28206 43494 28252 43546
rect 27956 43492 28012 43494
rect 28036 43492 28092 43494
rect 28116 43492 28172 43494
rect 28196 43492 28252 43494
rect 35070 54032 35126 54088
rect 32956 53882 33012 53884
rect 33036 53882 33092 53884
rect 33116 53882 33172 53884
rect 33196 53882 33252 53884
rect 32956 53830 33002 53882
rect 33002 53830 33012 53882
rect 33036 53830 33066 53882
rect 33066 53830 33078 53882
rect 33078 53830 33092 53882
rect 33116 53830 33130 53882
rect 33130 53830 33142 53882
rect 33142 53830 33172 53882
rect 33196 53830 33206 53882
rect 33206 53830 33252 53882
rect 32956 53828 33012 53830
rect 33036 53828 33092 53830
rect 33116 53828 33172 53830
rect 33196 53828 33252 53830
rect 32956 52794 33012 52796
rect 33036 52794 33092 52796
rect 33116 52794 33172 52796
rect 33196 52794 33252 52796
rect 32956 52742 33002 52794
rect 33002 52742 33012 52794
rect 33036 52742 33066 52794
rect 33066 52742 33078 52794
rect 33078 52742 33092 52794
rect 33116 52742 33130 52794
rect 33130 52742 33142 52794
rect 33142 52742 33172 52794
rect 33196 52742 33206 52794
rect 33206 52742 33252 52794
rect 32956 52740 33012 52742
rect 33036 52740 33092 52742
rect 33116 52740 33172 52742
rect 33196 52740 33252 52742
rect 32956 51706 33012 51708
rect 33036 51706 33092 51708
rect 33116 51706 33172 51708
rect 33196 51706 33252 51708
rect 32956 51654 33002 51706
rect 33002 51654 33012 51706
rect 33036 51654 33066 51706
rect 33066 51654 33078 51706
rect 33078 51654 33092 51706
rect 33116 51654 33130 51706
rect 33130 51654 33142 51706
rect 33142 51654 33172 51706
rect 33196 51654 33206 51706
rect 33206 51654 33252 51706
rect 32956 51652 33012 51654
rect 33036 51652 33092 51654
rect 33116 51652 33172 51654
rect 33196 51652 33252 51654
rect 32956 50618 33012 50620
rect 33036 50618 33092 50620
rect 33116 50618 33172 50620
rect 33196 50618 33252 50620
rect 32956 50566 33002 50618
rect 33002 50566 33012 50618
rect 33036 50566 33066 50618
rect 33066 50566 33078 50618
rect 33078 50566 33092 50618
rect 33116 50566 33130 50618
rect 33130 50566 33142 50618
rect 33142 50566 33172 50618
rect 33196 50566 33206 50618
rect 33206 50566 33252 50618
rect 32956 50564 33012 50566
rect 33036 50564 33092 50566
rect 33116 50564 33172 50566
rect 33196 50564 33252 50566
rect 32956 49530 33012 49532
rect 33036 49530 33092 49532
rect 33116 49530 33172 49532
rect 33196 49530 33252 49532
rect 32956 49478 33002 49530
rect 33002 49478 33012 49530
rect 33036 49478 33066 49530
rect 33066 49478 33078 49530
rect 33078 49478 33092 49530
rect 33116 49478 33130 49530
rect 33130 49478 33142 49530
rect 33142 49478 33172 49530
rect 33196 49478 33206 49530
rect 33206 49478 33252 49530
rect 32956 49476 33012 49478
rect 33036 49476 33092 49478
rect 33116 49476 33172 49478
rect 33196 49476 33252 49478
rect 29826 43288 29882 43344
rect 27956 42458 28012 42460
rect 28036 42458 28092 42460
rect 28116 42458 28172 42460
rect 28196 42458 28252 42460
rect 27956 42406 28002 42458
rect 28002 42406 28012 42458
rect 28036 42406 28066 42458
rect 28066 42406 28078 42458
rect 28078 42406 28092 42458
rect 28116 42406 28130 42458
rect 28130 42406 28142 42458
rect 28142 42406 28172 42458
rect 28196 42406 28206 42458
rect 28206 42406 28252 42458
rect 27956 42404 28012 42406
rect 28036 42404 28092 42406
rect 28116 42404 28172 42406
rect 28196 42404 28252 42406
rect 27956 41370 28012 41372
rect 28036 41370 28092 41372
rect 28116 41370 28172 41372
rect 28196 41370 28252 41372
rect 27956 41318 28002 41370
rect 28002 41318 28012 41370
rect 28036 41318 28066 41370
rect 28066 41318 28078 41370
rect 28078 41318 28092 41370
rect 28116 41318 28130 41370
rect 28130 41318 28142 41370
rect 28142 41318 28172 41370
rect 28196 41318 28206 41370
rect 28206 41318 28252 41370
rect 27956 41316 28012 41318
rect 28036 41316 28092 41318
rect 28116 41316 28172 41318
rect 28196 41316 28252 41318
rect 27956 40282 28012 40284
rect 28036 40282 28092 40284
rect 28116 40282 28172 40284
rect 28196 40282 28252 40284
rect 27956 40230 28002 40282
rect 28002 40230 28012 40282
rect 28036 40230 28066 40282
rect 28066 40230 28078 40282
rect 28078 40230 28092 40282
rect 28116 40230 28130 40282
rect 28130 40230 28142 40282
rect 28142 40230 28172 40282
rect 28196 40230 28206 40282
rect 28206 40230 28252 40282
rect 27956 40228 28012 40230
rect 28036 40228 28092 40230
rect 28116 40228 28172 40230
rect 28196 40228 28252 40230
rect 27956 39194 28012 39196
rect 28036 39194 28092 39196
rect 28116 39194 28172 39196
rect 28196 39194 28252 39196
rect 27956 39142 28002 39194
rect 28002 39142 28012 39194
rect 28036 39142 28066 39194
rect 28066 39142 28078 39194
rect 28078 39142 28092 39194
rect 28116 39142 28130 39194
rect 28130 39142 28142 39194
rect 28142 39142 28172 39194
rect 28196 39142 28206 39194
rect 28206 39142 28252 39194
rect 27956 39140 28012 39142
rect 28036 39140 28092 39142
rect 28116 39140 28172 39142
rect 28196 39140 28252 39142
rect 27956 38106 28012 38108
rect 28036 38106 28092 38108
rect 28116 38106 28172 38108
rect 28196 38106 28252 38108
rect 27956 38054 28002 38106
rect 28002 38054 28012 38106
rect 28036 38054 28066 38106
rect 28066 38054 28078 38106
rect 28078 38054 28092 38106
rect 28116 38054 28130 38106
rect 28130 38054 28142 38106
rect 28142 38054 28172 38106
rect 28196 38054 28206 38106
rect 28206 38054 28252 38106
rect 27956 38052 28012 38054
rect 28036 38052 28092 38054
rect 28116 38052 28172 38054
rect 28196 38052 28252 38054
rect 27956 37018 28012 37020
rect 28036 37018 28092 37020
rect 28116 37018 28172 37020
rect 28196 37018 28252 37020
rect 27956 36966 28002 37018
rect 28002 36966 28012 37018
rect 28036 36966 28066 37018
rect 28066 36966 28078 37018
rect 28078 36966 28092 37018
rect 28116 36966 28130 37018
rect 28130 36966 28142 37018
rect 28142 36966 28172 37018
rect 28196 36966 28206 37018
rect 28206 36966 28252 37018
rect 27956 36964 28012 36966
rect 28036 36964 28092 36966
rect 28116 36964 28172 36966
rect 28196 36964 28252 36966
rect 27956 35930 28012 35932
rect 28036 35930 28092 35932
rect 28116 35930 28172 35932
rect 28196 35930 28252 35932
rect 27956 35878 28002 35930
rect 28002 35878 28012 35930
rect 28036 35878 28066 35930
rect 28066 35878 28078 35930
rect 28078 35878 28092 35930
rect 28116 35878 28130 35930
rect 28130 35878 28142 35930
rect 28142 35878 28172 35930
rect 28196 35878 28206 35930
rect 28206 35878 28252 35930
rect 27956 35876 28012 35878
rect 28036 35876 28092 35878
rect 28116 35876 28172 35878
rect 28196 35876 28252 35878
rect 27956 34842 28012 34844
rect 28036 34842 28092 34844
rect 28116 34842 28172 34844
rect 28196 34842 28252 34844
rect 27956 34790 28002 34842
rect 28002 34790 28012 34842
rect 28036 34790 28066 34842
rect 28066 34790 28078 34842
rect 28078 34790 28092 34842
rect 28116 34790 28130 34842
rect 28130 34790 28142 34842
rect 28142 34790 28172 34842
rect 28196 34790 28206 34842
rect 28206 34790 28252 34842
rect 27956 34788 28012 34790
rect 28036 34788 28092 34790
rect 28116 34788 28172 34790
rect 28196 34788 28252 34790
rect 27956 33754 28012 33756
rect 28036 33754 28092 33756
rect 28116 33754 28172 33756
rect 28196 33754 28252 33756
rect 27956 33702 28002 33754
rect 28002 33702 28012 33754
rect 28036 33702 28066 33754
rect 28066 33702 28078 33754
rect 28078 33702 28092 33754
rect 28116 33702 28130 33754
rect 28130 33702 28142 33754
rect 28142 33702 28172 33754
rect 28196 33702 28206 33754
rect 28206 33702 28252 33754
rect 27956 33700 28012 33702
rect 28036 33700 28092 33702
rect 28116 33700 28172 33702
rect 28196 33700 28252 33702
rect 27956 32666 28012 32668
rect 28036 32666 28092 32668
rect 28116 32666 28172 32668
rect 28196 32666 28252 32668
rect 27956 32614 28002 32666
rect 28002 32614 28012 32666
rect 28036 32614 28066 32666
rect 28066 32614 28078 32666
rect 28078 32614 28092 32666
rect 28116 32614 28130 32666
rect 28130 32614 28142 32666
rect 28142 32614 28172 32666
rect 28196 32614 28206 32666
rect 28206 32614 28252 32666
rect 27956 32612 28012 32614
rect 28036 32612 28092 32614
rect 28116 32612 28172 32614
rect 28196 32612 28252 32614
rect 27956 31578 28012 31580
rect 28036 31578 28092 31580
rect 28116 31578 28172 31580
rect 28196 31578 28252 31580
rect 27956 31526 28002 31578
rect 28002 31526 28012 31578
rect 28036 31526 28066 31578
rect 28066 31526 28078 31578
rect 28078 31526 28092 31578
rect 28116 31526 28130 31578
rect 28130 31526 28142 31578
rect 28142 31526 28172 31578
rect 28196 31526 28206 31578
rect 28206 31526 28252 31578
rect 27956 31524 28012 31526
rect 28036 31524 28092 31526
rect 28116 31524 28172 31526
rect 28196 31524 28252 31526
rect 27956 30490 28012 30492
rect 28036 30490 28092 30492
rect 28116 30490 28172 30492
rect 28196 30490 28252 30492
rect 27956 30438 28002 30490
rect 28002 30438 28012 30490
rect 28036 30438 28066 30490
rect 28066 30438 28078 30490
rect 28078 30438 28092 30490
rect 28116 30438 28130 30490
rect 28130 30438 28142 30490
rect 28142 30438 28172 30490
rect 28196 30438 28206 30490
rect 28206 30438 28252 30490
rect 27956 30436 28012 30438
rect 28036 30436 28092 30438
rect 28116 30436 28172 30438
rect 28196 30436 28252 30438
rect 27956 29402 28012 29404
rect 28036 29402 28092 29404
rect 28116 29402 28172 29404
rect 28196 29402 28252 29404
rect 27956 29350 28002 29402
rect 28002 29350 28012 29402
rect 28036 29350 28066 29402
rect 28066 29350 28078 29402
rect 28078 29350 28092 29402
rect 28116 29350 28130 29402
rect 28130 29350 28142 29402
rect 28142 29350 28172 29402
rect 28196 29350 28206 29402
rect 28206 29350 28252 29402
rect 27956 29348 28012 29350
rect 28036 29348 28092 29350
rect 28116 29348 28172 29350
rect 28196 29348 28252 29350
rect 27956 28314 28012 28316
rect 28036 28314 28092 28316
rect 28116 28314 28172 28316
rect 28196 28314 28252 28316
rect 27956 28262 28002 28314
rect 28002 28262 28012 28314
rect 28036 28262 28066 28314
rect 28066 28262 28078 28314
rect 28078 28262 28092 28314
rect 28116 28262 28130 28314
rect 28130 28262 28142 28314
rect 28142 28262 28172 28314
rect 28196 28262 28206 28314
rect 28206 28262 28252 28314
rect 27956 28260 28012 28262
rect 28036 28260 28092 28262
rect 28116 28260 28172 28262
rect 28196 28260 28252 28262
rect 27956 27226 28012 27228
rect 28036 27226 28092 27228
rect 28116 27226 28172 27228
rect 28196 27226 28252 27228
rect 27956 27174 28002 27226
rect 28002 27174 28012 27226
rect 28036 27174 28066 27226
rect 28066 27174 28078 27226
rect 28078 27174 28092 27226
rect 28116 27174 28130 27226
rect 28130 27174 28142 27226
rect 28142 27174 28172 27226
rect 28196 27174 28206 27226
rect 28206 27174 28252 27226
rect 27956 27172 28012 27174
rect 28036 27172 28092 27174
rect 28116 27172 28172 27174
rect 28196 27172 28252 27174
rect 27956 26138 28012 26140
rect 28036 26138 28092 26140
rect 28116 26138 28172 26140
rect 28196 26138 28252 26140
rect 27956 26086 28002 26138
rect 28002 26086 28012 26138
rect 28036 26086 28066 26138
rect 28066 26086 28078 26138
rect 28078 26086 28092 26138
rect 28116 26086 28130 26138
rect 28130 26086 28142 26138
rect 28142 26086 28172 26138
rect 28196 26086 28206 26138
rect 28206 26086 28252 26138
rect 27956 26084 28012 26086
rect 28036 26084 28092 26086
rect 28116 26084 28172 26086
rect 28196 26084 28252 26086
rect 27956 25050 28012 25052
rect 28036 25050 28092 25052
rect 28116 25050 28172 25052
rect 28196 25050 28252 25052
rect 27956 24998 28002 25050
rect 28002 24998 28012 25050
rect 28036 24998 28066 25050
rect 28066 24998 28078 25050
rect 28078 24998 28092 25050
rect 28116 24998 28130 25050
rect 28130 24998 28142 25050
rect 28142 24998 28172 25050
rect 28196 24998 28206 25050
rect 28206 24998 28252 25050
rect 27956 24996 28012 24998
rect 28036 24996 28092 24998
rect 28116 24996 28172 24998
rect 28196 24996 28252 24998
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 32956 48442 33012 48444
rect 33036 48442 33092 48444
rect 33116 48442 33172 48444
rect 33196 48442 33252 48444
rect 32956 48390 33002 48442
rect 33002 48390 33012 48442
rect 33036 48390 33066 48442
rect 33066 48390 33078 48442
rect 33078 48390 33092 48442
rect 33116 48390 33130 48442
rect 33130 48390 33142 48442
rect 33142 48390 33172 48442
rect 33196 48390 33206 48442
rect 33206 48390 33252 48442
rect 32956 48388 33012 48390
rect 33036 48388 33092 48390
rect 33116 48388 33172 48390
rect 33196 48388 33252 48390
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 32956 47354 33012 47356
rect 33036 47354 33092 47356
rect 33116 47354 33172 47356
rect 33196 47354 33252 47356
rect 32956 47302 33002 47354
rect 33002 47302 33012 47354
rect 33036 47302 33066 47354
rect 33066 47302 33078 47354
rect 33078 47302 33092 47354
rect 33116 47302 33130 47354
rect 33130 47302 33142 47354
rect 33142 47302 33172 47354
rect 33196 47302 33206 47354
rect 33206 47302 33252 47354
rect 32956 47300 33012 47302
rect 33036 47300 33092 47302
rect 33116 47300 33172 47302
rect 33196 47300 33252 47302
rect 32956 46266 33012 46268
rect 33036 46266 33092 46268
rect 33116 46266 33172 46268
rect 33196 46266 33252 46268
rect 32956 46214 33002 46266
rect 33002 46214 33012 46266
rect 33036 46214 33066 46266
rect 33066 46214 33078 46266
rect 33078 46214 33092 46266
rect 33116 46214 33130 46266
rect 33130 46214 33142 46266
rect 33142 46214 33172 46266
rect 33196 46214 33206 46266
rect 33206 46214 33252 46266
rect 32956 46212 33012 46214
rect 33036 46212 33092 46214
rect 33116 46212 33172 46214
rect 33196 46212 33252 46214
rect 32956 45178 33012 45180
rect 33036 45178 33092 45180
rect 33116 45178 33172 45180
rect 33196 45178 33252 45180
rect 32956 45126 33002 45178
rect 33002 45126 33012 45178
rect 33036 45126 33066 45178
rect 33066 45126 33078 45178
rect 33078 45126 33092 45178
rect 33116 45126 33130 45178
rect 33130 45126 33142 45178
rect 33142 45126 33172 45178
rect 33196 45126 33206 45178
rect 33206 45126 33252 45178
rect 32956 45124 33012 45126
rect 33036 45124 33092 45126
rect 33116 45124 33172 45126
rect 33196 45124 33252 45126
rect 32956 44090 33012 44092
rect 33036 44090 33092 44092
rect 33116 44090 33172 44092
rect 33196 44090 33252 44092
rect 32956 44038 33002 44090
rect 33002 44038 33012 44090
rect 33036 44038 33066 44090
rect 33066 44038 33078 44090
rect 33078 44038 33092 44090
rect 33116 44038 33130 44090
rect 33130 44038 33142 44090
rect 33142 44038 33172 44090
rect 33196 44038 33206 44090
rect 33206 44038 33252 44090
rect 32956 44036 33012 44038
rect 33036 44036 33092 44038
rect 33116 44036 33172 44038
rect 33196 44036 33252 44038
rect 32956 43002 33012 43004
rect 33036 43002 33092 43004
rect 33116 43002 33172 43004
rect 33196 43002 33252 43004
rect 32956 42950 33002 43002
rect 33002 42950 33012 43002
rect 33036 42950 33066 43002
rect 33066 42950 33078 43002
rect 33078 42950 33092 43002
rect 33116 42950 33130 43002
rect 33130 42950 33142 43002
rect 33142 42950 33172 43002
rect 33196 42950 33206 43002
rect 33206 42950 33252 43002
rect 32956 42948 33012 42950
rect 33036 42948 33092 42950
rect 33116 42948 33172 42950
rect 33196 42948 33252 42950
rect 32956 41914 33012 41916
rect 33036 41914 33092 41916
rect 33116 41914 33172 41916
rect 33196 41914 33252 41916
rect 32956 41862 33002 41914
rect 33002 41862 33012 41914
rect 33036 41862 33066 41914
rect 33066 41862 33078 41914
rect 33078 41862 33092 41914
rect 33116 41862 33130 41914
rect 33130 41862 33142 41914
rect 33142 41862 33172 41914
rect 33196 41862 33206 41914
rect 33206 41862 33252 41914
rect 32956 41860 33012 41862
rect 33036 41860 33092 41862
rect 33116 41860 33172 41862
rect 33196 41860 33252 41862
rect 32956 40826 33012 40828
rect 33036 40826 33092 40828
rect 33116 40826 33172 40828
rect 33196 40826 33252 40828
rect 32956 40774 33002 40826
rect 33002 40774 33012 40826
rect 33036 40774 33066 40826
rect 33066 40774 33078 40826
rect 33078 40774 33092 40826
rect 33116 40774 33130 40826
rect 33130 40774 33142 40826
rect 33142 40774 33172 40826
rect 33196 40774 33206 40826
rect 33206 40774 33252 40826
rect 32956 40772 33012 40774
rect 33036 40772 33092 40774
rect 33116 40772 33172 40774
rect 33196 40772 33252 40774
rect 32956 39738 33012 39740
rect 33036 39738 33092 39740
rect 33116 39738 33172 39740
rect 33196 39738 33252 39740
rect 32956 39686 33002 39738
rect 33002 39686 33012 39738
rect 33036 39686 33066 39738
rect 33066 39686 33078 39738
rect 33078 39686 33092 39738
rect 33116 39686 33130 39738
rect 33130 39686 33142 39738
rect 33142 39686 33172 39738
rect 33196 39686 33206 39738
rect 33206 39686 33252 39738
rect 32956 39684 33012 39686
rect 33036 39684 33092 39686
rect 33116 39684 33172 39686
rect 33196 39684 33252 39686
rect 32956 38650 33012 38652
rect 33036 38650 33092 38652
rect 33116 38650 33172 38652
rect 33196 38650 33252 38652
rect 32956 38598 33002 38650
rect 33002 38598 33012 38650
rect 33036 38598 33066 38650
rect 33066 38598 33078 38650
rect 33078 38598 33092 38650
rect 33116 38598 33130 38650
rect 33130 38598 33142 38650
rect 33142 38598 33172 38650
rect 33196 38598 33206 38650
rect 33206 38598 33252 38650
rect 32956 38596 33012 38598
rect 33036 38596 33092 38598
rect 33116 38596 33172 38598
rect 33196 38596 33252 38598
rect 32956 37562 33012 37564
rect 33036 37562 33092 37564
rect 33116 37562 33172 37564
rect 33196 37562 33252 37564
rect 32956 37510 33002 37562
rect 33002 37510 33012 37562
rect 33036 37510 33066 37562
rect 33066 37510 33078 37562
rect 33078 37510 33092 37562
rect 33116 37510 33130 37562
rect 33130 37510 33142 37562
rect 33142 37510 33172 37562
rect 33196 37510 33206 37562
rect 33206 37510 33252 37562
rect 32956 37508 33012 37510
rect 33036 37508 33092 37510
rect 33116 37508 33172 37510
rect 33196 37508 33252 37510
rect 32956 36474 33012 36476
rect 33036 36474 33092 36476
rect 33116 36474 33172 36476
rect 33196 36474 33252 36476
rect 32956 36422 33002 36474
rect 33002 36422 33012 36474
rect 33036 36422 33066 36474
rect 33066 36422 33078 36474
rect 33078 36422 33092 36474
rect 33116 36422 33130 36474
rect 33130 36422 33142 36474
rect 33142 36422 33172 36474
rect 33196 36422 33206 36474
rect 33206 36422 33252 36474
rect 32956 36420 33012 36422
rect 33036 36420 33092 36422
rect 33116 36420 33172 36422
rect 33196 36420 33252 36422
rect 32956 35386 33012 35388
rect 33036 35386 33092 35388
rect 33116 35386 33172 35388
rect 33196 35386 33252 35388
rect 32956 35334 33002 35386
rect 33002 35334 33012 35386
rect 33036 35334 33066 35386
rect 33066 35334 33078 35386
rect 33078 35334 33092 35386
rect 33116 35334 33130 35386
rect 33130 35334 33142 35386
rect 33142 35334 33172 35386
rect 33196 35334 33206 35386
rect 33206 35334 33252 35386
rect 32956 35332 33012 35334
rect 33036 35332 33092 35334
rect 33116 35332 33172 35334
rect 33196 35332 33252 35334
rect 32956 34298 33012 34300
rect 33036 34298 33092 34300
rect 33116 34298 33172 34300
rect 33196 34298 33252 34300
rect 32956 34246 33002 34298
rect 33002 34246 33012 34298
rect 33036 34246 33066 34298
rect 33066 34246 33078 34298
rect 33078 34246 33092 34298
rect 33116 34246 33130 34298
rect 33130 34246 33142 34298
rect 33142 34246 33172 34298
rect 33196 34246 33206 34298
rect 33206 34246 33252 34298
rect 32956 34244 33012 34246
rect 33036 34244 33092 34246
rect 33116 34244 33172 34246
rect 33196 34244 33252 34246
rect 32956 33210 33012 33212
rect 33036 33210 33092 33212
rect 33116 33210 33172 33212
rect 33196 33210 33252 33212
rect 32956 33158 33002 33210
rect 33002 33158 33012 33210
rect 33036 33158 33066 33210
rect 33066 33158 33078 33210
rect 33078 33158 33092 33210
rect 33116 33158 33130 33210
rect 33130 33158 33142 33210
rect 33142 33158 33172 33210
rect 33196 33158 33206 33210
rect 33206 33158 33252 33210
rect 32956 33156 33012 33158
rect 33036 33156 33092 33158
rect 33116 33156 33172 33158
rect 33196 33156 33252 33158
rect 32956 32122 33012 32124
rect 33036 32122 33092 32124
rect 33116 32122 33172 32124
rect 33196 32122 33252 32124
rect 32956 32070 33002 32122
rect 33002 32070 33012 32122
rect 33036 32070 33066 32122
rect 33066 32070 33078 32122
rect 33078 32070 33092 32122
rect 33116 32070 33130 32122
rect 33130 32070 33142 32122
rect 33142 32070 33172 32122
rect 33196 32070 33206 32122
rect 33206 32070 33252 32122
rect 32956 32068 33012 32070
rect 33036 32068 33092 32070
rect 33116 32068 33172 32070
rect 33196 32068 33252 32070
rect 32956 31034 33012 31036
rect 33036 31034 33092 31036
rect 33116 31034 33172 31036
rect 33196 31034 33252 31036
rect 32956 30982 33002 31034
rect 33002 30982 33012 31034
rect 33036 30982 33066 31034
rect 33066 30982 33078 31034
rect 33078 30982 33092 31034
rect 33116 30982 33130 31034
rect 33130 30982 33142 31034
rect 33142 30982 33172 31034
rect 33196 30982 33206 31034
rect 33206 30982 33252 31034
rect 32956 30980 33012 30982
rect 33036 30980 33092 30982
rect 33116 30980 33172 30982
rect 33196 30980 33252 30982
rect 32956 29946 33012 29948
rect 33036 29946 33092 29948
rect 33116 29946 33172 29948
rect 33196 29946 33252 29948
rect 32956 29894 33002 29946
rect 33002 29894 33012 29946
rect 33036 29894 33066 29946
rect 33066 29894 33078 29946
rect 33078 29894 33092 29946
rect 33116 29894 33130 29946
rect 33130 29894 33142 29946
rect 33142 29894 33172 29946
rect 33196 29894 33206 29946
rect 33206 29894 33252 29946
rect 32956 29892 33012 29894
rect 33036 29892 33092 29894
rect 33116 29892 33172 29894
rect 33196 29892 33252 29894
rect 32956 28858 33012 28860
rect 33036 28858 33092 28860
rect 33116 28858 33172 28860
rect 33196 28858 33252 28860
rect 32956 28806 33002 28858
rect 33002 28806 33012 28858
rect 33036 28806 33066 28858
rect 33066 28806 33078 28858
rect 33078 28806 33092 28858
rect 33116 28806 33130 28858
rect 33130 28806 33142 28858
rect 33142 28806 33172 28858
rect 33196 28806 33206 28858
rect 33206 28806 33252 28858
rect 32956 28804 33012 28806
rect 33036 28804 33092 28806
rect 33116 28804 33172 28806
rect 33196 28804 33252 28806
rect 32956 27770 33012 27772
rect 33036 27770 33092 27772
rect 33116 27770 33172 27772
rect 33196 27770 33252 27772
rect 32956 27718 33002 27770
rect 33002 27718 33012 27770
rect 33036 27718 33066 27770
rect 33066 27718 33078 27770
rect 33078 27718 33092 27770
rect 33116 27718 33130 27770
rect 33130 27718 33142 27770
rect 33142 27718 33172 27770
rect 33196 27718 33206 27770
rect 33206 27718 33252 27770
rect 32956 27716 33012 27718
rect 33036 27716 33092 27718
rect 33116 27716 33172 27718
rect 33196 27716 33252 27718
rect 32956 26682 33012 26684
rect 33036 26682 33092 26684
rect 33116 26682 33172 26684
rect 33196 26682 33252 26684
rect 32956 26630 33002 26682
rect 33002 26630 33012 26682
rect 33036 26630 33066 26682
rect 33066 26630 33078 26682
rect 33078 26630 33092 26682
rect 33116 26630 33130 26682
rect 33130 26630 33142 26682
rect 33142 26630 33172 26682
rect 33196 26630 33206 26682
rect 33206 26630 33252 26682
rect 32956 26628 33012 26630
rect 33036 26628 33092 26630
rect 33116 26628 33172 26630
rect 33196 26628 33252 26630
rect 32956 25594 33012 25596
rect 33036 25594 33092 25596
rect 33116 25594 33172 25596
rect 33196 25594 33252 25596
rect 32956 25542 33002 25594
rect 33002 25542 33012 25594
rect 33036 25542 33066 25594
rect 33066 25542 33078 25594
rect 33078 25542 33092 25594
rect 33116 25542 33130 25594
rect 33130 25542 33142 25594
rect 33142 25542 33172 25594
rect 33196 25542 33206 25594
rect 33206 25542 33252 25594
rect 32956 25540 33012 25542
rect 33036 25540 33092 25542
rect 33116 25540 33172 25542
rect 33196 25540 33252 25542
rect 37956 54426 38012 54428
rect 38036 54426 38092 54428
rect 38116 54426 38172 54428
rect 38196 54426 38252 54428
rect 37956 54374 38002 54426
rect 38002 54374 38012 54426
rect 38036 54374 38066 54426
rect 38066 54374 38078 54426
rect 38078 54374 38092 54426
rect 38116 54374 38130 54426
rect 38130 54374 38142 54426
rect 38142 54374 38172 54426
rect 38196 54374 38206 54426
rect 38206 54374 38252 54426
rect 37956 54372 38012 54374
rect 38036 54372 38092 54374
rect 38116 54372 38172 54374
rect 38196 54372 38252 54374
rect 34242 41112 34298 41168
rect 37956 53338 38012 53340
rect 38036 53338 38092 53340
rect 38116 53338 38172 53340
rect 38196 53338 38252 53340
rect 37956 53286 38002 53338
rect 38002 53286 38012 53338
rect 38036 53286 38066 53338
rect 38066 53286 38078 53338
rect 38078 53286 38092 53338
rect 38116 53286 38130 53338
rect 38130 53286 38142 53338
rect 38142 53286 38172 53338
rect 38196 53286 38206 53338
rect 38206 53286 38252 53338
rect 37956 53284 38012 53286
rect 38036 53284 38092 53286
rect 38116 53284 38172 53286
rect 38196 53284 38252 53286
rect 37956 52250 38012 52252
rect 38036 52250 38092 52252
rect 38116 52250 38172 52252
rect 38196 52250 38252 52252
rect 37956 52198 38002 52250
rect 38002 52198 38012 52250
rect 38036 52198 38066 52250
rect 38066 52198 38078 52250
rect 38078 52198 38092 52250
rect 38116 52198 38130 52250
rect 38130 52198 38142 52250
rect 38142 52198 38172 52250
rect 38196 52198 38206 52250
rect 38206 52198 38252 52250
rect 37956 52196 38012 52198
rect 38036 52196 38092 52198
rect 38116 52196 38172 52198
rect 38196 52196 38252 52198
rect 37956 51162 38012 51164
rect 38036 51162 38092 51164
rect 38116 51162 38172 51164
rect 38196 51162 38252 51164
rect 37956 51110 38002 51162
rect 38002 51110 38012 51162
rect 38036 51110 38066 51162
rect 38066 51110 38078 51162
rect 38078 51110 38092 51162
rect 38116 51110 38130 51162
rect 38130 51110 38142 51162
rect 38142 51110 38172 51162
rect 38196 51110 38206 51162
rect 38206 51110 38252 51162
rect 37956 51108 38012 51110
rect 38036 51108 38092 51110
rect 38116 51108 38172 51110
rect 38196 51108 38252 51110
rect 37956 50074 38012 50076
rect 38036 50074 38092 50076
rect 38116 50074 38172 50076
rect 38196 50074 38252 50076
rect 37956 50022 38002 50074
rect 38002 50022 38012 50074
rect 38036 50022 38066 50074
rect 38066 50022 38078 50074
rect 38078 50022 38092 50074
rect 38116 50022 38130 50074
rect 38130 50022 38142 50074
rect 38142 50022 38172 50074
rect 38196 50022 38206 50074
rect 38206 50022 38252 50074
rect 37956 50020 38012 50022
rect 38036 50020 38092 50022
rect 38116 50020 38172 50022
rect 38196 50020 38252 50022
rect 37956 48986 38012 48988
rect 38036 48986 38092 48988
rect 38116 48986 38172 48988
rect 38196 48986 38252 48988
rect 37956 48934 38002 48986
rect 38002 48934 38012 48986
rect 38036 48934 38066 48986
rect 38066 48934 38078 48986
rect 38078 48934 38092 48986
rect 38116 48934 38130 48986
rect 38130 48934 38142 48986
rect 38142 48934 38172 48986
rect 38196 48934 38206 48986
rect 38206 48934 38252 48986
rect 37956 48932 38012 48934
rect 38036 48932 38092 48934
rect 38116 48932 38172 48934
rect 38196 48932 38252 48934
rect 37956 47898 38012 47900
rect 38036 47898 38092 47900
rect 38116 47898 38172 47900
rect 38196 47898 38252 47900
rect 37956 47846 38002 47898
rect 38002 47846 38012 47898
rect 38036 47846 38066 47898
rect 38066 47846 38078 47898
rect 38078 47846 38092 47898
rect 38116 47846 38130 47898
rect 38130 47846 38142 47898
rect 38142 47846 38172 47898
rect 38196 47846 38206 47898
rect 38206 47846 38252 47898
rect 37956 47844 38012 47846
rect 38036 47844 38092 47846
rect 38116 47844 38172 47846
rect 38196 47844 38252 47846
rect 37956 46810 38012 46812
rect 38036 46810 38092 46812
rect 38116 46810 38172 46812
rect 38196 46810 38252 46812
rect 37956 46758 38002 46810
rect 38002 46758 38012 46810
rect 38036 46758 38066 46810
rect 38066 46758 38078 46810
rect 38078 46758 38092 46810
rect 38116 46758 38130 46810
rect 38130 46758 38142 46810
rect 38142 46758 38172 46810
rect 38196 46758 38206 46810
rect 38206 46758 38252 46810
rect 37956 46756 38012 46758
rect 38036 46756 38092 46758
rect 38116 46756 38172 46758
rect 38196 46756 38252 46758
rect 37956 45722 38012 45724
rect 38036 45722 38092 45724
rect 38116 45722 38172 45724
rect 38196 45722 38252 45724
rect 37956 45670 38002 45722
rect 38002 45670 38012 45722
rect 38036 45670 38066 45722
rect 38066 45670 38078 45722
rect 38078 45670 38092 45722
rect 38116 45670 38130 45722
rect 38130 45670 38142 45722
rect 38142 45670 38172 45722
rect 38196 45670 38206 45722
rect 38206 45670 38252 45722
rect 37956 45668 38012 45670
rect 38036 45668 38092 45670
rect 38116 45668 38172 45670
rect 38196 45668 38252 45670
rect 37956 44634 38012 44636
rect 38036 44634 38092 44636
rect 38116 44634 38172 44636
rect 38196 44634 38252 44636
rect 37956 44582 38002 44634
rect 38002 44582 38012 44634
rect 38036 44582 38066 44634
rect 38066 44582 38078 44634
rect 38078 44582 38092 44634
rect 38116 44582 38130 44634
rect 38130 44582 38142 44634
rect 38142 44582 38172 44634
rect 38196 44582 38206 44634
rect 38206 44582 38252 44634
rect 37956 44580 38012 44582
rect 38036 44580 38092 44582
rect 38116 44580 38172 44582
rect 38196 44580 38252 44582
rect 37956 43546 38012 43548
rect 38036 43546 38092 43548
rect 38116 43546 38172 43548
rect 38196 43546 38252 43548
rect 37956 43494 38002 43546
rect 38002 43494 38012 43546
rect 38036 43494 38066 43546
rect 38066 43494 38078 43546
rect 38078 43494 38092 43546
rect 38116 43494 38130 43546
rect 38130 43494 38142 43546
rect 38142 43494 38172 43546
rect 38196 43494 38206 43546
rect 38206 43494 38252 43546
rect 37956 43492 38012 43494
rect 38036 43492 38092 43494
rect 38116 43492 38172 43494
rect 38196 43492 38252 43494
rect 37956 42458 38012 42460
rect 38036 42458 38092 42460
rect 38116 42458 38172 42460
rect 38196 42458 38252 42460
rect 37956 42406 38002 42458
rect 38002 42406 38012 42458
rect 38036 42406 38066 42458
rect 38066 42406 38078 42458
rect 38078 42406 38092 42458
rect 38116 42406 38130 42458
rect 38130 42406 38142 42458
rect 38142 42406 38172 42458
rect 38196 42406 38206 42458
rect 38206 42406 38252 42458
rect 37956 42404 38012 42406
rect 38036 42404 38092 42406
rect 38116 42404 38172 42406
rect 38196 42404 38252 42406
rect 37956 41370 38012 41372
rect 38036 41370 38092 41372
rect 38116 41370 38172 41372
rect 38196 41370 38252 41372
rect 37956 41318 38002 41370
rect 38002 41318 38012 41370
rect 38036 41318 38066 41370
rect 38066 41318 38078 41370
rect 38078 41318 38092 41370
rect 38116 41318 38130 41370
rect 38130 41318 38142 41370
rect 38142 41318 38172 41370
rect 38196 41318 38206 41370
rect 38206 41318 38252 41370
rect 37956 41316 38012 41318
rect 38036 41316 38092 41318
rect 38116 41316 38172 41318
rect 38196 41316 38252 41318
rect 37956 40282 38012 40284
rect 38036 40282 38092 40284
rect 38116 40282 38172 40284
rect 38196 40282 38252 40284
rect 37956 40230 38002 40282
rect 38002 40230 38012 40282
rect 38036 40230 38066 40282
rect 38066 40230 38078 40282
rect 38078 40230 38092 40282
rect 38116 40230 38130 40282
rect 38130 40230 38142 40282
rect 38142 40230 38172 40282
rect 38196 40230 38206 40282
rect 38206 40230 38252 40282
rect 37956 40228 38012 40230
rect 38036 40228 38092 40230
rect 38116 40228 38172 40230
rect 38196 40228 38252 40230
rect 42956 53882 43012 53884
rect 43036 53882 43092 53884
rect 43116 53882 43172 53884
rect 43196 53882 43252 53884
rect 42956 53830 43002 53882
rect 43002 53830 43012 53882
rect 43036 53830 43066 53882
rect 43066 53830 43078 53882
rect 43078 53830 43092 53882
rect 43116 53830 43130 53882
rect 43130 53830 43142 53882
rect 43142 53830 43172 53882
rect 43196 53830 43206 53882
rect 43206 53830 43252 53882
rect 42956 53828 43012 53830
rect 43036 53828 43092 53830
rect 43116 53828 43172 53830
rect 43196 53828 43252 53830
rect 42956 52794 43012 52796
rect 43036 52794 43092 52796
rect 43116 52794 43172 52796
rect 43196 52794 43252 52796
rect 42956 52742 43002 52794
rect 43002 52742 43012 52794
rect 43036 52742 43066 52794
rect 43066 52742 43078 52794
rect 43078 52742 43092 52794
rect 43116 52742 43130 52794
rect 43130 52742 43142 52794
rect 43142 52742 43172 52794
rect 43196 52742 43206 52794
rect 43206 52742 43252 52794
rect 42956 52740 43012 52742
rect 43036 52740 43092 52742
rect 43116 52740 43172 52742
rect 43196 52740 43252 52742
rect 42956 51706 43012 51708
rect 43036 51706 43092 51708
rect 43116 51706 43172 51708
rect 43196 51706 43252 51708
rect 42956 51654 43002 51706
rect 43002 51654 43012 51706
rect 43036 51654 43066 51706
rect 43066 51654 43078 51706
rect 43078 51654 43092 51706
rect 43116 51654 43130 51706
rect 43130 51654 43142 51706
rect 43142 51654 43172 51706
rect 43196 51654 43206 51706
rect 43206 51654 43252 51706
rect 42956 51652 43012 51654
rect 43036 51652 43092 51654
rect 43116 51652 43172 51654
rect 43196 51652 43252 51654
rect 42956 50618 43012 50620
rect 43036 50618 43092 50620
rect 43116 50618 43172 50620
rect 43196 50618 43252 50620
rect 42956 50566 43002 50618
rect 43002 50566 43012 50618
rect 43036 50566 43066 50618
rect 43066 50566 43078 50618
rect 43078 50566 43092 50618
rect 43116 50566 43130 50618
rect 43130 50566 43142 50618
rect 43142 50566 43172 50618
rect 43196 50566 43206 50618
rect 43206 50566 43252 50618
rect 42956 50564 43012 50566
rect 43036 50564 43092 50566
rect 43116 50564 43172 50566
rect 43196 50564 43252 50566
rect 42956 49530 43012 49532
rect 43036 49530 43092 49532
rect 43116 49530 43172 49532
rect 43196 49530 43252 49532
rect 42956 49478 43002 49530
rect 43002 49478 43012 49530
rect 43036 49478 43066 49530
rect 43066 49478 43078 49530
rect 43078 49478 43092 49530
rect 43116 49478 43130 49530
rect 43130 49478 43142 49530
rect 43142 49478 43172 49530
rect 43196 49478 43206 49530
rect 43206 49478 43252 49530
rect 42956 49476 43012 49478
rect 43036 49476 43092 49478
rect 43116 49476 43172 49478
rect 43196 49476 43252 49478
rect 42956 48442 43012 48444
rect 43036 48442 43092 48444
rect 43116 48442 43172 48444
rect 43196 48442 43252 48444
rect 42956 48390 43002 48442
rect 43002 48390 43012 48442
rect 43036 48390 43066 48442
rect 43066 48390 43078 48442
rect 43078 48390 43092 48442
rect 43116 48390 43130 48442
rect 43130 48390 43142 48442
rect 43142 48390 43172 48442
rect 43196 48390 43206 48442
rect 43206 48390 43252 48442
rect 42956 48388 43012 48390
rect 43036 48388 43092 48390
rect 43116 48388 43172 48390
rect 43196 48388 43252 48390
rect 42956 47354 43012 47356
rect 43036 47354 43092 47356
rect 43116 47354 43172 47356
rect 43196 47354 43252 47356
rect 42956 47302 43002 47354
rect 43002 47302 43012 47354
rect 43036 47302 43066 47354
rect 43066 47302 43078 47354
rect 43078 47302 43092 47354
rect 43116 47302 43130 47354
rect 43130 47302 43142 47354
rect 43142 47302 43172 47354
rect 43196 47302 43206 47354
rect 43206 47302 43252 47354
rect 42956 47300 43012 47302
rect 43036 47300 43092 47302
rect 43116 47300 43172 47302
rect 43196 47300 43252 47302
rect 42956 46266 43012 46268
rect 43036 46266 43092 46268
rect 43116 46266 43172 46268
rect 43196 46266 43252 46268
rect 42956 46214 43002 46266
rect 43002 46214 43012 46266
rect 43036 46214 43066 46266
rect 43066 46214 43078 46266
rect 43078 46214 43092 46266
rect 43116 46214 43130 46266
rect 43130 46214 43142 46266
rect 43142 46214 43172 46266
rect 43196 46214 43206 46266
rect 43206 46214 43252 46266
rect 42956 46212 43012 46214
rect 43036 46212 43092 46214
rect 43116 46212 43172 46214
rect 43196 46212 43252 46214
rect 42956 45178 43012 45180
rect 43036 45178 43092 45180
rect 43116 45178 43172 45180
rect 43196 45178 43252 45180
rect 42956 45126 43002 45178
rect 43002 45126 43012 45178
rect 43036 45126 43066 45178
rect 43066 45126 43078 45178
rect 43078 45126 43092 45178
rect 43116 45126 43130 45178
rect 43130 45126 43142 45178
rect 43142 45126 43172 45178
rect 43196 45126 43206 45178
rect 43206 45126 43252 45178
rect 42956 45124 43012 45126
rect 43036 45124 43092 45126
rect 43116 45124 43172 45126
rect 43196 45124 43252 45126
rect 42956 44090 43012 44092
rect 43036 44090 43092 44092
rect 43116 44090 43172 44092
rect 43196 44090 43252 44092
rect 42956 44038 43002 44090
rect 43002 44038 43012 44090
rect 43036 44038 43066 44090
rect 43066 44038 43078 44090
rect 43078 44038 43092 44090
rect 43116 44038 43130 44090
rect 43130 44038 43142 44090
rect 43142 44038 43172 44090
rect 43196 44038 43206 44090
rect 43206 44038 43252 44090
rect 42956 44036 43012 44038
rect 43036 44036 43092 44038
rect 43116 44036 43172 44038
rect 43196 44036 43252 44038
rect 42956 43002 43012 43004
rect 43036 43002 43092 43004
rect 43116 43002 43172 43004
rect 43196 43002 43252 43004
rect 42956 42950 43002 43002
rect 43002 42950 43012 43002
rect 43036 42950 43066 43002
rect 43066 42950 43078 43002
rect 43078 42950 43092 43002
rect 43116 42950 43130 43002
rect 43130 42950 43142 43002
rect 43142 42950 43172 43002
rect 43196 42950 43206 43002
rect 43206 42950 43252 43002
rect 42956 42948 43012 42950
rect 43036 42948 43092 42950
rect 43116 42948 43172 42950
rect 43196 42948 43252 42950
rect 40222 42744 40278 42800
rect 38934 42608 38990 42664
rect 42956 41914 43012 41916
rect 43036 41914 43092 41916
rect 43116 41914 43172 41916
rect 43196 41914 43252 41916
rect 42956 41862 43002 41914
rect 43002 41862 43012 41914
rect 43036 41862 43066 41914
rect 43066 41862 43078 41914
rect 43078 41862 43092 41914
rect 43116 41862 43130 41914
rect 43130 41862 43142 41914
rect 43142 41862 43172 41914
rect 43196 41862 43206 41914
rect 43206 41862 43252 41914
rect 42956 41860 43012 41862
rect 43036 41860 43092 41862
rect 43116 41860 43172 41862
rect 43196 41860 43252 41862
rect 42956 40826 43012 40828
rect 43036 40826 43092 40828
rect 43116 40826 43172 40828
rect 43196 40826 43252 40828
rect 42956 40774 43002 40826
rect 43002 40774 43012 40826
rect 43036 40774 43066 40826
rect 43066 40774 43078 40826
rect 43078 40774 43092 40826
rect 43116 40774 43130 40826
rect 43130 40774 43142 40826
rect 43142 40774 43172 40826
rect 43196 40774 43206 40826
rect 43206 40774 43252 40826
rect 42956 40772 43012 40774
rect 43036 40772 43092 40774
rect 43116 40772 43172 40774
rect 43196 40772 43252 40774
rect 47956 54426 48012 54428
rect 48036 54426 48092 54428
rect 48116 54426 48172 54428
rect 48196 54426 48252 54428
rect 47956 54374 48002 54426
rect 48002 54374 48012 54426
rect 48036 54374 48066 54426
rect 48066 54374 48078 54426
rect 48078 54374 48092 54426
rect 48116 54374 48130 54426
rect 48130 54374 48142 54426
rect 48142 54374 48172 54426
rect 48196 54374 48206 54426
rect 48206 54374 48252 54426
rect 47956 54372 48012 54374
rect 48036 54372 48092 54374
rect 48116 54372 48172 54374
rect 48196 54372 48252 54374
rect 49054 54576 49110 54632
rect 47956 53338 48012 53340
rect 48036 53338 48092 53340
rect 48116 53338 48172 53340
rect 48196 53338 48252 53340
rect 47956 53286 48002 53338
rect 48002 53286 48012 53338
rect 48036 53286 48066 53338
rect 48066 53286 48078 53338
rect 48078 53286 48092 53338
rect 48116 53286 48130 53338
rect 48130 53286 48142 53338
rect 48142 53286 48172 53338
rect 48196 53286 48206 53338
rect 48206 53286 48252 53338
rect 47956 53284 48012 53286
rect 48036 53284 48092 53286
rect 48116 53284 48172 53286
rect 48196 53284 48252 53286
rect 47956 52250 48012 52252
rect 48036 52250 48092 52252
rect 48116 52250 48172 52252
rect 48196 52250 48252 52252
rect 47956 52198 48002 52250
rect 48002 52198 48012 52250
rect 48036 52198 48066 52250
rect 48066 52198 48078 52250
rect 48078 52198 48092 52250
rect 48116 52198 48130 52250
rect 48130 52198 48142 52250
rect 48142 52198 48172 52250
rect 48196 52198 48206 52250
rect 48206 52198 48252 52250
rect 47956 52196 48012 52198
rect 48036 52196 48092 52198
rect 48116 52196 48172 52198
rect 48196 52196 48252 52198
rect 47956 51162 48012 51164
rect 48036 51162 48092 51164
rect 48116 51162 48172 51164
rect 48196 51162 48252 51164
rect 47956 51110 48002 51162
rect 48002 51110 48012 51162
rect 48036 51110 48066 51162
rect 48066 51110 48078 51162
rect 48078 51110 48092 51162
rect 48116 51110 48130 51162
rect 48130 51110 48142 51162
rect 48142 51110 48172 51162
rect 48196 51110 48206 51162
rect 48206 51110 48252 51162
rect 47956 51108 48012 51110
rect 48036 51108 48092 51110
rect 48116 51108 48172 51110
rect 48196 51108 48252 51110
rect 47956 50074 48012 50076
rect 48036 50074 48092 50076
rect 48116 50074 48172 50076
rect 48196 50074 48252 50076
rect 47956 50022 48002 50074
rect 48002 50022 48012 50074
rect 48036 50022 48066 50074
rect 48066 50022 48078 50074
rect 48078 50022 48092 50074
rect 48116 50022 48130 50074
rect 48130 50022 48142 50074
rect 48142 50022 48172 50074
rect 48196 50022 48206 50074
rect 48206 50022 48252 50074
rect 47956 50020 48012 50022
rect 48036 50020 48092 50022
rect 48116 50020 48172 50022
rect 48196 50020 48252 50022
rect 47956 48986 48012 48988
rect 48036 48986 48092 48988
rect 48116 48986 48172 48988
rect 48196 48986 48252 48988
rect 47956 48934 48002 48986
rect 48002 48934 48012 48986
rect 48036 48934 48066 48986
rect 48066 48934 48078 48986
rect 48078 48934 48092 48986
rect 48116 48934 48130 48986
rect 48130 48934 48142 48986
rect 48142 48934 48172 48986
rect 48196 48934 48206 48986
rect 48206 48934 48252 48986
rect 47956 48932 48012 48934
rect 48036 48932 48092 48934
rect 48116 48932 48172 48934
rect 48196 48932 48252 48934
rect 47956 47898 48012 47900
rect 48036 47898 48092 47900
rect 48116 47898 48172 47900
rect 48196 47898 48252 47900
rect 47956 47846 48002 47898
rect 48002 47846 48012 47898
rect 48036 47846 48066 47898
rect 48066 47846 48078 47898
rect 48078 47846 48092 47898
rect 48116 47846 48130 47898
rect 48130 47846 48142 47898
rect 48142 47846 48172 47898
rect 48196 47846 48206 47898
rect 48206 47846 48252 47898
rect 47956 47844 48012 47846
rect 48036 47844 48092 47846
rect 48116 47844 48172 47846
rect 48196 47844 48252 47846
rect 47956 46810 48012 46812
rect 48036 46810 48092 46812
rect 48116 46810 48172 46812
rect 48196 46810 48252 46812
rect 47956 46758 48002 46810
rect 48002 46758 48012 46810
rect 48036 46758 48066 46810
rect 48066 46758 48078 46810
rect 48078 46758 48092 46810
rect 48116 46758 48130 46810
rect 48130 46758 48142 46810
rect 48142 46758 48172 46810
rect 48196 46758 48206 46810
rect 48206 46758 48252 46810
rect 47956 46756 48012 46758
rect 48036 46756 48092 46758
rect 48116 46756 48172 46758
rect 48196 46756 48252 46758
rect 42956 39738 43012 39740
rect 43036 39738 43092 39740
rect 43116 39738 43172 39740
rect 43196 39738 43252 39740
rect 42956 39686 43002 39738
rect 43002 39686 43012 39738
rect 43036 39686 43066 39738
rect 43066 39686 43078 39738
rect 43078 39686 43092 39738
rect 43116 39686 43130 39738
rect 43130 39686 43142 39738
rect 43142 39686 43172 39738
rect 43196 39686 43206 39738
rect 43206 39686 43252 39738
rect 42956 39684 43012 39686
rect 43036 39684 43092 39686
rect 43116 39684 43172 39686
rect 43196 39684 43252 39686
rect 37956 39194 38012 39196
rect 38036 39194 38092 39196
rect 38116 39194 38172 39196
rect 38196 39194 38252 39196
rect 37956 39142 38002 39194
rect 38002 39142 38012 39194
rect 38036 39142 38066 39194
rect 38066 39142 38078 39194
rect 38078 39142 38092 39194
rect 38116 39142 38130 39194
rect 38130 39142 38142 39194
rect 38142 39142 38172 39194
rect 38196 39142 38206 39194
rect 38206 39142 38252 39194
rect 37956 39140 38012 39142
rect 38036 39140 38092 39142
rect 38116 39140 38172 39142
rect 38196 39140 38252 39142
rect 42956 38650 43012 38652
rect 43036 38650 43092 38652
rect 43116 38650 43172 38652
rect 43196 38650 43252 38652
rect 42956 38598 43002 38650
rect 43002 38598 43012 38650
rect 43036 38598 43066 38650
rect 43066 38598 43078 38650
rect 43078 38598 43092 38650
rect 43116 38598 43130 38650
rect 43130 38598 43142 38650
rect 43142 38598 43172 38650
rect 43196 38598 43206 38650
rect 43206 38598 43252 38650
rect 42956 38596 43012 38598
rect 43036 38596 43092 38598
rect 43116 38596 43172 38598
rect 43196 38596 43252 38598
rect 37956 38106 38012 38108
rect 38036 38106 38092 38108
rect 38116 38106 38172 38108
rect 38196 38106 38252 38108
rect 37956 38054 38002 38106
rect 38002 38054 38012 38106
rect 38036 38054 38066 38106
rect 38066 38054 38078 38106
rect 38078 38054 38092 38106
rect 38116 38054 38130 38106
rect 38130 38054 38142 38106
rect 38142 38054 38172 38106
rect 38196 38054 38206 38106
rect 38206 38054 38252 38106
rect 37956 38052 38012 38054
rect 38036 38052 38092 38054
rect 38116 38052 38172 38054
rect 38196 38052 38252 38054
rect 42956 37562 43012 37564
rect 43036 37562 43092 37564
rect 43116 37562 43172 37564
rect 43196 37562 43252 37564
rect 42956 37510 43002 37562
rect 43002 37510 43012 37562
rect 43036 37510 43066 37562
rect 43066 37510 43078 37562
rect 43078 37510 43092 37562
rect 43116 37510 43130 37562
rect 43130 37510 43142 37562
rect 43142 37510 43172 37562
rect 43196 37510 43206 37562
rect 43206 37510 43252 37562
rect 42956 37508 43012 37510
rect 43036 37508 43092 37510
rect 43116 37508 43172 37510
rect 43196 37508 43252 37510
rect 37956 37018 38012 37020
rect 38036 37018 38092 37020
rect 38116 37018 38172 37020
rect 38196 37018 38252 37020
rect 37956 36966 38002 37018
rect 38002 36966 38012 37018
rect 38036 36966 38066 37018
rect 38066 36966 38078 37018
rect 38078 36966 38092 37018
rect 38116 36966 38130 37018
rect 38130 36966 38142 37018
rect 38142 36966 38172 37018
rect 38196 36966 38206 37018
rect 38206 36966 38252 37018
rect 37956 36964 38012 36966
rect 38036 36964 38092 36966
rect 38116 36964 38172 36966
rect 38196 36964 38252 36966
rect 42956 36474 43012 36476
rect 43036 36474 43092 36476
rect 43116 36474 43172 36476
rect 43196 36474 43252 36476
rect 42956 36422 43002 36474
rect 43002 36422 43012 36474
rect 43036 36422 43066 36474
rect 43066 36422 43078 36474
rect 43078 36422 43092 36474
rect 43116 36422 43130 36474
rect 43130 36422 43142 36474
rect 43142 36422 43172 36474
rect 43196 36422 43206 36474
rect 43206 36422 43252 36474
rect 42956 36420 43012 36422
rect 43036 36420 43092 36422
rect 43116 36420 43172 36422
rect 43196 36420 43252 36422
rect 37956 35930 38012 35932
rect 38036 35930 38092 35932
rect 38116 35930 38172 35932
rect 38196 35930 38252 35932
rect 37956 35878 38002 35930
rect 38002 35878 38012 35930
rect 38036 35878 38066 35930
rect 38066 35878 38078 35930
rect 38078 35878 38092 35930
rect 38116 35878 38130 35930
rect 38130 35878 38142 35930
rect 38142 35878 38172 35930
rect 38196 35878 38206 35930
rect 38206 35878 38252 35930
rect 37956 35876 38012 35878
rect 38036 35876 38092 35878
rect 38116 35876 38172 35878
rect 38196 35876 38252 35878
rect 42956 35386 43012 35388
rect 43036 35386 43092 35388
rect 43116 35386 43172 35388
rect 43196 35386 43252 35388
rect 42956 35334 43002 35386
rect 43002 35334 43012 35386
rect 43036 35334 43066 35386
rect 43066 35334 43078 35386
rect 43078 35334 43092 35386
rect 43116 35334 43130 35386
rect 43130 35334 43142 35386
rect 43142 35334 43172 35386
rect 43196 35334 43206 35386
rect 43206 35334 43252 35386
rect 42956 35332 43012 35334
rect 43036 35332 43092 35334
rect 43116 35332 43172 35334
rect 43196 35332 43252 35334
rect 37956 34842 38012 34844
rect 38036 34842 38092 34844
rect 38116 34842 38172 34844
rect 38196 34842 38252 34844
rect 37956 34790 38002 34842
rect 38002 34790 38012 34842
rect 38036 34790 38066 34842
rect 38066 34790 38078 34842
rect 38078 34790 38092 34842
rect 38116 34790 38130 34842
rect 38130 34790 38142 34842
rect 38142 34790 38172 34842
rect 38196 34790 38206 34842
rect 38206 34790 38252 34842
rect 37956 34788 38012 34790
rect 38036 34788 38092 34790
rect 38116 34788 38172 34790
rect 38196 34788 38252 34790
rect 42956 34298 43012 34300
rect 43036 34298 43092 34300
rect 43116 34298 43172 34300
rect 43196 34298 43252 34300
rect 42956 34246 43002 34298
rect 43002 34246 43012 34298
rect 43036 34246 43066 34298
rect 43066 34246 43078 34298
rect 43078 34246 43092 34298
rect 43116 34246 43130 34298
rect 43130 34246 43142 34298
rect 43142 34246 43172 34298
rect 43196 34246 43206 34298
rect 43206 34246 43252 34298
rect 42956 34244 43012 34246
rect 43036 34244 43092 34246
rect 43116 34244 43172 34246
rect 43196 34244 43252 34246
rect 37956 33754 38012 33756
rect 38036 33754 38092 33756
rect 38116 33754 38172 33756
rect 38196 33754 38252 33756
rect 37956 33702 38002 33754
rect 38002 33702 38012 33754
rect 38036 33702 38066 33754
rect 38066 33702 38078 33754
rect 38078 33702 38092 33754
rect 38116 33702 38130 33754
rect 38130 33702 38142 33754
rect 38142 33702 38172 33754
rect 38196 33702 38206 33754
rect 38206 33702 38252 33754
rect 37956 33700 38012 33702
rect 38036 33700 38092 33702
rect 38116 33700 38172 33702
rect 38196 33700 38252 33702
rect 42956 33210 43012 33212
rect 43036 33210 43092 33212
rect 43116 33210 43172 33212
rect 43196 33210 43252 33212
rect 42956 33158 43002 33210
rect 43002 33158 43012 33210
rect 43036 33158 43066 33210
rect 43066 33158 43078 33210
rect 43078 33158 43092 33210
rect 43116 33158 43130 33210
rect 43130 33158 43142 33210
rect 43142 33158 43172 33210
rect 43196 33158 43206 33210
rect 43206 33158 43252 33210
rect 42956 33156 43012 33158
rect 43036 33156 43092 33158
rect 43116 33156 43172 33158
rect 43196 33156 43252 33158
rect 37956 32666 38012 32668
rect 38036 32666 38092 32668
rect 38116 32666 38172 32668
rect 38196 32666 38252 32668
rect 37956 32614 38002 32666
rect 38002 32614 38012 32666
rect 38036 32614 38066 32666
rect 38066 32614 38078 32666
rect 38078 32614 38092 32666
rect 38116 32614 38130 32666
rect 38130 32614 38142 32666
rect 38142 32614 38172 32666
rect 38196 32614 38206 32666
rect 38206 32614 38252 32666
rect 37956 32612 38012 32614
rect 38036 32612 38092 32614
rect 38116 32612 38172 32614
rect 38196 32612 38252 32614
rect 42956 32122 43012 32124
rect 43036 32122 43092 32124
rect 43116 32122 43172 32124
rect 43196 32122 43252 32124
rect 42956 32070 43002 32122
rect 43002 32070 43012 32122
rect 43036 32070 43066 32122
rect 43066 32070 43078 32122
rect 43078 32070 43092 32122
rect 43116 32070 43130 32122
rect 43130 32070 43142 32122
rect 43142 32070 43172 32122
rect 43196 32070 43206 32122
rect 43206 32070 43252 32122
rect 42956 32068 43012 32070
rect 43036 32068 43092 32070
rect 43116 32068 43172 32070
rect 43196 32068 43252 32070
rect 37956 31578 38012 31580
rect 38036 31578 38092 31580
rect 38116 31578 38172 31580
rect 38196 31578 38252 31580
rect 37956 31526 38002 31578
rect 38002 31526 38012 31578
rect 38036 31526 38066 31578
rect 38066 31526 38078 31578
rect 38078 31526 38092 31578
rect 38116 31526 38130 31578
rect 38130 31526 38142 31578
rect 38142 31526 38172 31578
rect 38196 31526 38206 31578
rect 38206 31526 38252 31578
rect 37956 31524 38012 31526
rect 38036 31524 38092 31526
rect 38116 31524 38172 31526
rect 38196 31524 38252 31526
rect 42956 31034 43012 31036
rect 43036 31034 43092 31036
rect 43116 31034 43172 31036
rect 43196 31034 43252 31036
rect 42956 30982 43002 31034
rect 43002 30982 43012 31034
rect 43036 30982 43066 31034
rect 43066 30982 43078 31034
rect 43078 30982 43092 31034
rect 43116 30982 43130 31034
rect 43130 30982 43142 31034
rect 43142 30982 43172 31034
rect 43196 30982 43206 31034
rect 43206 30982 43252 31034
rect 42956 30980 43012 30982
rect 43036 30980 43092 30982
rect 43116 30980 43172 30982
rect 43196 30980 43252 30982
rect 37956 30490 38012 30492
rect 38036 30490 38092 30492
rect 38116 30490 38172 30492
rect 38196 30490 38252 30492
rect 37956 30438 38002 30490
rect 38002 30438 38012 30490
rect 38036 30438 38066 30490
rect 38066 30438 38078 30490
rect 38078 30438 38092 30490
rect 38116 30438 38130 30490
rect 38130 30438 38142 30490
rect 38142 30438 38172 30490
rect 38196 30438 38206 30490
rect 38206 30438 38252 30490
rect 37956 30436 38012 30438
rect 38036 30436 38092 30438
rect 38116 30436 38172 30438
rect 38196 30436 38252 30438
rect 42956 29946 43012 29948
rect 43036 29946 43092 29948
rect 43116 29946 43172 29948
rect 43196 29946 43252 29948
rect 42956 29894 43002 29946
rect 43002 29894 43012 29946
rect 43036 29894 43066 29946
rect 43066 29894 43078 29946
rect 43078 29894 43092 29946
rect 43116 29894 43130 29946
rect 43130 29894 43142 29946
rect 43142 29894 43172 29946
rect 43196 29894 43206 29946
rect 43206 29894 43252 29946
rect 42956 29892 43012 29894
rect 43036 29892 43092 29894
rect 43116 29892 43172 29894
rect 43196 29892 43252 29894
rect 37956 29402 38012 29404
rect 38036 29402 38092 29404
rect 38116 29402 38172 29404
rect 38196 29402 38252 29404
rect 37956 29350 38002 29402
rect 38002 29350 38012 29402
rect 38036 29350 38066 29402
rect 38066 29350 38078 29402
rect 38078 29350 38092 29402
rect 38116 29350 38130 29402
rect 38130 29350 38142 29402
rect 38142 29350 38172 29402
rect 38196 29350 38206 29402
rect 38206 29350 38252 29402
rect 37956 29348 38012 29350
rect 38036 29348 38092 29350
rect 38116 29348 38172 29350
rect 38196 29348 38252 29350
rect 42956 28858 43012 28860
rect 43036 28858 43092 28860
rect 43116 28858 43172 28860
rect 43196 28858 43252 28860
rect 42956 28806 43002 28858
rect 43002 28806 43012 28858
rect 43036 28806 43066 28858
rect 43066 28806 43078 28858
rect 43078 28806 43092 28858
rect 43116 28806 43130 28858
rect 43130 28806 43142 28858
rect 43142 28806 43172 28858
rect 43196 28806 43206 28858
rect 43206 28806 43252 28858
rect 42956 28804 43012 28806
rect 43036 28804 43092 28806
rect 43116 28804 43172 28806
rect 43196 28804 43252 28806
rect 37956 28314 38012 28316
rect 38036 28314 38092 28316
rect 38116 28314 38172 28316
rect 38196 28314 38252 28316
rect 37956 28262 38002 28314
rect 38002 28262 38012 28314
rect 38036 28262 38066 28314
rect 38066 28262 38078 28314
rect 38078 28262 38092 28314
rect 38116 28262 38130 28314
rect 38130 28262 38142 28314
rect 38142 28262 38172 28314
rect 38196 28262 38206 28314
rect 38206 28262 38252 28314
rect 37956 28260 38012 28262
rect 38036 28260 38092 28262
rect 38116 28260 38172 28262
rect 38196 28260 38252 28262
rect 42956 27770 43012 27772
rect 43036 27770 43092 27772
rect 43116 27770 43172 27772
rect 43196 27770 43252 27772
rect 42956 27718 43002 27770
rect 43002 27718 43012 27770
rect 43036 27718 43066 27770
rect 43066 27718 43078 27770
rect 43078 27718 43092 27770
rect 43116 27718 43130 27770
rect 43130 27718 43142 27770
rect 43142 27718 43172 27770
rect 43196 27718 43206 27770
rect 43206 27718 43252 27770
rect 42956 27716 43012 27718
rect 43036 27716 43092 27718
rect 43116 27716 43172 27718
rect 43196 27716 43252 27718
rect 37956 27226 38012 27228
rect 38036 27226 38092 27228
rect 38116 27226 38172 27228
rect 38196 27226 38252 27228
rect 37956 27174 38002 27226
rect 38002 27174 38012 27226
rect 38036 27174 38066 27226
rect 38066 27174 38078 27226
rect 38078 27174 38092 27226
rect 38116 27174 38130 27226
rect 38130 27174 38142 27226
rect 38142 27174 38172 27226
rect 38196 27174 38206 27226
rect 38206 27174 38252 27226
rect 37956 27172 38012 27174
rect 38036 27172 38092 27174
rect 38116 27172 38172 27174
rect 38196 27172 38252 27174
rect 42956 26682 43012 26684
rect 43036 26682 43092 26684
rect 43116 26682 43172 26684
rect 43196 26682 43252 26684
rect 42956 26630 43002 26682
rect 43002 26630 43012 26682
rect 43036 26630 43066 26682
rect 43066 26630 43078 26682
rect 43078 26630 43092 26682
rect 43116 26630 43130 26682
rect 43130 26630 43142 26682
rect 43142 26630 43172 26682
rect 43196 26630 43206 26682
rect 43206 26630 43252 26682
rect 42956 26628 43012 26630
rect 43036 26628 43092 26630
rect 43116 26628 43172 26630
rect 43196 26628 43252 26630
rect 37956 26138 38012 26140
rect 38036 26138 38092 26140
rect 38116 26138 38172 26140
rect 38196 26138 38252 26140
rect 37956 26086 38002 26138
rect 38002 26086 38012 26138
rect 38036 26086 38066 26138
rect 38066 26086 38078 26138
rect 38078 26086 38092 26138
rect 38116 26086 38130 26138
rect 38130 26086 38142 26138
rect 38142 26086 38172 26138
rect 38196 26086 38206 26138
rect 38206 26086 38252 26138
rect 37956 26084 38012 26086
rect 38036 26084 38092 26086
rect 38116 26084 38172 26086
rect 38196 26084 38252 26086
rect 42956 25594 43012 25596
rect 43036 25594 43092 25596
rect 43116 25594 43172 25596
rect 43196 25594 43252 25596
rect 42956 25542 43002 25594
rect 43002 25542 43012 25594
rect 43036 25542 43066 25594
rect 43066 25542 43078 25594
rect 43078 25542 43092 25594
rect 43116 25542 43130 25594
rect 43130 25542 43142 25594
rect 43142 25542 43172 25594
rect 43196 25542 43206 25594
rect 43206 25542 43252 25594
rect 42956 25540 43012 25542
rect 43036 25540 43092 25542
rect 43116 25540 43172 25542
rect 43196 25540 43252 25542
rect 37956 25050 38012 25052
rect 38036 25050 38092 25052
rect 38116 25050 38172 25052
rect 38196 25050 38252 25052
rect 37956 24998 38002 25050
rect 38002 24998 38012 25050
rect 38036 24998 38066 25050
rect 38066 24998 38078 25050
rect 38078 24998 38092 25050
rect 38116 24998 38130 25050
rect 38130 24998 38142 25050
rect 38142 24998 38172 25050
rect 38196 24998 38206 25050
rect 38206 24998 38252 25050
rect 37956 24996 38012 24998
rect 38036 24996 38092 24998
rect 38116 24996 38172 24998
rect 38196 24996 38252 24998
rect 47956 45722 48012 45724
rect 48036 45722 48092 45724
rect 48116 45722 48172 45724
rect 48196 45722 48252 45724
rect 47956 45670 48002 45722
rect 48002 45670 48012 45722
rect 48036 45670 48066 45722
rect 48066 45670 48078 45722
rect 48078 45670 48092 45722
rect 48116 45670 48130 45722
rect 48130 45670 48142 45722
rect 48142 45670 48172 45722
rect 48196 45670 48206 45722
rect 48206 45670 48252 45722
rect 47956 45668 48012 45670
rect 48036 45668 48092 45670
rect 48116 45668 48172 45670
rect 48196 45668 48252 45670
rect 47956 44634 48012 44636
rect 48036 44634 48092 44636
rect 48116 44634 48172 44636
rect 48196 44634 48252 44636
rect 47956 44582 48002 44634
rect 48002 44582 48012 44634
rect 48036 44582 48066 44634
rect 48066 44582 48078 44634
rect 48078 44582 48092 44634
rect 48116 44582 48130 44634
rect 48130 44582 48142 44634
rect 48142 44582 48172 44634
rect 48196 44582 48206 44634
rect 48206 44582 48252 44634
rect 47956 44580 48012 44582
rect 48036 44580 48092 44582
rect 48116 44580 48172 44582
rect 48196 44580 48252 44582
rect 47956 43546 48012 43548
rect 48036 43546 48092 43548
rect 48116 43546 48172 43548
rect 48196 43546 48252 43548
rect 47956 43494 48002 43546
rect 48002 43494 48012 43546
rect 48036 43494 48066 43546
rect 48066 43494 48078 43546
rect 48078 43494 48092 43546
rect 48116 43494 48130 43546
rect 48130 43494 48142 43546
rect 48142 43494 48172 43546
rect 48196 43494 48206 43546
rect 48206 43494 48252 43546
rect 47956 43492 48012 43494
rect 48036 43492 48092 43494
rect 48116 43492 48172 43494
rect 48196 43492 48252 43494
rect 47956 42458 48012 42460
rect 48036 42458 48092 42460
rect 48116 42458 48172 42460
rect 48196 42458 48252 42460
rect 47956 42406 48002 42458
rect 48002 42406 48012 42458
rect 48036 42406 48066 42458
rect 48066 42406 48078 42458
rect 48078 42406 48092 42458
rect 48116 42406 48130 42458
rect 48130 42406 48142 42458
rect 48142 42406 48172 42458
rect 48196 42406 48206 42458
rect 48206 42406 48252 42458
rect 47956 42404 48012 42406
rect 48036 42404 48092 42406
rect 48116 42404 48172 42406
rect 48196 42404 48252 42406
rect 47956 41370 48012 41372
rect 48036 41370 48092 41372
rect 48116 41370 48172 41372
rect 48196 41370 48252 41372
rect 47956 41318 48002 41370
rect 48002 41318 48012 41370
rect 48036 41318 48066 41370
rect 48066 41318 48078 41370
rect 48078 41318 48092 41370
rect 48116 41318 48130 41370
rect 48130 41318 48142 41370
rect 48142 41318 48172 41370
rect 48196 41318 48206 41370
rect 48206 41318 48252 41370
rect 47956 41316 48012 41318
rect 48036 41316 48092 41318
rect 48116 41316 48172 41318
rect 48196 41316 48252 41318
rect 47956 40282 48012 40284
rect 48036 40282 48092 40284
rect 48116 40282 48172 40284
rect 48196 40282 48252 40284
rect 47956 40230 48002 40282
rect 48002 40230 48012 40282
rect 48036 40230 48066 40282
rect 48066 40230 48078 40282
rect 48078 40230 48092 40282
rect 48116 40230 48130 40282
rect 48130 40230 48142 40282
rect 48142 40230 48172 40282
rect 48196 40230 48206 40282
rect 48206 40230 48252 40282
rect 47956 40228 48012 40230
rect 48036 40228 48092 40230
rect 48116 40228 48172 40230
rect 48196 40228 48252 40230
rect 47956 39194 48012 39196
rect 48036 39194 48092 39196
rect 48116 39194 48172 39196
rect 48196 39194 48252 39196
rect 47956 39142 48002 39194
rect 48002 39142 48012 39194
rect 48036 39142 48066 39194
rect 48066 39142 48078 39194
rect 48078 39142 48092 39194
rect 48116 39142 48130 39194
rect 48130 39142 48142 39194
rect 48142 39142 48172 39194
rect 48196 39142 48206 39194
rect 48206 39142 48252 39194
rect 47956 39140 48012 39142
rect 48036 39140 48092 39142
rect 48116 39140 48172 39142
rect 48196 39140 48252 39142
rect 49054 52436 49056 52456
rect 49056 52436 49108 52456
rect 49108 52436 49110 52456
rect 49054 52400 49110 52436
rect 49054 50260 49056 50280
rect 49056 50260 49108 50280
rect 49108 50260 49110 50280
rect 49054 50224 49110 50260
rect 48962 48068 49018 48104
rect 48962 48048 48964 48068
rect 48964 48048 49016 48068
rect 49016 48048 49018 48068
rect 49146 45908 49148 45928
rect 49148 45908 49200 45928
rect 49200 45908 49202 45928
rect 49146 45872 49202 45908
rect 47956 38106 48012 38108
rect 48036 38106 48092 38108
rect 48116 38106 48172 38108
rect 48196 38106 48252 38108
rect 47956 38054 48002 38106
rect 48002 38054 48012 38106
rect 48036 38054 48066 38106
rect 48066 38054 48078 38106
rect 48078 38054 48092 38106
rect 48116 38054 48130 38106
rect 48130 38054 48142 38106
rect 48142 38054 48172 38106
rect 48196 38054 48206 38106
rect 48206 38054 48252 38106
rect 47956 38052 48012 38054
rect 48036 38052 48092 38054
rect 48116 38052 48172 38054
rect 48196 38052 48252 38054
rect 47956 37018 48012 37020
rect 48036 37018 48092 37020
rect 48116 37018 48172 37020
rect 48196 37018 48252 37020
rect 47956 36966 48002 37018
rect 48002 36966 48012 37018
rect 48036 36966 48066 37018
rect 48066 36966 48078 37018
rect 48078 36966 48092 37018
rect 48116 36966 48130 37018
rect 48130 36966 48142 37018
rect 48142 36966 48172 37018
rect 48196 36966 48206 37018
rect 48206 36966 48252 37018
rect 47956 36964 48012 36966
rect 48036 36964 48092 36966
rect 48116 36964 48172 36966
rect 48196 36964 48252 36966
rect 47956 35930 48012 35932
rect 48036 35930 48092 35932
rect 48116 35930 48172 35932
rect 48196 35930 48252 35932
rect 47956 35878 48002 35930
rect 48002 35878 48012 35930
rect 48036 35878 48066 35930
rect 48066 35878 48078 35930
rect 48078 35878 48092 35930
rect 48116 35878 48130 35930
rect 48130 35878 48142 35930
rect 48142 35878 48172 35930
rect 48196 35878 48206 35930
rect 48206 35878 48252 35930
rect 47956 35876 48012 35878
rect 48036 35876 48092 35878
rect 48116 35876 48172 35878
rect 48196 35876 48252 35878
rect 47956 34842 48012 34844
rect 48036 34842 48092 34844
rect 48116 34842 48172 34844
rect 48196 34842 48252 34844
rect 47956 34790 48002 34842
rect 48002 34790 48012 34842
rect 48036 34790 48066 34842
rect 48066 34790 48078 34842
rect 48078 34790 48092 34842
rect 48116 34790 48130 34842
rect 48130 34790 48142 34842
rect 48142 34790 48172 34842
rect 48196 34790 48206 34842
rect 48206 34790 48252 34842
rect 47956 34788 48012 34790
rect 48036 34788 48092 34790
rect 48116 34788 48172 34790
rect 48196 34788 48252 34790
rect 47956 33754 48012 33756
rect 48036 33754 48092 33756
rect 48116 33754 48172 33756
rect 48196 33754 48252 33756
rect 47956 33702 48002 33754
rect 48002 33702 48012 33754
rect 48036 33702 48066 33754
rect 48066 33702 48078 33754
rect 48078 33702 48092 33754
rect 48116 33702 48130 33754
rect 48130 33702 48142 33754
rect 48142 33702 48172 33754
rect 48196 33702 48206 33754
rect 48206 33702 48252 33754
rect 47956 33700 48012 33702
rect 48036 33700 48092 33702
rect 48116 33700 48172 33702
rect 48196 33700 48252 33702
rect 47956 32666 48012 32668
rect 48036 32666 48092 32668
rect 48116 32666 48172 32668
rect 48196 32666 48252 32668
rect 47956 32614 48002 32666
rect 48002 32614 48012 32666
rect 48036 32614 48066 32666
rect 48066 32614 48078 32666
rect 48078 32614 48092 32666
rect 48116 32614 48130 32666
rect 48130 32614 48142 32666
rect 48142 32614 48172 32666
rect 48196 32614 48206 32666
rect 48206 32614 48252 32666
rect 47956 32612 48012 32614
rect 48036 32612 48092 32614
rect 48116 32612 48172 32614
rect 48196 32612 48252 32614
rect 47956 31578 48012 31580
rect 48036 31578 48092 31580
rect 48116 31578 48172 31580
rect 48196 31578 48252 31580
rect 47956 31526 48002 31578
rect 48002 31526 48012 31578
rect 48036 31526 48066 31578
rect 48066 31526 48078 31578
rect 48078 31526 48092 31578
rect 48116 31526 48130 31578
rect 48130 31526 48142 31578
rect 48142 31526 48172 31578
rect 48196 31526 48206 31578
rect 48206 31526 48252 31578
rect 47956 31524 48012 31526
rect 48036 31524 48092 31526
rect 48116 31524 48172 31526
rect 48196 31524 48252 31526
rect 47956 30490 48012 30492
rect 48036 30490 48092 30492
rect 48116 30490 48172 30492
rect 48196 30490 48252 30492
rect 47956 30438 48002 30490
rect 48002 30438 48012 30490
rect 48036 30438 48066 30490
rect 48066 30438 48078 30490
rect 48078 30438 48092 30490
rect 48116 30438 48130 30490
rect 48130 30438 48142 30490
rect 48142 30438 48172 30490
rect 48196 30438 48206 30490
rect 48206 30438 48252 30490
rect 47956 30436 48012 30438
rect 48036 30436 48092 30438
rect 48116 30436 48172 30438
rect 48196 30436 48252 30438
rect 47956 29402 48012 29404
rect 48036 29402 48092 29404
rect 48116 29402 48172 29404
rect 48196 29402 48252 29404
rect 47956 29350 48002 29402
rect 48002 29350 48012 29402
rect 48036 29350 48066 29402
rect 48066 29350 48078 29402
rect 48078 29350 48092 29402
rect 48116 29350 48130 29402
rect 48130 29350 48142 29402
rect 48142 29350 48172 29402
rect 48196 29350 48206 29402
rect 48206 29350 48252 29402
rect 47956 29348 48012 29350
rect 48036 29348 48092 29350
rect 48116 29348 48172 29350
rect 48196 29348 48252 29350
rect 47956 28314 48012 28316
rect 48036 28314 48092 28316
rect 48116 28314 48172 28316
rect 48196 28314 48252 28316
rect 47956 28262 48002 28314
rect 48002 28262 48012 28314
rect 48036 28262 48066 28314
rect 48066 28262 48078 28314
rect 48078 28262 48092 28314
rect 48116 28262 48130 28314
rect 48130 28262 48142 28314
rect 48142 28262 48172 28314
rect 48196 28262 48206 28314
rect 48206 28262 48252 28314
rect 47956 28260 48012 28262
rect 48036 28260 48092 28262
rect 48116 28260 48172 28262
rect 48196 28260 48252 28262
rect 47956 27226 48012 27228
rect 48036 27226 48092 27228
rect 48116 27226 48172 27228
rect 48196 27226 48252 27228
rect 47956 27174 48002 27226
rect 48002 27174 48012 27226
rect 48036 27174 48066 27226
rect 48066 27174 48078 27226
rect 48078 27174 48092 27226
rect 48116 27174 48130 27226
rect 48130 27174 48142 27226
rect 48142 27174 48172 27226
rect 48196 27174 48206 27226
rect 48206 27174 48252 27226
rect 47956 27172 48012 27174
rect 48036 27172 48092 27174
rect 48116 27172 48172 27174
rect 48196 27172 48252 27174
rect 47956 26138 48012 26140
rect 48036 26138 48092 26140
rect 48116 26138 48172 26140
rect 48196 26138 48252 26140
rect 47956 26086 48002 26138
rect 48002 26086 48012 26138
rect 48036 26086 48066 26138
rect 48066 26086 48078 26138
rect 48078 26086 48092 26138
rect 48116 26086 48130 26138
rect 48130 26086 48142 26138
rect 48142 26086 48172 26138
rect 48196 26086 48206 26138
rect 48206 26086 48252 26138
rect 47956 26084 48012 26086
rect 48036 26084 48092 26086
rect 48116 26084 48172 26086
rect 48196 26084 48252 26086
rect 47956 25050 48012 25052
rect 48036 25050 48092 25052
rect 48116 25050 48172 25052
rect 48196 25050 48252 25052
rect 47956 24998 48002 25050
rect 48002 24998 48012 25050
rect 48036 24998 48066 25050
rect 48066 24998 48078 25050
rect 48078 24998 48092 25050
rect 48116 24998 48130 25050
rect 48130 24998 48142 25050
rect 48142 24998 48172 25050
rect 48196 24998 48206 25050
rect 48206 24998 48252 25050
rect 47956 24996 48012 24998
rect 48036 24996 48092 24998
rect 48116 24996 48172 24998
rect 48196 24996 48252 24998
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
<< metal3 >>
rect 0 54634 800 54664
rect 3417 54634 3483 54637
rect 0 54632 3483 54634
rect 0 54576 3422 54632
rect 3478 54576 3483 54632
rect 0 54574 3483 54576
rect 0 54544 800 54574
rect 3417 54571 3483 54574
rect 49049 54634 49115 54637
rect 50200 54634 51000 54664
rect 49049 54632 51000 54634
rect 49049 54576 49054 54632
rect 49110 54576 51000 54632
rect 49049 54574 51000 54576
rect 49049 54571 49115 54574
rect 50200 54544 51000 54574
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 27946 54432 28262 54433
rect 27946 54368 27952 54432
rect 28016 54368 28032 54432
rect 28096 54368 28112 54432
rect 28176 54368 28192 54432
rect 28256 54368 28262 54432
rect 27946 54367 28262 54368
rect 37946 54432 38262 54433
rect 37946 54368 37952 54432
rect 38016 54368 38032 54432
rect 38096 54368 38112 54432
rect 38176 54368 38192 54432
rect 38256 54368 38262 54432
rect 37946 54367 38262 54368
rect 47946 54432 48262 54433
rect 47946 54368 47952 54432
rect 48016 54368 48032 54432
rect 48096 54368 48112 54432
rect 48176 54368 48192 54432
rect 48256 54368 48262 54432
rect 47946 54367 48262 54368
rect 11094 54028 11100 54092
rect 11164 54090 11170 54092
rect 35065 54090 35131 54093
rect 11164 54088 35131 54090
rect 11164 54032 35070 54088
rect 35126 54032 35131 54088
rect 11164 54030 35131 54032
rect 11164 54028 11170 54030
rect 35065 54027 35131 54030
rect 2946 53888 3262 53889
rect 0 53818 800 53848
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 32946 53888 33262 53889
rect 32946 53824 32952 53888
rect 33016 53824 33032 53888
rect 33096 53824 33112 53888
rect 33176 53824 33192 53888
rect 33256 53824 33262 53888
rect 32946 53823 33262 53824
rect 42946 53888 43262 53889
rect 42946 53824 42952 53888
rect 43016 53824 43032 53888
rect 43096 53824 43112 53888
rect 43176 53824 43192 53888
rect 43256 53824 43262 53888
rect 42946 53823 43262 53824
rect 2773 53818 2839 53821
rect 0 53816 2839 53818
rect 0 53760 2778 53816
rect 2834 53760 2839 53816
rect 0 53758 2839 53760
rect 0 53728 800 53758
rect 2773 53755 2839 53758
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 27946 53344 28262 53345
rect 27946 53280 27952 53344
rect 28016 53280 28032 53344
rect 28096 53280 28112 53344
rect 28176 53280 28192 53344
rect 28256 53280 28262 53344
rect 27946 53279 28262 53280
rect 37946 53344 38262 53345
rect 37946 53280 37952 53344
rect 38016 53280 38032 53344
rect 38096 53280 38112 53344
rect 38176 53280 38192 53344
rect 38256 53280 38262 53344
rect 37946 53279 38262 53280
rect 47946 53344 48262 53345
rect 47946 53280 47952 53344
rect 48016 53280 48032 53344
rect 48096 53280 48112 53344
rect 48176 53280 48192 53344
rect 48256 53280 48262 53344
rect 47946 53279 48262 53280
rect 0 53002 800 53032
rect 3601 53002 3667 53005
rect 0 53000 3667 53002
rect 0 52944 3606 53000
rect 3662 52944 3667 53000
rect 0 52942 3667 52944
rect 0 52912 800 52942
rect 3601 52939 3667 52942
rect 2946 52800 3262 52801
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 32946 52800 33262 52801
rect 32946 52736 32952 52800
rect 33016 52736 33032 52800
rect 33096 52736 33112 52800
rect 33176 52736 33192 52800
rect 33256 52736 33262 52800
rect 32946 52735 33262 52736
rect 42946 52800 43262 52801
rect 42946 52736 42952 52800
rect 43016 52736 43032 52800
rect 43096 52736 43112 52800
rect 43176 52736 43192 52800
rect 43256 52736 43262 52800
rect 42946 52735 43262 52736
rect 49049 52458 49115 52461
rect 50200 52458 51000 52488
rect 49049 52456 51000 52458
rect 49049 52400 49054 52456
rect 49110 52400 51000 52456
rect 49049 52398 51000 52400
rect 49049 52395 49115 52398
rect 50200 52368 51000 52398
rect 7946 52256 8262 52257
rect 0 52186 800 52216
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 27946 52256 28262 52257
rect 27946 52192 27952 52256
rect 28016 52192 28032 52256
rect 28096 52192 28112 52256
rect 28176 52192 28192 52256
rect 28256 52192 28262 52256
rect 27946 52191 28262 52192
rect 37946 52256 38262 52257
rect 37946 52192 37952 52256
rect 38016 52192 38032 52256
rect 38096 52192 38112 52256
rect 38176 52192 38192 52256
rect 38256 52192 38262 52256
rect 37946 52191 38262 52192
rect 47946 52256 48262 52257
rect 47946 52192 47952 52256
rect 48016 52192 48032 52256
rect 48096 52192 48112 52256
rect 48176 52192 48192 52256
rect 48256 52192 48262 52256
rect 47946 52191 48262 52192
rect 3325 52186 3391 52189
rect 0 52184 3391 52186
rect 0 52128 3330 52184
rect 3386 52128 3391 52184
rect 0 52126 3391 52128
rect 0 52096 800 52126
rect 3325 52123 3391 52126
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 32946 51712 33262 51713
rect 32946 51648 32952 51712
rect 33016 51648 33032 51712
rect 33096 51648 33112 51712
rect 33176 51648 33192 51712
rect 33256 51648 33262 51712
rect 32946 51647 33262 51648
rect 42946 51712 43262 51713
rect 42946 51648 42952 51712
rect 43016 51648 43032 51712
rect 43096 51648 43112 51712
rect 43176 51648 43192 51712
rect 43256 51648 43262 51712
rect 42946 51647 43262 51648
rect 0 51370 800 51400
rect 1301 51370 1367 51373
rect 0 51368 1367 51370
rect 0 51312 1306 51368
rect 1362 51312 1367 51368
rect 0 51310 1367 51312
rect 0 51280 800 51310
rect 1301 51307 1367 51310
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 27946 51168 28262 51169
rect 27946 51104 27952 51168
rect 28016 51104 28032 51168
rect 28096 51104 28112 51168
rect 28176 51104 28192 51168
rect 28256 51104 28262 51168
rect 27946 51103 28262 51104
rect 37946 51168 38262 51169
rect 37946 51104 37952 51168
rect 38016 51104 38032 51168
rect 38096 51104 38112 51168
rect 38176 51104 38192 51168
rect 38256 51104 38262 51168
rect 37946 51103 38262 51104
rect 47946 51168 48262 51169
rect 47946 51104 47952 51168
rect 48016 51104 48032 51168
rect 48096 51104 48112 51168
rect 48176 51104 48192 51168
rect 48256 51104 48262 51168
rect 47946 51103 48262 51104
rect 2946 50624 3262 50625
rect 0 50554 800 50584
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 32946 50624 33262 50625
rect 32946 50560 32952 50624
rect 33016 50560 33032 50624
rect 33096 50560 33112 50624
rect 33176 50560 33192 50624
rect 33256 50560 33262 50624
rect 32946 50559 33262 50560
rect 42946 50624 43262 50625
rect 42946 50560 42952 50624
rect 43016 50560 43032 50624
rect 43096 50560 43112 50624
rect 43176 50560 43192 50624
rect 43256 50560 43262 50624
rect 42946 50559 43262 50560
rect 1301 50554 1367 50557
rect 0 50552 1367 50554
rect 0 50496 1306 50552
rect 1362 50496 1367 50552
rect 0 50494 1367 50496
rect 0 50464 800 50494
rect 1301 50491 1367 50494
rect 49049 50282 49115 50285
rect 50200 50282 51000 50312
rect 49049 50280 51000 50282
rect 49049 50224 49054 50280
rect 49110 50224 51000 50280
rect 49049 50222 51000 50224
rect 49049 50219 49115 50222
rect 50200 50192 51000 50222
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 27946 50080 28262 50081
rect 27946 50016 27952 50080
rect 28016 50016 28032 50080
rect 28096 50016 28112 50080
rect 28176 50016 28192 50080
rect 28256 50016 28262 50080
rect 27946 50015 28262 50016
rect 37946 50080 38262 50081
rect 37946 50016 37952 50080
rect 38016 50016 38032 50080
rect 38096 50016 38112 50080
rect 38176 50016 38192 50080
rect 38256 50016 38262 50080
rect 37946 50015 38262 50016
rect 47946 50080 48262 50081
rect 47946 50016 47952 50080
rect 48016 50016 48032 50080
rect 48096 50016 48112 50080
rect 48176 50016 48192 50080
rect 48256 50016 48262 50080
rect 47946 50015 48262 50016
rect 0 49738 800 49768
rect 1301 49738 1367 49741
rect 0 49736 1367 49738
rect 0 49680 1306 49736
rect 1362 49680 1367 49736
rect 0 49678 1367 49680
rect 0 49648 800 49678
rect 1301 49675 1367 49678
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 32946 49536 33262 49537
rect 32946 49472 32952 49536
rect 33016 49472 33032 49536
rect 33096 49472 33112 49536
rect 33176 49472 33192 49536
rect 33256 49472 33262 49536
rect 32946 49471 33262 49472
rect 42946 49536 43262 49537
rect 42946 49472 42952 49536
rect 43016 49472 43032 49536
rect 43096 49472 43112 49536
rect 43176 49472 43192 49536
rect 43256 49472 43262 49536
rect 42946 49471 43262 49472
rect 7946 48992 8262 48993
rect 0 48922 800 48952
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 27946 48992 28262 48993
rect 27946 48928 27952 48992
rect 28016 48928 28032 48992
rect 28096 48928 28112 48992
rect 28176 48928 28192 48992
rect 28256 48928 28262 48992
rect 27946 48927 28262 48928
rect 37946 48992 38262 48993
rect 37946 48928 37952 48992
rect 38016 48928 38032 48992
rect 38096 48928 38112 48992
rect 38176 48928 38192 48992
rect 38256 48928 38262 48992
rect 37946 48927 38262 48928
rect 47946 48992 48262 48993
rect 47946 48928 47952 48992
rect 48016 48928 48032 48992
rect 48096 48928 48112 48992
rect 48176 48928 48192 48992
rect 48256 48928 48262 48992
rect 47946 48927 48262 48928
rect 1301 48922 1367 48925
rect 0 48920 1367 48922
rect 0 48864 1306 48920
rect 1362 48864 1367 48920
rect 0 48862 1367 48864
rect 0 48832 800 48862
rect 1301 48859 1367 48862
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 32946 48448 33262 48449
rect 32946 48384 32952 48448
rect 33016 48384 33032 48448
rect 33096 48384 33112 48448
rect 33176 48384 33192 48448
rect 33256 48384 33262 48448
rect 32946 48383 33262 48384
rect 42946 48448 43262 48449
rect 42946 48384 42952 48448
rect 43016 48384 43032 48448
rect 43096 48384 43112 48448
rect 43176 48384 43192 48448
rect 43256 48384 43262 48448
rect 42946 48383 43262 48384
rect 0 48106 800 48136
rect 1301 48106 1367 48109
rect 0 48104 1367 48106
rect 0 48048 1306 48104
rect 1362 48048 1367 48104
rect 0 48046 1367 48048
rect 0 48016 800 48046
rect 1301 48043 1367 48046
rect 17861 48106 17927 48109
rect 18413 48106 18479 48109
rect 17861 48104 18479 48106
rect 17861 48048 17866 48104
rect 17922 48048 18418 48104
rect 18474 48048 18479 48104
rect 17861 48046 18479 48048
rect 17861 48043 17927 48046
rect 18413 48043 18479 48046
rect 48957 48106 49023 48109
rect 50200 48106 51000 48136
rect 48957 48104 51000 48106
rect 48957 48048 48962 48104
rect 49018 48048 51000 48104
rect 48957 48046 51000 48048
rect 48957 48043 49023 48046
rect 50200 48016 51000 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 27946 47904 28262 47905
rect 27946 47840 27952 47904
rect 28016 47840 28032 47904
rect 28096 47840 28112 47904
rect 28176 47840 28192 47904
rect 28256 47840 28262 47904
rect 27946 47839 28262 47840
rect 37946 47904 38262 47905
rect 37946 47840 37952 47904
rect 38016 47840 38032 47904
rect 38096 47840 38112 47904
rect 38176 47840 38192 47904
rect 38256 47840 38262 47904
rect 37946 47839 38262 47840
rect 47946 47904 48262 47905
rect 47946 47840 47952 47904
rect 48016 47840 48032 47904
rect 48096 47840 48112 47904
rect 48176 47840 48192 47904
rect 48256 47840 48262 47904
rect 47946 47839 48262 47840
rect 2946 47360 3262 47361
rect 0 47290 800 47320
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 32946 47360 33262 47361
rect 32946 47296 32952 47360
rect 33016 47296 33032 47360
rect 33096 47296 33112 47360
rect 33176 47296 33192 47360
rect 33256 47296 33262 47360
rect 32946 47295 33262 47296
rect 42946 47360 43262 47361
rect 42946 47296 42952 47360
rect 43016 47296 43032 47360
rect 43096 47296 43112 47360
rect 43176 47296 43192 47360
rect 43256 47296 43262 47360
rect 42946 47295 43262 47296
rect 1301 47290 1367 47293
rect 0 47288 1367 47290
rect 0 47232 1306 47288
rect 1362 47232 1367 47288
rect 0 47230 1367 47232
rect 0 47200 800 47230
rect 1301 47227 1367 47230
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 27946 46816 28262 46817
rect 27946 46752 27952 46816
rect 28016 46752 28032 46816
rect 28096 46752 28112 46816
rect 28176 46752 28192 46816
rect 28256 46752 28262 46816
rect 27946 46751 28262 46752
rect 37946 46816 38262 46817
rect 37946 46752 37952 46816
rect 38016 46752 38032 46816
rect 38096 46752 38112 46816
rect 38176 46752 38192 46816
rect 38256 46752 38262 46816
rect 37946 46751 38262 46752
rect 47946 46816 48262 46817
rect 47946 46752 47952 46816
rect 48016 46752 48032 46816
rect 48096 46752 48112 46816
rect 48176 46752 48192 46816
rect 48256 46752 48262 46816
rect 47946 46751 48262 46752
rect 0 46474 800 46504
rect 1301 46474 1367 46477
rect 0 46472 1367 46474
rect 0 46416 1306 46472
rect 1362 46416 1367 46472
rect 0 46414 1367 46416
rect 0 46384 800 46414
rect 1301 46411 1367 46414
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 32946 46272 33262 46273
rect 32946 46208 32952 46272
rect 33016 46208 33032 46272
rect 33096 46208 33112 46272
rect 33176 46208 33192 46272
rect 33256 46208 33262 46272
rect 32946 46207 33262 46208
rect 42946 46272 43262 46273
rect 42946 46208 42952 46272
rect 43016 46208 43032 46272
rect 43096 46208 43112 46272
rect 43176 46208 43192 46272
rect 43256 46208 43262 46272
rect 42946 46207 43262 46208
rect 49141 45930 49207 45933
rect 50200 45930 51000 45960
rect 49141 45928 51000 45930
rect 49141 45872 49146 45928
rect 49202 45872 51000 45928
rect 49141 45870 51000 45872
rect 49141 45867 49207 45870
rect 50200 45840 51000 45870
rect 7946 45728 8262 45729
rect 0 45658 800 45688
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 27946 45728 28262 45729
rect 27946 45664 27952 45728
rect 28016 45664 28032 45728
rect 28096 45664 28112 45728
rect 28176 45664 28192 45728
rect 28256 45664 28262 45728
rect 27946 45663 28262 45664
rect 37946 45728 38262 45729
rect 37946 45664 37952 45728
rect 38016 45664 38032 45728
rect 38096 45664 38112 45728
rect 38176 45664 38192 45728
rect 38256 45664 38262 45728
rect 37946 45663 38262 45664
rect 47946 45728 48262 45729
rect 47946 45664 47952 45728
rect 48016 45664 48032 45728
rect 48096 45664 48112 45728
rect 48176 45664 48192 45728
rect 48256 45664 48262 45728
rect 47946 45663 48262 45664
rect 1301 45658 1367 45661
rect 0 45656 1367 45658
rect 0 45600 1306 45656
rect 1362 45600 1367 45656
rect 0 45598 1367 45600
rect 0 45568 800 45598
rect 1301 45595 1367 45598
rect 3509 45522 3575 45525
rect 15929 45522 15995 45525
rect 20437 45522 20503 45525
rect 23749 45522 23815 45525
rect 3509 45520 23815 45522
rect 3509 45464 3514 45520
rect 3570 45464 15934 45520
rect 15990 45464 20442 45520
rect 20498 45464 23754 45520
rect 23810 45464 23815 45520
rect 3509 45462 23815 45464
rect 3509 45459 3575 45462
rect 15929 45459 15995 45462
rect 20437 45459 20503 45462
rect 23749 45459 23815 45462
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 32946 45184 33262 45185
rect 32946 45120 32952 45184
rect 33016 45120 33032 45184
rect 33096 45120 33112 45184
rect 33176 45120 33192 45184
rect 33256 45120 33262 45184
rect 32946 45119 33262 45120
rect 42946 45184 43262 45185
rect 42946 45120 42952 45184
rect 43016 45120 43032 45184
rect 43096 45120 43112 45184
rect 43176 45120 43192 45184
rect 43256 45120 43262 45184
rect 42946 45119 43262 45120
rect 0 44842 800 44872
rect 1301 44842 1367 44845
rect 0 44840 1367 44842
rect 0 44784 1306 44840
rect 1362 44784 1367 44840
rect 0 44782 1367 44784
rect 0 44752 800 44782
rect 1301 44779 1367 44782
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 27946 44640 28262 44641
rect 27946 44576 27952 44640
rect 28016 44576 28032 44640
rect 28096 44576 28112 44640
rect 28176 44576 28192 44640
rect 28256 44576 28262 44640
rect 27946 44575 28262 44576
rect 37946 44640 38262 44641
rect 37946 44576 37952 44640
rect 38016 44576 38032 44640
rect 38096 44576 38112 44640
rect 38176 44576 38192 44640
rect 38256 44576 38262 44640
rect 37946 44575 38262 44576
rect 47946 44640 48262 44641
rect 47946 44576 47952 44640
rect 48016 44576 48032 44640
rect 48096 44576 48112 44640
rect 48176 44576 48192 44640
rect 48256 44576 48262 44640
rect 47946 44575 48262 44576
rect 2946 44096 3262 44097
rect 0 44026 800 44056
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 32946 44096 33262 44097
rect 32946 44032 32952 44096
rect 33016 44032 33032 44096
rect 33096 44032 33112 44096
rect 33176 44032 33192 44096
rect 33256 44032 33262 44096
rect 32946 44031 33262 44032
rect 42946 44096 43262 44097
rect 42946 44032 42952 44096
rect 43016 44032 43032 44096
rect 43096 44032 43112 44096
rect 43176 44032 43192 44096
rect 43256 44032 43262 44096
rect 42946 44031 43262 44032
rect 2037 44026 2103 44029
rect 0 44024 2103 44026
rect 0 43968 2042 44024
rect 2098 43968 2103 44024
rect 0 43966 2103 43968
rect 0 43936 800 43966
rect 2037 43963 2103 43966
rect 7946 43552 8262 43553
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 27946 43552 28262 43553
rect 27946 43488 27952 43552
rect 28016 43488 28032 43552
rect 28096 43488 28112 43552
rect 28176 43488 28192 43552
rect 28256 43488 28262 43552
rect 27946 43487 28262 43488
rect 37946 43552 38262 43553
rect 37946 43488 37952 43552
rect 38016 43488 38032 43552
rect 38096 43488 38112 43552
rect 38176 43488 38192 43552
rect 38256 43488 38262 43552
rect 37946 43487 38262 43488
rect 47946 43552 48262 43553
rect 47946 43488 47952 43552
rect 48016 43488 48032 43552
rect 48096 43488 48112 43552
rect 48176 43488 48192 43552
rect 48256 43488 48262 43552
rect 47946 43487 48262 43488
rect 29821 43346 29887 43349
rect 12390 43344 29887 43346
rect 12390 43288 29826 43344
rect 29882 43288 29887 43344
rect 12390 43286 29887 43288
rect 0 43210 800 43240
rect 1301 43210 1367 43213
rect 9213 43212 9279 43213
rect 9213 43210 9260 43212
rect 0 43208 1367 43210
rect 0 43152 1306 43208
rect 1362 43152 1367 43208
rect 0 43150 1367 43152
rect 9168 43208 9260 43210
rect 9324 43210 9330 43212
rect 12390 43210 12450 43286
rect 29821 43283 29887 43286
rect 9168 43152 9218 43208
rect 9168 43150 9260 43152
rect 0 43120 800 43150
rect 1301 43147 1367 43150
rect 9213 43148 9260 43150
rect 9324 43150 12450 43210
rect 9324 43148 9330 43150
rect 9213 43147 9279 43148
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 32946 43008 33262 43009
rect 32946 42944 32952 43008
rect 33016 42944 33032 43008
rect 33096 42944 33112 43008
rect 33176 42944 33192 43008
rect 33256 42944 33262 43008
rect 32946 42943 33262 42944
rect 42946 43008 43262 43009
rect 42946 42944 42952 43008
rect 43016 42944 43032 43008
rect 43096 42944 43112 43008
rect 43176 42944 43192 43008
rect 43256 42944 43262 43008
rect 42946 42943 43262 42944
rect 20713 42802 20779 42805
rect 40217 42802 40283 42805
rect 20713 42800 40283 42802
rect 20713 42744 20718 42800
rect 20774 42744 40222 42800
rect 40278 42744 40283 42800
rect 20713 42742 40283 42744
rect 20713 42739 20779 42742
rect 40217 42739 40283 42742
rect 18689 42666 18755 42669
rect 38929 42666 38995 42669
rect 18689 42664 38995 42666
rect 18689 42608 18694 42664
rect 18750 42608 38934 42664
rect 38990 42608 38995 42664
rect 18689 42606 38995 42608
rect 18689 42603 18755 42606
rect 38929 42603 38995 42606
rect 7946 42464 8262 42465
rect 0 42394 800 42424
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 27946 42464 28262 42465
rect 27946 42400 27952 42464
rect 28016 42400 28032 42464
rect 28096 42400 28112 42464
rect 28176 42400 28192 42464
rect 28256 42400 28262 42464
rect 27946 42399 28262 42400
rect 37946 42464 38262 42465
rect 37946 42400 37952 42464
rect 38016 42400 38032 42464
rect 38096 42400 38112 42464
rect 38176 42400 38192 42464
rect 38256 42400 38262 42464
rect 37946 42399 38262 42400
rect 47946 42464 48262 42465
rect 47946 42400 47952 42464
rect 48016 42400 48032 42464
rect 48096 42400 48112 42464
rect 48176 42400 48192 42464
rect 48256 42400 48262 42464
rect 47946 42399 48262 42400
rect 1301 42394 1367 42397
rect 0 42392 1367 42394
rect 0 42336 1306 42392
rect 1362 42336 1367 42392
rect 0 42334 1367 42336
rect 0 42304 800 42334
rect 1301 42331 1367 42334
rect 18781 41988 18847 41989
rect 18781 41984 18828 41988
rect 18892 41986 18898 41988
rect 18781 41928 18786 41984
rect 18781 41924 18828 41928
rect 18892 41926 18938 41986
rect 18892 41924 18898 41926
rect 18781 41923 18847 41924
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 32946 41920 33262 41921
rect 32946 41856 32952 41920
rect 33016 41856 33032 41920
rect 33096 41856 33112 41920
rect 33176 41856 33192 41920
rect 33256 41856 33262 41920
rect 32946 41855 33262 41856
rect 42946 41920 43262 41921
rect 42946 41856 42952 41920
rect 43016 41856 43032 41920
rect 43096 41856 43112 41920
rect 43176 41856 43192 41920
rect 43256 41856 43262 41920
rect 42946 41855 43262 41856
rect 14365 41850 14431 41853
rect 17493 41850 17559 41853
rect 14365 41848 17559 41850
rect 14365 41792 14370 41848
rect 14426 41792 17498 41848
rect 17554 41792 17559 41848
rect 14365 41790 17559 41792
rect 14365 41787 14431 41790
rect 17493 41787 17559 41790
rect 14733 41714 14799 41717
rect 20989 41714 21055 41717
rect 14733 41712 21055 41714
rect 14733 41656 14738 41712
rect 14794 41656 20994 41712
rect 21050 41656 21055 41712
rect 14733 41654 21055 41656
rect 14733 41651 14799 41654
rect 20989 41651 21055 41654
rect 0 41578 800 41608
rect 1301 41578 1367 41581
rect 0 41576 1367 41578
rect 0 41520 1306 41576
rect 1362 41520 1367 41576
rect 0 41518 1367 41520
rect 0 41488 800 41518
rect 1301 41515 1367 41518
rect 18229 41578 18295 41581
rect 18505 41578 18571 41581
rect 18229 41576 18571 41578
rect 18229 41520 18234 41576
rect 18290 41520 18510 41576
rect 18566 41520 18571 41576
rect 18229 41518 18571 41520
rect 18229 41515 18295 41518
rect 18505 41515 18571 41518
rect 19609 41442 19675 41445
rect 23749 41442 23815 41445
rect 19609 41440 23815 41442
rect 19609 41384 19614 41440
rect 19670 41384 23754 41440
rect 23810 41384 23815 41440
rect 19609 41382 23815 41384
rect 19609 41379 19675 41382
rect 23749 41379 23815 41382
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 27946 41376 28262 41377
rect 27946 41312 27952 41376
rect 28016 41312 28032 41376
rect 28096 41312 28112 41376
rect 28176 41312 28192 41376
rect 28256 41312 28262 41376
rect 27946 41311 28262 41312
rect 37946 41376 38262 41377
rect 37946 41312 37952 41376
rect 38016 41312 38032 41376
rect 38096 41312 38112 41376
rect 38176 41312 38192 41376
rect 38256 41312 38262 41376
rect 37946 41311 38262 41312
rect 47946 41376 48262 41377
rect 47946 41312 47952 41376
rect 48016 41312 48032 41376
rect 48096 41312 48112 41376
rect 48176 41312 48192 41376
rect 48256 41312 48262 41376
rect 47946 41311 48262 41312
rect 12065 41170 12131 41173
rect 12617 41170 12683 41173
rect 34237 41170 34303 41173
rect 12065 41168 34303 41170
rect 12065 41112 12070 41168
rect 12126 41112 12622 41168
rect 12678 41112 34242 41168
rect 34298 41112 34303 41168
rect 12065 41110 34303 41112
rect 12065 41107 12131 41110
rect 12617 41107 12683 41110
rect 34237 41107 34303 41110
rect 10777 41034 10843 41037
rect 14917 41034 14983 41037
rect 10777 41032 14983 41034
rect 10777 40976 10782 41032
rect 10838 40976 14922 41032
rect 14978 40976 14983 41032
rect 10777 40974 14983 40976
rect 10777 40971 10843 40974
rect 14917 40971 14983 40974
rect 10685 40900 10751 40901
rect 10685 40898 10732 40900
rect 10640 40896 10732 40898
rect 10640 40840 10690 40896
rect 10640 40838 10732 40840
rect 10685 40836 10732 40838
rect 10796 40836 10802 40900
rect 10685 40835 10751 40836
rect 2946 40832 3262 40833
rect 0 40762 800 40792
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 32946 40832 33262 40833
rect 32946 40768 32952 40832
rect 33016 40768 33032 40832
rect 33096 40768 33112 40832
rect 33176 40768 33192 40832
rect 33256 40768 33262 40832
rect 32946 40767 33262 40768
rect 42946 40832 43262 40833
rect 42946 40768 42952 40832
rect 43016 40768 43032 40832
rect 43096 40768 43112 40832
rect 43176 40768 43192 40832
rect 43256 40768 43262 40832
rect 42946 40767 43262 40768
rect 1301 40762 1367 40765
rect 0 40760 1367 40762
rect 0 40704 1306 40760
rect 1362 40704 1367 40760
rect 0 40702 1367 40704
rect 0 40672 800 40702
rect 1301 40699 1367 40702
rect 12249 40626 12315 40629
rect 12985 40626 13051 40629
rect 12249 40624 13051 40626
rect 12249 40568 12254 40624
rect 12310 40568 12990 40624
rect 13046 40568 13051 40624
rect 12249 40566 13051 40568
rect 12249 40563 12315 40566
rect 12985 40563 13051 40566
rect 9857 40490 9923 40493
rect 18505 40490 18571 40493
rect 9857 40488 18571 40490
rect 9857 40432 9862 40488
rect 9918 40432 18510 40488
rect 18566 40432 18571 40488
rect 9857 40430 18571 40432
rect 9857 40427 9923 40430
rect 18505 40427 18571 40430
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 27946 40288 28262 40289
rect 27946 40224 27952 40288
rect 28016 40224 28032 40288
rect 28096 40224 28112 40288
rect 28176 40224 28192 40288
rect 28256 40224 28262 40288
rect 27946 40223 28262 40224
rect 37946 40288 38262 40289
rect 37946 40224 37952 40288
rect 38016 40224 38032 40288
rect 38096 40224 38112 40288
rect 38176 40224 38192 40288
rect 38256 40224 38262 40288
rect 37946 40223 38262 40224
rect 47946 40288 48262 40289
rect 47946 40224 47952 40288
rect 48016 40224 48032 40288
rect 48096 40224 48112 40288
rect 48176 40224 48192 40288
rect 48256 40224 48262 40288
rect 47946 40223 48262 40224
rect 12157 40218 12223 40221
rect 12341 40218 12407 40221
rect 12157 40216 12407 40218
rect 12157 40160 12162 40216
rect 12218 40160 12346 40216
rect 12402 40160 12407 40216
rect 12157 40158 12407 40160
rect 12157 40155 12223 40158
rect 12341 40155 12407 40158
rect 10961 40082 11027 40085
rect 18873 40082 18939 40085
rect 10961 40080 18939 40082
rect 10961 40024 10966 40080
rect 11022 40024 18878 40080
rect 18934 40024 18939 40080
rect 10961 40022 18939 40024
rect 10961 40019 11027 40022
rect 18873 40019 18939 40022
rect 0 39946 800 39976
rect 2037 39946 2103 39949
rect 0 39944 2103 39946
rect 0 39888 2042 39944
rect 2098 39888 2103 39944
rect 0 39886 2103 39888
rect 0 39856 800 39886
rect 2037 39883 2103 39886
rect 12249 39946 12315 39949
rect 12433 39946 12499 39949
rect 12249 39944 12499 39946
rect 12249 39888 12254 39944
rect 12310 39888 12438 39944
rect 12494 39888 12499 39944
rect 12249 39886 12499 39888
rect 12249 39883 12315 39886
rect 12433 39883 12499 39886
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 32946 39744 33262 39745
rect 32946 39680 32952 39744
rect 33016 39680 33032 39744
rect 33096 39680 33112 39744
rect 33176 39680 33192 39744
rect 33256 39680 33262 39744
rect 32946 39679 33262 39680
rect 42946 39744 43262 39745
rect 42946 39680 42952 39744
rect 43016 39680 43032 39744
rect 43096 39680 43112 39744
rect 43176 39680 43192 39744
rect 43256 39680 43262 39744
rect 42946 39679 43262 39680
rect 10501 39538 10567 39541
rect 12893 39538 12959 39541
rect 10501 39536 12959 39538
rect 10501 39480 10506 39536
rect 10562 39480 12898 39536
rect 12954 39480 12959 39536
rect 10501 39478 12959 39480
rect 10501 39475 10567 39478
rect 12893 39475 12959 39478
rect 13077 39538 13143 39541
rect 18689 39538 18755 39541
rect 13077 39536 18755 39538
rect 13077 39480 13082 39536
rect 13138 39480 18694 39536
rect 18750 39480 18755 39536
rect 13077 39478 18755 39480
rect 13077 39475 13143 39478
rect 18689 39475 18755 39478
rect 12525 39266 12591 39269
rect 13537 39266 13603 39269
rect 12525 39264 13603 39266
rect 12525 39208 12530 39264
rect 12586 39208 13542 39264
rect 13598 39208 13603 39264
rect 12525 39206 13603 39208
rect 12525 39203 12591 39206
rect 13537 39203 13603 39206
rect 7946 39200 8262 39201
rect 0 39130 800 39160
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 27946 39200 28262 39201
rect 27946 39136 27952 39200
rect 28016 39136 28032 39200
rect 28096 39136 28112 39200
rect 28176 39136 28192 39200
rect 28256 39136 28262 39200
rect 27946 39135 28262 39136
rect 37946 39200 38262 39201
rect 37946 39136 37952 39200
rect 38016 39136 38032 39200
rect 38096 39136 38112 39200
rect 38176 39136 38192 39200
rect 38256 39136 38262 39200
rect 37946 39135 38262 39136
rect 47946 39200 48262 39201
rect 47946 39136 47952 39200
rect 48016 39136 48032 39200
rect 48096 39136 48112 39200
rect 48176 39136 48192 39200
rect 48256 39136 48262 39200
rect 47946 39135 48262 39136
rect 1301 39130 1367 39133
rect 0 39128 1367 39130
rect 0 39072 1306 39128
rect 1362 39072 1367 39128
rect 0 39070 1367 39072
rect 0 39040 800 39070
rect 1301 39067 1367 39070
rect 12985 39130 13051 39133
rect 13629 39130 13695 39133
rect 12985 39128 13695 39130
rect 12985 39072 12990 39128
rect 13046 39072 13634 39128
rect 13690 39072 13695 39128
rect 12985 39070 13695 39072
rect 12985 39067 13051 39070
rect 13629 39067 13695 39070
rect 12065 38994 12131 38997
rect 18229 38994 18295 38997
rect 12065 38992 18295 38994
rect 12065 38936 12070 38992
rect 12126 38936 18234 38992
rect 18290 38936 18295 38992
rect 12065 38934 18295 38936
rect 12065 38931 12131 38934
rect 18229 38931 18295 38934
rect 11881 38858 11947 38861
rect 14181 38858 14247 38861
rect 11881 38856 14247 38858
rect 11881 38800 11886 38856
rect 11942 38800 14186 38856
rect 14242 38800 14247 38856
rect 11881 38798 14247 38800
rect 11881 38795 11947 38798
rect 14181 38795 14247 38798
rect 9121 38722 9187 38725
rect 12525 38722 12591 38725
rect 9121 38720 12591 38722
rect 9121 38664 9126 38720
rect 9182 38664 12530 38720
rect 12586 38664 12591 38720
rect 9121 38662 12591 38664
rect 9121 38659 9187 38662
rect 12525 38659 12591 38662
rect 19425 38722 19491 38725
rect 21357 38722 21423 38725
rect 19425 38720 21423 38722
rect 19425 38664 19430 38720
rect 19486 38664 21362 38720
rect 21418 38664 21423 38720
rect 19425 38662 21423 38664
rect 19425 38659 19491 38662
rect 21357 38659 21423 38662
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 32946 38656 33262 38657
rect 32946 38592 32952 38656
rect 33016 38592 33032 38656
rect 33096 38592 33112 38656
rect 33176 38592 33192 38656
rect 33256 38592 33262 38656
rect 32946 38591 33262 38592
rect 42946 38656 43262 38657
rect 42946 38592 42952 38656
rect 43016 38592 43032 38656
rect 43096 38592 43112 38656
rect 43176 38592 43192 38656
rect 43256 38592 43262 38656
rect 42946 38591 43262 38592
rect 0 38314 800 38344
rect 1301 38314 1367 38317
rect 0 38312 1367 38314
rect 0 38256 1306 38312
rect 1362 38256 1367 38312
rect 0 38254 1367 38256
rect 0 38224 800 38254
rect 1301 38251 1367 38254
rect 10869 38180 10935 38181
rect 10869 38178 10916 38180
rect 10824 38176 10916 38178
rect 10824 38120 10874 38176
rect 10824 38118 10916 38120
rect 10869 38116 10916 38118
rect 10980 38116 10986 38180
rect 15377 38178 15443 38181
rect 15929 38178 15995 38181
rect 17217 38178 17283 38181
rect 17769 38178 17835 38181
rect 15377 38176 17835 38178
rect 15377 38120 15382 38176
rect 15438 38120 15934 38176
rect 15990 38120 17222 38176
rect 17278 38120 17774 38176
rect 17830 38120 17835 38176
rect 15377 38118 17835 38120
rect 10869 38115 10935 38116
rect 15377 38115 15443 38118
rect 15929 38115 15995 38118
rect 17217 38115 17283 38118
rect 17769 38115 17835 38118
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 27946 38112 28262 38113
rect 27946 38048 27952 38112
rect 28016 38048 28032 38112
rect 28096 38048 28112 38112
rect 28176 38048 28192 38112
rect 28256 38048 28262 38112
rect 27946 38047 28262 38048
rect 37946 38112 38262 38113
rect 37946 38048 37952 38112
rect 38016 38048 38032 38112
rect 38096 38048 38112 38112
rect 38176 38048 38192 38112
rect 38256 38048 38262 38112
rect 37946 38047 38262 38048
rect 47946 38112 48262 38113
rect 47946 38048 47952 38112
rect 48016 38048 48032 38112
rect 48096 38048 48112 38112
rect 48176 38048 48192 38112
rect 48256 38048 48262 38112
rect 47946 38047 48262 38048
rect 13813 38042 13879 38045
rect 16941 38042 17007 38045
rect 13813 38040 17007 38042
rect 13813 37984 13818 38040
rect 13874 37984 16946 38040
rect 17002 37984 17007 38040
rect 13813 37982 17007 37984
rect 13813 37979 13879 37982
rect 16941 37979 17007 37982
rect 23473 37906 23539 37909
rect 18462 37904 23539 37906
rect 18462 37848 23478 37904
rect 23534 37848 23539 37904
rect 18462 37846 23539 37848
rect 18462 37773 18522 37846
rect 23473 37843 23539 37846
rect 12985 37770 13051 37773
rect 18413 37770 18522 37773
rect 12985 37768 18522 37770
rect 12985 37712 12990 37768
rect 13046 37712 18418 37768
rect 18474 37712 18522 37768
rect 12985 37710 18522 37712
rect 12985 37707 13051 37710
rect 18413 37707 18479 37710
rect 2946 37568 3262 37569
rect 0 37498 800 37528
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 32946 37568 33262 37569
rect 32946 37504 32952 37568
rect 33016 37504 33032 37568
rect 33096 37504 33112 37568
rect 33176 37504 33192 37568
rect 33256 37504 33262 37568
rect 32946 37503 33262 37504
rect 42946 37568 43262 37569
rect 42946 37504 42952 37568
rect 43016 37504 43032 37568
rect 43096 37504 43112 37568
rect 43176 37504 43192 37568
rect 43256 37504 43262 37568
rect 42946 37503 43262 37504
rect 1301 37498 1367 37501
rect 0 37496 1367 37498
rect 0 37440 1306 37496
rect 1362 37440 1367 37496
rect 0 37438 1367 37440
rect 0 37408 800 37438
rect 1301 37435 1367 37438
rect 7373 37498 7439 37501
rect 9305 37498 9371 37501
rect 9673 37498 9739 37501
rect 7373 37496 9739 37498
rect 7373 37440 7378 37496
rect 7434 37440 9310 37496
rect 9366 37440 9678 37496
rect 9734 37440 9739 37496
rect 7373 37438 9739 37440
rect 7373 37435 7439 37438
rect 9305 37435 9371 37438
rect 9673 37435 9739 37438
rect 6269 37362 6335 37365
rect 9029 37362 9095 37365
rect 6269 37360 9095 37362
rect 6269 37304 6274 37360
rect 6330 37304 9034 37360
rect 9090 37304 9095 37360
rect 6269 37302 9095 37304
rect 6269 37299 6335 37302
rect 9029 37299 9095 37302
rect 11053 37228 11119 37229
rect 11053 37226 11100 37228
rect 11008 37224 11100 37226
rect 11008 37168 11058 37224
rect 11008 37166 11100 37168
rect 11053 37164 11100 37166
rect 11164 37164 11170 37228
rect 17769 37226 17835 37229
rect 18781 37226 18847 37229
rect 17769 37224 18847 37226
rect 17769 37168 17774 37224
rect 17830 37168 18786 37224
rect 18842 37168 18847 37224
rect 17769 37166 18847 37168
rect 11053 37163 11119 37164
rect 17769 37163 17835 37166
rect 18781 37163 18847 37166
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 27946 37024 28262 37025
rect 27946 36960 27952 37024
rect 28016 36960 28032 37024
rect 28096 36960 28112 37024
rect 28176 36960 28192 37024
rect 28256 36960 28262 37024
rect 27946 36959 28262 36960
rect 37946 37024 38262 37025
rect 37946 36960 37952 37024
rect 38016 36960 38032 37024
rect 38096 36960 38112 37024
rect 38176 36960 38192 37024
rect 38256 36960 38262 37024
rect 37946 36959 38262 36960
rect 47946 37024 48262 37025
rect 47946 36960 47952 37024
rect 48016 36960 48032 37024
rect 48096 36960 48112 37024
rect 48176 36960 48192 37024
rect 48256 36960 48262 37024
rect 47946 36959 48262 36960
rect 9254 36892 9260 36956
rect 9324 36954 9330 36956
rect 9581 36954 9647 36957
rect 9324 36952 9647 36954
rect 9324 36896 9586 36952
rect 9642 36896 9647 36952
rect 9324 36894 9647 36896
rect 9324 36892 9330 36894
rect 9581 36891 9647 36894
rect 7465 36818 7531 36821
rect 12249 36818 12315 36821
rect 7465 36816 12315 36818
rect 7465 36760 7470 36816
rect 7526 36760 12254 36816
rect 12310 36760 12315 36816
rect 7465 36758 12315 36760
rect 7465 36755 7531 36758
rect 12249 36755 12315 36758
rect 0 36682 800 36712
rect 1301 36682 1367 36685
rect 0 36680 1367 36682
rect 0 36624 1306 36680
rect 1362 36624 1367 36680
rect 0 36622 1367 36624
rect 0 36592 800 36622
rect 1301 36619 1367 36622
rect 7097 36682 7163 36685
rect 7230 36682 7236 36684
rect 7097 36680 7236 36682
rect 7097 36624 7102 36680
rect 7158 36624 7236 36680
rect 7097 36622 7236 36624
rect 7097 36619 7163 36622
rect 7230 36620 7236 36622
rect 7300 36682 7306 36684
rect 8201 36682 8267 36685
rect 7300 36680 8267 36682
rect 7300 36624 8206 36680
rect 8262 36624 8267 36680
rect 7300 36622 8267 36624
rect 7300 36620 7306 36622
rect 8201 36619 8267 36622
rect 9438 36620 9444 36684
rect 9508 36682 9514 36684
rect 9581 36682 9647 36685
rect 9508 36680 9647 36682
rect 9508 36624 9586 36680
rect 9642 36624 9647 36680
rect 9508 36622 9647 36624
rect 9508 36620 9514 36622
rect 9581 36619 9647 36622
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 32946 36480 33262 36481
rect 32946 36416 32952 36480
rect 33016 36416 33032 36480
rect 33096 36416 33112 36480
rect 33176 36416 33192 36480
rect 33256 36416 33262 36480
rect 32946 36415 33262 36416
rect 42946 36480 43262 36481
rect 42946 36416 42952 36480
rect 43016 36416 43032 36480
rect 43096 36416 43112 36480
rect 43176 36416 43192 36480
rect 43256 36416 43262 36480
rect 42946 36415 43262 36416
rect 7946 35936 8262 35937
rect 0 35866 800 35896
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 27946 35936 28262 35937
rect 27946 35872 27952 35936
rect 28016 35872 28032 35936
rect 28096 35872 28112 35936
rect 28176 35872 28192 35936
rect 28256 35872 28262 35936
rect 27946 35871 28262 35872
rect 37946 35936 38262 35937
rect 37946 35872 37952 35936
rect 38016 35872 38032 35936
rect 38096 35872 38112 35936
rect 38176 35872 38192 35936
rect 38256 35872 38262 35936
rect 37946 35871 38262 35872
rect 47946 35936 48262 35937
rect 47946 35872 47952 35936
rect 48016 35872 48032 35936
rect 48096 35872 48112 35936
rect 48176 35872 48192 35936
rect 48256 35872 48262 35936
rect 47946 35871 48262 35872
rect 2773 35866 2839 35869
rect 0 35864 2839 35866
rect 0 35808 2778 35864
rect 2834 35808 2839 35864
rect 0 35806 2839 35808
rect 0 35776 800 35806
rect 2773 35803 2839 35806
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 32946 35392 33262 35393
rect 32946 35328 32952 35392
rect 33016 35328 33032 35392
rect 33096 35328 33112 35392
rect 33176 35328 33192 35392
rect 33256 35328 33262 35392
rect 32946 35327 33262 35328
rect 42946 35392 43262 35393
rect 42946 35328 42952 35392
rect 43016 35328 43032 35392
rect 43096 35328 43112 35392
rect 43176 35328 43192 35392
rect 43256 35328 43262 35392
rect 42946 35327 43262 35328
rect 0 35050 800 35080
rect 1301 35050 1367 35053
rect 0 35048 1367 35050
rect 0 34992 1306 35048
rect 1362 34992 1367 35048
rect 0 34990 1367 34992
rect 0 34960 800 34990
rect 1301 34987 1367 34990
rect 8109 35050 8175 35053
rect 13353 35050 13419 35053
rect 8109 35048 13419 35050
rect 8109 34992 8114 35048
rect 8170 34992 13358 35048
rect 13414 34992 13419 35048
rect 8109 34990 13419 34992
rect 8109 34987 8175 34990
rect 13353 34987 13419 34990
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 27946 34848 28262 34849
rect 27946 34784 27952 34848
rect 28016 34784 28032 34848
rect 28096 34784 28112 34848
rect 28176 34784 28192 34848
rect 28256 34784 28262 34848
rect 27946 34783 28262 34784
rect 37946 34848 38262 34849
rect 37946 34784 37952 34848
rect 38016 34784 38032 34848
rect 38096 34784 38112 34848
rect 38176 34784 38192 34848
rect 38256 34784 38262 34848
rect 37946 34783 38262 34784
rect 47946 34848 48262 34849
rect 47946 34784 47952 34848
rect 48016 34784 48032 34848
rect 48096 34784 48112 34848
rect 48176 34784 48192 34848
rect 48256 34784 48262 34848
rect 47946 34783 48262 34784
rect 2946 34304 3262 34305
rect 0 34234 800 34264
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 32946 34304 33262 34305
rect 32946 34240 32952 34304
rect 33016 34240 33032 34304
rect 33096 34240 33112 34304
rect 33176 34240 33192 34304
rect 33256 34240 33262 34304
rect 32946 34239 33262 34240
rect 42946 34304 43262 34305
rect 42946 34240 42952 34304
rect 43016 34240 43032 34304
rect 43096 34240 43112 34304
rect 43176 34240 43192 34304
rect 43256 34240 43262 34304
rect 42946 34239 43262 34240
rect 2037 34234 2103 34237
rect 0 34232 2103 34234
rect 0 34176 2042 34232
rect 2098 34176 2103 34232
rect 0 34174 2103 34176
rect 0 34144 800 34174
rect 2037 34171 2103 34174
rect 12617 33962 12683 33965
rect 14641 33962 14707 33965
rect 17401 33962 17467 33965
rect 17861 33962 17927 33965
rect 12617 33960 17927 33962
rect 12617 33904 12622 33960
rect 12678 33904 14646 33960
rect 14702 33904 17406 33960
rect 17462 33904 17866 33960
rect 17922 33904 17927 33960
rect 12617 33902 17927 33904
rect 12617 33899 12683 33902
rect 14641 33899 14707 33902
rect 17401 33899 17467 33902
rect 17861 33899 17927 33902
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 27946 33760 28262 33761
rect 27946 33696 27952 33760
rect 28016 33696 28032 33760
rect 28096 33696 28112 33760
rect 28176 33696 28192 33760
rect 28256 33696 28262 33760
rect 27946 33695 28262 33696
rect 37946 33760 38262 33761
rect 37946 33696 37952 33760
rect 38016 33696 38032 33760
rect 38096 33696 38112 33760
rect 38176 33696 38192 33760
rect 38256 33696 38262 33760
rect 37946 33695 38262 33696
rect 47946 33760 48262 33761
rect 47946 33696 47952 33760
rect 48016 33696 48032 33760
rect 48096 33696 48112 33760
rect 48176 33696 48192 33760
rect 48256 33696 48262 33760
rect 47946 33695 48262 33696
rect 0 33418 800 33448
rect 1301 33418 1367 33421
rect 0 33416 1367 33418
rect 0 33360 1306 33416
rect 1362 33360 1367 33416
rect 0 33358 1367 33360
rect 0 33328 800 33358
rect 1301 33355 1367 33358
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 32946 33216 33262 33217
rect 32946 33152 32952 33216
rect 33016 33152 33032 33216
rect 33096 33152 33112 33216
rect 33176 33152 33192 33216
rect 33256 33152 33262 33216
rect 32946 33151 33262 33152
rect 42946 33216 43262 33217
rect 42946 33152 42952 33216
rect 43016 33152 43032 33216
rect 43096 33152 43112 33216
rect 43176 33152 43192 33216
rect 43256 33152 43262 33216
rect 42946 33151 43262 33152
rect 10685 33148 10751 33149
rect 10685 33144 10732 33148
rect 10796 33146 10802 33148
rect 10685 33088 10690 33144
rect 10685 33084 10732 33088
rect 10796 33086 10842 33146
rect 10796 33084 10802 33086
rect 10685 33083 10751 33084
rect 7946 32672 8262 32673
rect 0 32602 800 32632
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 27946 32672 28262 32673
rect 27946 32608 27952 32672
rect 28016 32608 28032 32672
rect 28096 32608 28112 32672
rect 28176 32608 28192 32672
rect 28256 32608 28262 32672
rect 27946 32607 28262 32608
rect 37946 32672 38262 32673
rect 37946 32608 37952 32672
rect 38016 32608 38032 32672
rect 38096 32608 38112 32672
rect 38176 32608 38192 32672
rect 38256 32608 38262 32672
rect 37946 32607 38262 32608
rect 47946 32672 48262 32673
rect 47946 32608 47952 32672
rect 48016 32608 48032 32672
rect 48096 32608 48112 32672
rect 48176 32608 48192 32672
rect 48256 32608 48262 32672
rect 47946 32607 48262 32608
rect 1301 32602 1367 32605
rect 0 32600 1367 32602
rect 0 32544 1306 32600
rect 1362 32544 1367 32600
rect 0 32542 1367 32544
rect 0 32512 800 32542
rect 1301 32539 1367 32542
rect 9213 32602 9279 32605
rect 15469 32602 15535 32605
rect 9213 32600 15535 32602
rect 9213 32544 9218 32600
rect 9274 32544 15474 32600
rect 15530 32544 15535 32600
rect 9213 32542 15535 32544
rect 9213 32539 9279 32542
rect 15469 32539 15535 32542
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 32946 32128 33262 32129
rect 32946 32064 32952 32128
rect 33016 32064 33032 32128
rect 33096 32064 33112 32128
rect 33176 32064 33192 32128
rect 33256 32064 33262 32128
rect 32946 32063 33262 32064
rect 42946 32128 43262 32129
rect 42946 32064 42952 32128
rect 43016 32064 43032 32128
rect 43096 32064 43112 32128
rect 43176 32064 43192 32128
rect 43256 32064 43262 32128
rect 42946 32063 43262 32064
rect 0 31786 800 31816
rect 1301 31786 1367 31789
rect 0 31784 1367 31786
rect 0 31728 1306 31784
rect 1362 31728 1367 31784
rect 0 31726 1367 31728
rect 0 31696 800 31726
rect 1301 31723 1367 31726
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 27946 31584 28262 31585
rect 27946 31520 27952 31584
rect 28016 31520 28032 31584
rect 28096 31520 28112 31584
rect 28176 31520 28192 31584
rect 28256 31520 28262 31584
rect 27946 31519 28262 31520
rect 37946 31584 38262 31585
rect 37946 31520 37952 31584
rect 38016 31520 38032 31584
rect 38096 31520 38112 31584
rect 38176 31520 38192 31584
rect 38256 31520 38262 31584
rect 37946 31519 38262 31520
rect 47946 31584 48262 31585
rect 47946 31520 47952 31584
rect 48016 31520 48032 31584
rect 48096 31520 48112 31584
rect 48176 31520 48192 31584
rect 48256 31520 48262 31584
rect 47946 31519 48262 31520
rect 2946 31040 3262 31041
rect 0 30970 800 31000
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 32946 31040 33262 31041
rect 32946 30976 32952 31040
rect 33016 30976 33032 31040
rect 33096 30976 33112 31040
rect 33176 30976 33192 31040
rect 33256 30976 33262 31040
rect 32946 30975 33262 30976
rect 42946 31040 43262 31041
rect 42946 30976 42952 31040
rect 43016 30976 43032 31040
rect 43096 30976 43112 31040
rect 43176 30976 43192 31040
rect 43256 30976 43262 31040
rect 42946 30975 43262 30976
rect 1301 30970 1367 30973
rect 0 30968 1367 30970
rect 0 30912 1306 30968
rect 1362 30912 1367 30968
rect 0 30910 1367 30912
rect 0 30880 800 30910
rect 1301 30907 1367 30910
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 27946 30496 28262 30497
rect 27946 30432 27952 30496
rect 28016 30432 28032 30496
rect 28096 30432 28112 30496
rect 28176 30432 28192 30496
rect 28256 30432 28262 30496
rect 27946 30431 28262 30432
rect 37946 30496 38262 30497
rect 37946 30432 37952 30496
rect 38016 30432 38032 30496
rect 38096 30432 38112 30496
rect 38176 30432 38192 30496
rect 38256 30432 38262 30496
rect 37946 30431 38262 30432
rect 47946 30496 48262 30497
rect 47946 30432 47952 30496
rect 48016 30432 48032 30496
rect 48096 30432 48112 30496
rect 48176 30432 48192 30496
rect 48256 30432 48262 30496
rect 47946 30431 48262 30432
rect 0 30154 800 30184
rect 1301 30154 1367 30157
rect 0 30152 1367 30154
rect 0 30096 1306 30152
rect 1362 30096 1367 30152
rect 0 30094 1367 30096
rect 0 30064 800 30094
rect 1301 30091 1367 30094
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 32946 29952 33262 29953
rect 32946 29888 32952 29952
rect 33016 29888 33032 29952
rect 33096 29888 33112 29952
rect 33176 29888 33192 29952
rect 33256 29888 33262 29952
rect 32946 29887 33262 29888
rect 42946 29952 43262 29953
rect 42946 29888 42952 29952
rect 43016 29888 43032 29952
rect 43096 29888 43112 29952
rect 43176 29888 43192 29952
rect 43256 29888 43262 29952
rect 42946 29887 43262 29888
rect 7946 29408 8262 29409
rect 0 29338 800 29368
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 27946 29408 28262 29409
rect 27946 29344 27952 29408
rect 28016 29344 28032 29408
rect 28096 29344 28112 29408
rect 28176 29344 28192 29408
rect 28256 29344 28262 29408
rect 27946 29343 28262 29344
rect 37946 29408 38262 29409
rect 37946 29344 37952 29408
rect 38016 29344 38032 29408
rect 38096 29344 38112 29408
rect 38176 29344 38192 29408
rect 38256 29344 38262 29408
rect 37946 29343 38262 29344
rect 47946 29408 48262 29409
rect 47946 29344 47952 29408
rect 48016 29344 48032 29408
rect 48096 29344 48112 29408
rect 48176 29344 48192 29408
rect 48256 29344 48262 29408
rect 47946 29343 48262 29344
rect 1301 29338 1367 29341
rect 0 29336 1367 29338
rect 0 29280 1306 29336
rect 1362 29280 1367 29336
rect 0 29278 1367 29280
rect 0 29248 800 29278
rect 1301 29275 1367 29278
rect 13905 29202 13971 29205
rect 13494 29200 13971 29202
rect 13494 29144 13910 29200
rect 13966 29144 13971 29200
rect 13494 29142 13971 29144
rect 11237 29066 11303 29069
rect 12617 29066 12683 29069
rect 11237 29064 12683 29066
rect 11237 29008 11242 29064
rect 11298 29008 12622 29064
rect 12678 29008 12683 29064
rect 13261 29010 13327 29013
rect 11237 29006 12683 29008
rect 11237 29003 11303 29006
rect 12617 29003 12683 29006
rect 12758 29008 13327 29010
rect 12758 28952 13266 29008
rect 13322 28952 13327 29008
rect 12758 28950 13327 28952
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 10869 28794 10935 28797
rect 12758 28794 12818 28950
rect 13261 28947 13327 28950
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 10869 28792 12818 28794
rect 10869 28736 10874 28792
rect 10930 28736 12818 28792
rect 10869 28734 12818 28736
rect 13494 28794 13554 29142
rect 13905 29139 13971 29142
rect 13813 29010 13879 29013
rect 13813 29008 13922 29010
rect 13813 28952 13818 29008
rect 13874 28952 13922 29008
rect 13813 28947 13922 28952
rect 13862 28930 13922 28947
rect 13997 28930 14063 28933
rect 13862 28928 14063 28930
rect 13862 28872 14002 28928
rect 14058 28872 14063 28928
rect 13862 28870 14063 28872
rect 13997 28867 14063 28870
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 32946 28864 33262 28865
rect 32946 28800 32952 28864
rect 33016 28800 33032 28864
rect 33096 28800 33112 28864
rect 33176 28800 33192 28864
rect 33256 28800 33262 28864
rect 32946 28799 33262 28800
rect 42946 28864 43262 28865
rect 42946 28800 42952 28864
rect 43016 28800 43032 28864
rect 43096 28800 43112 28864
rect 43176 28800 43192 28864
rect 43256 28800 43262 28864
rect 42946 28799 43262 28800
rect 13813 28794 13879 28797
rect 13494 28792 13879 28794
rect 13494 28736 13818 28792
rect 13874 28736 13879 28792
rect 13494 28734 13879 28736
rect 10869 28731 10935 28734
rect 13813 28731 13879 28734
rect 1761 28658 1827 28661
rect 18822 28658 18828 28660
rect 1761 28656 18828 28658
rect 1761 28600 1766 28656
rect 1822 28600 18828 28656
rect 1761 28598 18828 28600
rect 1761 28595 1827 28598
rect 18822 28596 18828 28598
rect 18892 28596 18898 28660
rect 0 28522 800 28552
rect 1301 28522 1367 28525
rect 0 28520 1367 28522
rect 0 28464 1306 28520
rect 1362 28464 1367 28520
rect 0 28462 1367 28464
rect 0 28432 800 28462
rect 1301 28459 1367 28462
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 27946 28320 28262 28321
rect 27946 28256 27952 28320
rect 28016 28256 28032 28320
rect 28096 28256 28112 28320
rect 28176 28256 28192 28320
rect 28256 28256 28262 28320
rect 27946 28255 28262 28256
rect 37946 28320 38262 28321
rect 37946 28256 37952 28320
rect 38016 28256 38032 28320
rect 38096 28256 38112 28320
rect 38176 28256 38192 28320
rect 38256 28256 38262 28320
rect 37946 28255 38262 28256
rect 47946 28320 48262 28321
rect 47946 28256 47952 28320
rect 48016 28256 48032 28320
rect 48096 28256 48112 28320
rect 48176 28256 48192 28320
rect 48256 28256 48262 28320
rect 47946 28255 48262 28256
rect 2946 27776 3262 27777
rect 0 27706 800 27736
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 32946 27776 33262 27777
rect 32946 27712 32952 27776
rect 33016 27712 33032 27776
rect 33096 27712 33112 27776
rect 33176 27712 33192 27776
rect 33256 27712 33262 27776
rect 32946 27711 33262 27712
rect 42946 27776 43262 27777
rect 42946 27712 42952 27776
rect 43016 27712 43032 27776
rect 43096 27712 43112 27776
rect 43176 27712 43192 27776
rect 43256 27712 43262 27776
rect 42946 27711 43262 27712
rect 1301 27706 1367 27709
rect 0 27704 1367 27706
rect 0 27648 1306 27704
rect 1362 27648 1367 27704
rect 0 27646 1367 27648
rect 0 27616 800 27646
rect 1301 27643 1367 27646
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 27946 27232 28262 27233
rect 27946 27168 27952 27232
rect 28016 27168 28032 27232
rect 28096 27168 28112 27232
rect 28176 27168 28192 27232
rect 28256 27168 28262 27232
rect 27946 27167 28262 27168
rect 37946 27232 38262 27233
rect 37946 27168 37952 27232
rect 38016 27168 38032 27232
rect 38096 27168 38112 27232
rect 38176 27168 38192 27232
rect 38256 27168 38262 27232
rect 37946 27167 38262 27168
rect 47946 27232 48262 27233
rect 47946 27168 47952 27232
rect 48016 27168 48032 27232
rect 48096 27168 48112 27232
rect 48176 27168 48192 27232
rect 48256 27168 48262 27232
rect 47946 27167 48262 27168
rect 0 26890 800 26920
rect 933 26890 999 26893
rect 0 26888 999 26890
rect 0 26832 938 26888
rect 994 26832 999 26888
rect 0 26830 999 26832
rect 0 26800 800 26830
rect 933 26827 999 26830
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 32946 26688 33262 26689
rect 32946 26624 32952 26688
rect 33016 26624 33032 26688
rect 33096 26624 33112 26688
rect 33176 26624 33192 26688
rect 33256 26624 33262 26688
rect 32946 26623 33262 26624
rect 42946 26688 43262 26689
rect 42946 26624 42952 26688
rect 43016 26624 43032 26688
rect 43096 26624 43112 26688
rect 43176 26624 43192 26688
rect 43256 26624 43262 26688
rect 42946 26623 43262 26624
rect 7946 26144 8262 26145
rect 0 26074 800 26104
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 27946 26144 28262 26145
rect 27946 26080 27952 26144
rect 28016 26080 28032 26144
rect 28096 26080 28112 26144
rect 28176 26080 28192 26144
rect 28256 26080 28262 26144
rect 27946 26079 28262 26080
rect 37946 26144 38262 26145
rect 37946 26080 37952 26144
rect 38016 26080 38032 26144
rect 38096 26080 38112 26144
rect 38176 26080 38192 26144
rect 38256 26080 38262 26144
rect 37946 26079 38262 26080
rect 47946 26144 48262 26145
rect 47946 26080 47952 26144
rect 48016 26080 48032 26144
rect 48096 26080 48112 26144
rect 48176 26080 48192 26144
rect 48256 26080 48262 26144
rect 47946 26079 48262 26080
rect 1577 26074 1643 26077
rect 0 26072 1643 26074
rect 0 26016 1582 26072
rect 1638 26016 1643 26072
rect 0 26014 1643 26016
rect 0 25984 800 26014
rect 1577 26011 1643 26014
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 32946 25600 33262 25601
rect 32946 25536 32952 25600
rect 33016 25536 33032 25600
rect 33096 25536 33112 25600
rect 33176 25536 33192 25600
rect 33256 25536 33262 25600
rect 32946 25535 33262 25536
rect 42946 25600 43262 25601
rect 42946 25536 42952 25600
rect 43016 25536 43032 25600
rect 43096 25536 43112 25600
rect 43176 25536 43192 25600
rect 43256 25536 43262 25600
rect 42946 25535 43262 25536
rect 0 25258 800 25288
rect 933 25258 999 25261
rect 0 25256 999 25258
rect 0 25200 938 25256
rect 994 25200 999 25256
rect 0 25198 999 25200
rect 0 25168 800 25198
rect 933 25195 999 25198
rect 7946 25056 8262 25057
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 27946 25056 28262 25057
rect 27946 24992 27952 25056
rect 28016 24992 28032 25056
rect 28096 24992 28112 25056
rect 28176 24992 28192 25056
rect 28256 24992 28262 25056
rect 27946 24991 28262 24992
rect 37946 25056 38262 25057
rect 37946 24992 37952 25056
rect 38016 24992 38032 25056
rect 38096 24992 38112 25056
rect 38176 24992 38192 25056
rect 38256 24992 38262 25056
rect 37946 24991 38262 24992
rect 47946 25056 48262 25057
rect 47946 24992 47952 25056
rect 48016 24992 48032 25056
rect 48096 24992 48112 25056
rect 48176 24992 48192 25056
rect 48256 24992 48262 25056
rect 47946 24991 48262 24992
rect 2946 24512 3262 24513
rect 0 24442 800 24472
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 933 24442 999 24445
rect 0 24440 999 24442
rect 0 24384 938 24440
rect 994 24384 999 24440
rect 0 24382 999 24384
rect 0 24352 800 24382
rect 933 24379 999 24382
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 0 23626 800 23656
rect 933 23626 999 23629
rect 0 23624 999 23626
rect 0 23568 938 23624
rect 994 23568 999 23624
rect 0 23566 999 23568
rect 0 23536 800 23566
rect 933 23563 999 23566
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 42946 23359 43262 23360
rect 7946 22880 8262 22881
rect 0 22810 800 22840
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 47946 22815 48262 22816
rect 933 22810 999 22813
rect 0 22808 999 22810
rect 0 22752 938 22808
rect 994 22752 999 22808
rect 0 22750 999 22752
rect 0 22720 800 22750
rect 933 22747 999 22750
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 0 21994 800 22024
rect 933 21994 999 21997
rect 0 21992 999 21994
rect 0 21936 938 21992
rect 994 21936 999 21992
rect 0 21934 999 21936
rect 0 21904 800 21934
rect 933 21931 999 21934
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 47946 21727 48262 21728
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 933 21178 999 21181
rect 0 21176 999 21178
rect 0 21120 938 21176
rect 994 21120 999 21176
rect 0 21118 999 21120
rect 0 21088 800 21118
rect 933 21115 999 21118
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 0 20362 800 20392
rect 933 20362 999 20365
rect 0 20360 999 20362
rect 0 20304 938 20360
rect 994 20304 999 20360
rect 0 20302 999 20304
rect 0 20272 800 20302
rect 933 20299 999 20302
rect 1853 20362 1919 20365
rect 7230 20362 7236 20364
rect 1853 20360 7236 20362
rect 1853 20304 1858 20360
rect 1914 20304 7236 20360
rect 1853 20302 7236 20304
rect 1853 20299 1919 20302
rect 7230 20300 7236 20302
rect 7300 20300 7306 20364
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 42946 20095 43262 20096
rect 7946 19616 8262 19617
rect 0 19546 800 19576
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 933 19546 999 19549
rect 0 19544 999 19546
rect 0 19488 938 19544
rect 994 19488 999 19544
rect 0 19486 999 19488
rect 0 19456 800 19486
rect 933 19483 999 19486
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 0 18730 800 18760
rect 933 18730 999 18733
rect 0 18728 999 18730
rect 0 18672 938 18728
rect 994 18672 999 18728
rect 0 18670 999 18672
rect 0 18640 800 18670
rect 933 18667 999 18670
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 47946 18463 48262 18464
rect 2946 17984 3262 17985
rect 0 17914 800 17944
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 1761 17914 1827 17917
rect 0 17912 1827 17914
rect 0 17856 1766 17912
rect 1822 17856 1827 17912
rect 0 17854 1827 17856
rect 0 17824 800 17854
rect 1761 17851 1827 17854
rect 1945 17778 2011 17781
rect 9438 17778 9444 17780
rect 1945 17776 9444 17778
rect 1945 17720 1950 17776
rect 2006 17720 9444 17776
rect 1945 17718 9444 17720
rect 1945 17715 2011 17718
rect 9438 17716 9444 17718
rect 9508 17716 9514 17780
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 0 17098 800 17128
rect 933 17098 999 17101
rect 0 17096 999 17098
rect 0 17040 938 17096
rect 994 17040 999 17096
rect 0 17038 999 17040
rect 0 17008 800 17038
rect 933 17035 999 17038
rect 1853 17098 1919 17101
rect 10910 17098 10916 17100
rect 1853 17096 10916 17098
rect 1853 17040 1858 17096
rect 1914 17040 10916 17096
rect 1853 17038 10916 17040
rect 1853 17035 1919 17038
rect 10910 17036 10916 17038
rect 10980 17036 10986 17100
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 42946 16831 43262 16832
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 933 16282 999 16285
rect 0 16280 999 16282
rect 0 16224 938 16280
rect 994 16224 999 16280
rect 0 16222 999 16224
rect 0 16192 800 16222
rect 933 16219 999 16222
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 0 15466 800 15496
rect 933 15466 999 15469
rect 0 15464 999 15466
rect 0 15408 938 15464
rect 994 15408 999 15464
rect 0 15406 999 15408
rect 0 15376 800 15406
rect 933 15403 999 15406
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 47946 15199 48262 15200
rect 2946 14720 3262 14721
rect 0 14650 800 14680
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 933 14650 999 14653
rect 0 14648 999 14650
rect 0 14592 938 14648
rect 994 14592 999 14648
rect 0 14590 999 14592
rect 0 14560 800 14590
rect 933 14587 999 14590
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 0 13834 800 13864
rect 933 13834 999 13837
rect 0 13832 999 13834
rect 0 13776 938 13832
rect 994 13776 999 13832
rect 0 13774 999 13776
rect 0 13744 800 13774
rect 933 13771 999 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 42946 13567 43262 13568
rect 7946 13088 8262 13089
rect 0 13018 800 13048
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 933 13018 999 13021
rect 0 13016 999 13018
rect 0 12960 938 13016
rect 994 12960 999 13016
rect 0 12958 999 12960
rect 0 12928 800 12958
rect 933 12955 999 12958
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 0 12202 800 12232
rect 933 12202 999 12205
rect 0 12200 999 12202
rect 0 12144 938 12200
rect 994 12144 999 12200
rect 0 12142 999 12144
rect 0 12112 800 12142
rect 933 12139 999 12142
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 47946 11935 48262 11936
rect 2946 11456 3262 11457
rect 0 11386 800 11416
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 933 11386 999 11389
rect 0 11384 999 11386
rect 0 11328 938 11384
rect 994 11328 999 11384
rect 0 11326 999 11328
rect 0 11296 800 11326
rect 933 11323 999 11326
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 0 10570 800 10600
rect 933 10570 999 10573
rect 0 10568 999 10570
rect 0 10512 938 10568
rect 994 10512 999 10568
rect 0 10510 999 10512
rect 0 10480 800 10510
rect 933 10507 999 10510
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 42946 10303 43262 10304
rect 7946 9824 8262 9825
rect 0 9754 800 9784
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 933 9754 999 9757
rect 0 9752 999 9754
rect 0 9696 938 9752
rect 994 9696 999 9752
rect 0 9694 999 9696
rect 0 9664 800 9694
rect 933 9691 999 9694
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 47946 8671 48262 8672
rect 2946 8192 3262 8193
rect 0 8122 800 8152
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 1761 8122 1827 8125
rect 0 8120 1827 8122
rect 0 8064 1766 8120
rect 1822 8064 1827 8120
rect 0 8062 1827 8064
rect 0 8032 800 8062
rect 1761 8059 1827 8062
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 0 7306 800 7336
rect 933 7306 999 7309
rect 0 7304 999 7306
rect 0 7248 938 7304
rect 994 7248 999 7304
rect 0 7246 999 7248
rect 0 7216 800 7246
rect 933 7243 999 7246
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 42946 7039 43262 7040
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 933 6490 999 6493
rect 0 6488 999 6490
rect 0 6432 938 6488
rect 994 6432 999 6488
rect 0 6430 999 6432
rect 0 6400 800 6430
rect 933 6427 999 6430
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 0 5674 800 5704
rect 933 5674 999 5677
rect 0 5672 999 5674
rect 0 5616 938 5672
rect 994 5616 999 5672
rect 0 5614 999 5616
rect 0 5584 800 5614
rect 933 5611 999 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 47946 5407 48262 5408
rect 2946 4928 3262 4929
rect 0 4858 800 4888
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4768 800 4798
rect 933 4795 999 4798
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 0 4042 800 4072
rect 933 4042 999 4045
rect 0 4040 999 4042
rect 0 3984 938 4040
rect 994 3984 999 4040
rect 0 3982 999 3984
rect 0 3952 800 3982
rect 933 3979 999 3982
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 42946 3775 43262 3776
rect 7946 3296 8262 3297
rect 0 3226 800 3256
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 933 3226 999 3229
rect 0 3224 999 3226
rect 0 3168 938 3224
rect 994 3168 999 3224
rect 0 3166 999 3168
rect 0 3136 800 3166
rect 933 3163 999 3166
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 47946 2143 48262 2144
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 27952 54428 28016 54432
rect 27952 54372 27956 54428
rect 27956 54372 28012 54428
rect 28012 54372 28016 54428
rect 27952 54368 28016 54372
rect 28032 54428 28096 54432
rect 28032 54372 28036 54428
rect 28036 54372 28092 54428
rect 28092 54372 28096 54428
rect 28032 54368 28096 54372
rect 28112 54428 28176 54432
rect 28112 54372 28116 54428
rect 28116 54372 28172 54428
rect 28172 54372 28176 54428
rect 28112 54368 28176 54372
rect 28192 54428 28256 54432
rect 28192 54372 28196 54428
rect 28196 54372 28252 54428
rect 28252 54372 28256 54428
rect 28192 54368 28256 54372
rect 37952 54428 38016 54432
rect 37952 54372 37956 54428
rect 37956 54372 38012 54428
rect 38012 54372 38016 54428
rect 37952 54368 38016 54372
rect 38032 54428 38096 54432
rect 38032 54372 38036 54428
rect 38036 54372 38092 54428
rect 38092 54372 38096 54428
rect 38032 54368 38096 54372
rect 38112 54428 38176 54432
rect 38112 54372 38116 54428
rect 38116 54372 38172 54428
rect 38172 54372 38176 54428
rect 38112 54368 38176 54372
rect 38192 54428 38256 54432
rect 38192 54372 38196 54428
rect 38196 54372 38252 54428
rect 38252 54372 38256 54428
rect 38192 54368 38256 54372
rect 47952 54428 48016 54432
rect 47952 54372 47956 54428
rect 47956 54372 48012 54428
rect 48012 54372 48016 54428
rect 47952 54368 48016 54372
rect 48032 54428 48096 54432
rect 48032 54372 48036 54428
rect 48036 54372 48092 54428
rect 48092 54372 48096 54428
rect 48032 54368 48096 54372
rect 48112 54428 48176 54432
rect 48112 54372 48116 54428
rect 48116 54372 48172 54428
rect 48172 54372 48176 54428
rect 48112 54368 48176 54372
rect 48192 54428 48256 54432
rect 48192 54372 48196 54428
rect 48196 54372 48252 54428
rect 48252 54372 48256 54428
rect 48192 54368 48256 54372
rect 11100 54028 11164 54092
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 32952 53884 33016 53888
rect 32952 53828 32956 53884
rect 32956 53828 33012 53884
rect 33012 53828 33016 53884
rect 32952 53824 33016 53828
rect 33032 53884 33096 53888
rect 33032 53828 33036 53884
rect 33036 53828 33092 53884
rect 33092 53828 33096 53884
rect 33032 53824 33096 53828
rect 33112 53884 33176 53888
rect 33112 53828 33116 53884
rect 33116 53828 33172 53884
rect 33172 53828 33176 53884
rect 33112 53824 33176 53828
rect 33192 53884 33256 53888
rect 33192 53828 33196 53884
rect 33196 53828 33252 53884
rect 33252 53828 33256 53884
rect 33192 53824 33256 53828
rect 42952 53884 43016 53888
rect 42952 53828 42956 53884
rect 42956 53828 43012 53884
rect 43012 53828 43016 53884
rect 42952 53824 43016 53828
rect 43032 53884 43096 53888
rect 43032 53828 43036 53884
rect 43036 53828 43092 53884
rect 43092 53828 43096 53884
rect 43032 53824 43096 53828
rect 43112 53884 43176 53888
rect 43112 53828 43116 53884
rect 43116 53828 43172 53884
rect 43172 53828 43176 53884
rect 43112 53824 43176 53828
rect 43192 53884 43256 53888
rect 43192 53828 43196 53884
rect 43196 53828 43252 53884
rect 43252 53828 43256 53884
rect 43192 53824 43256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 27952 53340 28016 53344
rect 27952 53284 27956 53340
rect 27956 53284 28012 53340
rect 28012 53284 28016 53340
rect 27952 53280 28016 53284
rect 28032 53340 28096 53344
rect 28032 53284 28036 53340
rect 28036 53284 28092 53340
rect 28092 53284 28096 53340
rect 28032 53280 28096 53284
rect 28112 53340 28176 53344
rect 28112 53284 28116 53340
rect 28116 53284 28172 53340
rect 28172 53284 28176 53340
rect 28112 53280 28176 53284
rect 28192 53340 28256 53344
rect 28192 53284 28196 53340
rect 28196 53284 28252 53340
rect 28252 53284 28256 53340
rect 28192 53280 28256 53284
rect 37952 53340 38016 53344
rect 37952 53284 37956 53340
rect 37956 53284 38012 53340
rect 38012 53284 38016 53340
rect 37952 53280 38016 53284
rect 38032 53340 38096 53344
rect 38032 53284 38036 53340
rect 38036 53284 38092 53340
rect 38092 53284 38096 53340
rect 38032 53280 38096 53284
rect 38112 53340 38176 53344
rect 38112 53284 38116 53340
rect 38116 53284 38172 53340
rect 38172 53284 38176 53340
rect 38112 53280 38176 53284
rect 38192 53340 38256 53344
rect 38192 53284 38196 53340
rect 38196 53284 38252 53340
rect 38252 53284 38256 53340
rect 38192 53280 38256 53284
rect 47952 53340 48016 53344
rect 47952 53284 47956 53340
rect 47956 53284 48012 53340
rect 48012 53284 48016 53340
rect 47952 53280 48016 53284
rect 48032 53340 48096 53344
rect 48032 53284 48036 53340
rect 48036 53284 48092 53340
rect 48092 53284 48096 53340
rect 48032 53280 48096 53284
rect 48112 53340 48176 53344
rect 48112 53284 48116 53340
rect 48116 53284 48172 53340
rect 48172 53284 48176 53340
rect 48112 53280 48176 53284
rect 48192 53340 48256 53344
rect 48192 53284 48196 53340
rect 48196 53284 48252 53340
rect 48252 53284 48256 53340
rect 48192 53280 48256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 32952 52796 33016 52800
rect 32952 52740 32956 52796
rect 32956 52740 33012 52796
rect 33012 52740 33016 52796
rect 32952 52736 33016 52740
rect 33032 52796 33096 52800
rect 33032 52740 33036 52796
rect 33036 52740 33092 52796
rect 33092 52740 33096 52796
rect 33032 52736 33096 52740
rect 33112 52796 33176 52800
rect 33112 52740 33116 52796
rect 33116 52740 33172 52796
rect 33172 52740 33176 52796
rect 33112 52736 33176 52740
rect 33192 52796 33256 52800
rect 33192 52740 33196 52796
rect 33196 52740 33252 52796
rect 33252 52740 33256 52796
rect 33192 52736 33256 52740
rect 42952 52796 43016 52800
rect 42952 52740 42956 52796
rect 42956 52740 43012 52796
rect 43012 52740 43016 52796
rect 42952 52736 43016 52740
rect 43032 52796 43096 52800
rect 43032 52740 43036 52796
rect 43036 52740 43092 52796
rect 43092 52740 43096 52796
rect 43032 52736 43096 52740
rect 43112 52796 43176 52800
rect 43112 52740 43116 52796
rect 43116 52740 43172 52796
rect 43172 52740 43176 52796
rect 43112 52736 43176 52740
rect 43192 52796 43256 52800
rect 43192 52740 43196 52796
rect 43196 52740 43252 52796
rect 43252 52740 43256 52796
rect 43192 52736 43256 52740
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 27952 52252 28016 52256
rect 27952 52196 27956 52252
rect 27956 52196 28012 52252
rect 28012 52196 28016 52252
rect 27952 52192 28016 52196
rect 28032 52252 28096 52256
rect 28032 52196 28036 52252
rect 28036 52196 28092 52252
rect 28092 52196 28096 52252
rect 28032 52192 28096 52196
rect 28112 52252 28176 52256
rect 28112 52196 28116 52252
rect 28116 52196 28172 52252
rect 28172 52196 28176 52252
rect 28112 52192 28176 52196
rect 28192 52252 28256 52256
rect 28192 52196 28196 52252
rect 28196 52196 28252 52252
rect 28252 52196 28256 52252
rect 28192 52192 28256 52196
rect 37952 52252 38016 52256
rect 37952 52196 37956 52252
rect 37956 52196 38012 52252
rect 38012 52196 38016 52252
rect 37952 52192 38016 52196
rect 38032 52252 38096 52256
rect 38032 52196 38036 52252
rect 38036 52196 38092 52252
rect 38092 52196 38096 52252
rect 38032 52192 38096 52196
rect 38112 52252 38176 52256
rect 38112 52196 38116 52252
rect 38116 52196 38172 52252
rect 38172 52196 38176 52252
rect 38112 52192 38176 52196
rect 38192 52252 38256 52256
rect 38192 52196 38196 52252
rect 38196 52196 38252 52252
rect 38252 52196 38256 52252
rect 38192 52192 38256 52196
rect 47952 52252 48016 52256
rect 47952 52196 47956 52252
rect 47956 52196 48012 52252
rect 48012 52196 48016 52252
rect 47952 52192 48016 52196
rect 48032 52252 48096 52256
rect 48032 52196 48036 52252
rect 48036 52196 48092 52252
rect 48092 52196 48096 52252
rect 48032 52192 48096 52196
rect 48112 52252 48176 52256
rect 48112 52196 48116 52252
rect 48116 52196 48172 52252
rect 48172 52196 48176 52252
rect 48112 52192 48176 52196
rect 48192 52252 48256 52256
rect 48192 52196 48196 52252
rect 48196 52196 48252 52252
rect 48252 52196 48256 52252
rect 48192 52192 48256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 32952 51708 33016 51712
rect 32952 51652 32956 51708
rect 32956 51652 33012 51708
rect 33012 51652 33016 51708
rect 32952 51648 33016 51652
rect 33032 51708 33096 51712
rect 33032 51652 33036 51708
rect 33036 51652 33092 51708
rect 33092 51652 33096 51708
rect 33032 51648 33096 51652
rect 33112 51708 33176 51712
rect 33112 51652 33116 51708
rect 33116 51652 33172 51708
rect 33172 51652 33176 51708
rect 33112 51648 33176 51652
rect 33192 51708 33256 51712
rect 33192 51652 33196 51708
rect 33196 51652 33252 51708
rect 33252 51652 33256 51708
rect 33192 51648 33256 51652
rect 42952 51708 43016 51712
rect 42952 51652 42956 51708
rect 42956 51652 43012 51708
rect 43012 51652 43016 51708
rect 42952 51648 43016 51652
rect 43032 51708 43096 51712
rect 43032 51652 43036 51708
rect 43036 51652 43092 51708
rect 43092 51652 43096 51708
rect 43032 51648 43096 51652
rect 43112 51708 43176 51712
rect 43112 51652 43116 51708
rect 43116 51652 43172 51708
rect 43172 51652 43176 51708
rect 43112 51648 43176 51652
rect 43192 51708 43256 51712
rect 43192 51652 43196 51708
rect 43196 51652 43252 51708
rect 43252 51652 43256 51708
rect 43192 51648 43256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 27952 51164 28016 51168
rect 27952 51108 27956 51164
rect 27956 51108 28012 51164
rect 28012 51108 28016 51164
rect 27952 51104 28016 51108
rect 28032 51164 28096 51168
rect 28032 51108 28036 51164
rect 28036 51108 28092 51164
rect 28092 51108 28096 51164
rect 28032 51104 28096 51108
rect 28112 51164 28176 51168
rect 28112 51108 28116 51164
rect 28116 51108 28172 51164
rect 28172 51108 28176 51164
rect 28112 51104 28176 51108
rect 28192 51164 28256 51168
rect 28192 51108 28196 51164
rect 28196 51108 28252 51164
rect 28252 51108 28256 51164
rect 28192 51104 28256 51108
rect 37952 51164 38016 51168
rect 37952 51108 37956 51164
rect 37956 51108 38012 51164
rect 38012 51108 38016 51164
rect 37952 51104 38016 51108
rect 38032 51164 38096 51168
rect 38032 51108 38036 51164
rect 38036 51108 38092 51164
rect 38092 51108 38096 51164
rect 38032 51104 38096 51108
rect 38112 51164 38176 51168
rect 38112 51108 38116 51164
rect 38116 51108 38172 51164
rect 38172 51108 38176 51164
rect 38112 51104 38176 51108
rect 38192 51164 38256 51168
rect 38192 51108 38196 51164
rect 38196 51108 38252 51164
rect 38252 51108 38256 51164
rect 38192 51104 38256 51108
rect 47952 51164 48016 51168
rect 47952 51108 47956 51164
rect 47956 51108 48012 51164
rect 48012 51108 48016 51164
rect 47952 51104 48016 51108
rect 48032 51164 48096 51168
rect 48032 51108 48036 51164
rect 48036 51108 48092 51164
rect 48092 51108 48096 51164
rect 48032 51104 48096 51108
rect 48112 51164 48176 51168
rect 48112 51108 48116 51164
rect 48116 51108 48172 51164
rect 48172 51108 48176 51164
rect 48112 51104 48176 51108
rect 48192 51164 48256 51168
rect 48192 51108 48196 51164
rect 48196 51108 48252 51164
rect 48252 51108 48256 51164
rect 48192 51104 48256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 32952 50620 33016 50624
rect 32952 50564 32956 50620
rect 32956 50564 33012 50620
rect 33012 50564 33016 50620
rect 32952 50560 33016 50564
rect 33032 50620 33096 50624
rect 33032 50564 33036 50620
rect 33036 50564 33092 50620
rect 33092 50564 33096 50620
rect 33032 50560 33096 50564
rect 33112 50620 33176 50624
rect 33112 50564 33116 50620
rect 33116 50564 33172 50620
rect 33172 50564 33176 50620
rect 33112 50560 33176 50564
rect 33192 50620 33256 50624
rect 33192 50564 33196 50620
rect 33196 50564 33252 50620
rect 33252 50564 33256 50620
rect 33192 50560 33256 50564
rect 42952 50620 43016 50624
rect 42952 50564 42956 50620
rect 42956 50564 43012 50620
rect 43012 50564 43016 50620
rect 42952 50560 43016 50564
rect 43032 50620 43096 50624
rect 43032 50564 43036 50620
rect 43036 50564 43092 50620
rect 43092 50564 43096 50620
rect 43032 50560 43096 50564
rect 43112 50620 43176 50624
rect 43112 50564 43116 50620
rect 43116 50564 43172 50620
rect 43172 50564 43176 50620
rect 43112 50560 43176 50564
rect 43192 50620 43256 50624
rect 43192 50564 43196 50620
rect 43196 50564 43252 50620
rect 43252 50564 43256 50620
rect 43192 50560 43256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 27952 50076 28016 50080
rect 27952 50020 27956 50076
rect 27956 50020 28012 50076
rect 28012 50020 28016 50076
rect 27952 50016 28016 50020
rect 28032 50076 28096 50080
rect 28032 50020 28036 50076
rect 28036 50020 28092 50076
rect 28092 50020 28096 50076
rect 28032 50016 28096 50020
rect 28112 50076 28176 50080
rect 28112 50020 28116 50076
rect 28116 50020 28172 50076
rect 28172 50020 28176 50076
rect 28112 50016 28176 50020
rect 28192 50076 28256 50080
rect 28192 50020 28196 50076
rect 28196 50020 28252 50076
rect 28252 50020 28256 50076
rect 28192 50016 28256 50020
rect 37952 50076 38016 50080
rect 37952 50020 37956 50076
rect 37956 50020 38012 50076
rect 38012 50020 38016 50076
rect 37952 50016 38016 50020
rect 38032 50076 38096 50080
rect 38032 50020 38036 50076
rect 38036 50020 38092 50076
rect 38092 50020 38096 50076
rect 38032 50016 38096 50020
rect 38112 50076 38176 50080
rect 38112 50020 38116 50076
rect 38116 50020 38172 50076
rect 38172 50020 38176 50076
rect 38112 50016 38176 50020
rect 38192 50076 38256 50080
rect 38192 50020 38196 50076
rect 38196 50020 38252 50076
rect 38252 50020 38256 50076
rect 38192 50016 38256 50020
rect 47952 50076 48016 50080
rect 47952 50020 47956 50076
rect 47956 50020 48012 50076
rect 48012 50020 48016 50076
rect 47952 50016 48016 50020
rect 48032 50076 48096 50080
rect 48032 50020 48036 50076
rect 48036 50020 48092 50076
rect 48092 50020 48096 50076
rect 48032 50016 48096 50020
rect 48112 50076 48176 50080
rect 48112 50020 48116 50076
rect 48116 50020 48172 50076
rect 48172 50020 48176 50076
rect 48112 50016 48176 50020
rect 48192 50076 48256 50080
rect 48192 50020 48196 50076
rect 48196 50020 48252 50076
rect 48252 50020 48256 50076
rect 48192 50016 48256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 32952 49532 33016 49536
rect 32952 49476 32956 49532
rect 32956 49476 33012 49532
rect 33012 49476 33016 49532
rect 32952 49472 33016 49476
rect 33032 49532 33096 49536
rect 33032 49476 33036 49532
rect 33036 49476 33092 49532
rect 33092 49476 33096 49532
rect 33032 49472 33096 49476
rect 33112 49532 33176 49536
rect 33112 49476 33116 49532
rect 33116 49476 33172 49532
rect 33172 49476 33176 49532
rect 33112 49472 33176 49476
rect 33192 49532 33256 49536
rect 33192 49476 33196 49532
rect 33196 49476 33252 49532
rect 33252 49476 33256 49532
rect 33192 49472 33256 49476
rect 42952 49532 43016 49536
rect 42952 49476 42956 49532
rect 42956 49476 43012 49532
rect 43012 49476 43016 49532
rect 42952 49472 43016 49476
rect 43032 49532 43096 49536
rect 43032 49476 43036 49532
rect 43036 49476 43092 49532
rect 43092 49476 43096 49532
rect 43032 49472 43096 49476
rect 43112 49532 43176 49536
rect 43112 49476 43116 49532
rect 43116 49476 43172 49532
rect 43172 49476 43176 49532
rect 43112 49472 43176 49476
rect 43192 49532 43256 49536
rect 43192 49476 43196 49532
rect 43196 49476 43252 49532
rect 43252 49476 43256 49532
rect 43192 49472 43256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 27952 48988 28016 48992
rect 27952 48932 27956 48988
rect 27956 48932 28012 48988
rect 28012 48932 28016 48988
rect 27952 48928 28016 48932
rect 28032 48988 28096 48992
rect 28032 48932 28036 48988
rect 28036 48932 28092 48988
rect 28092 48932 28096 48988
rect 28032 48928 28096 48932
rect 28112 48988 28176 48992
rect 28112 48932 28116 48988
rect 28116 48932 28172 48988
rect 28172 48932 28176 48988
rect 28112 48928 28176 48932
rect 28192 48988 28256 48992
rect 28192 48932 28196 48988
rect 28196 48932 28252 48988
rect 28252 48932 28256 48988
rect 28192 48928 28256 48932
rect 37952 48988 38016 48992
rect 37952 48932 37956 48988
rect 37956 48932 38012 48988
rect 38012 48932 38016 48988
rect 37952 48928 38016 48932
rect 38032 48988 38096 48992
rect 38032 48932 38036 48988
rect 38036 48932 38092 48988
rect 38092 48932 38096 48988
rect 38032 48928 38096 48932
rect 38112 48988 38176 48992
rect 38112 48932 38116 48988
rect 38116 48932 38172 48988
rect 38172 48932 38176 48988
rect 38112 48928 38176 48932
rect 38192 48988 38256 48992
rect 38192 48932 38196 48988
rect 38196 48932 38252 48988
rect 38252 48932 38256 48988
rect 38192 48928 38256 48932
rect 47952 48988 48016 48992
rect 47952 48932 47956 48988
rect 47956 48932 48012 48988
rect 48012 48932 48016 48988
rect 47952 48928 48016 48932
rect 48032 48988 48096 48992
rect 48032 48932 48036 48988
rect 48036 48932 48092 48988
rect 48092 48932 48096 48988
rect 48032 48928 48096 48932
rect 48112 48988 48176 48992
rect 48112 48932 48116 48988
rect 48116 48932 48172 48988
rect 48172 48932 48176 48988
rect 48112 48928 48176 48932
rect 48192 48988 48256 48992
rect 48192 48932 48196 48988
rect 48196 48932 48252 48988
rect 48252 48932 48256 48988
rect 48192 48928 48256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 32952 48444 33016 48448
rect 32952 48388 32956 48444
rect 32956 48388 33012 48444
rect 33012 48388 33016 48444
rect 32952 48384 33016 48388
rect 33032 48444 33096 48448
rect 33032 48388 33036 48444
rect 33036 48388 33092 48444
rect 33092 48388 33096 48444
rect 33032 48384 33096 48388
rect 33112 48444 33176 48448
rect 33112 48388 33116 48444
rect 33116 48388 33172 48444
rect 33172 48388 33176 48444
rect 33112 48384 33176 48388
rect 33192 48444 33256 48448
rect 33192 48388 33196 48444
rect 33196 48388 33252 48444
rect 33252 48388 33256 48444
rect 33192 48384 33256 48388
rect 42952 48444 43016 48448
rect 42952 48388 42956 48444
rect 42956 48388 43012 48444
rect 43012 48388 43016 48444
rect 42952 48384 43016 48388
rect 43032 48444 43096 48448
rect 43032 48388 43036 48444
rect 43036 48388 43092 48444
rect 43092 48388 43096 48444
rect 43032 48384 43096 48388
rect 43112 48444 43176 48448
rect 43112 48388 43116 48444
rect 43116 48388 43172 48444
rect 43172 48388 43176 48444
rect 43112 48384 43176 48388
rect 43192 48444 43256 48448
rect 43192 48388 43196 48444
rect 43196 48388 43252 48444
rect 43252 48388 43256 48444
rect 43192 48384 43256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 27952 47900 28016 47904
rect 27952 47844 27956 47900
rect 27956 47844 28012 47900
rect 28012 47844 28016 47900
rect 27952 47840 28016 47844
rect 28032 47900 28096 47904
rect 28032 47844 28036 47900
rect 28036 47844 28092 47900
rect 28092 47844 28096 47900
rect 28032 47840 28096 47844
rect 28112 47900 28176 47904
rect 28112 47844 28116 47900
rect 28116 47844 28172 47900
rect 28172 47844 28176 47900
rect 28112 47840 28176 47844
rect 28192 47900 28256 47904
rect 28192 47844 28196 47900
rect 28196 47844 28252 47900
rect 28252 47844 28256 47900
rect 28192 47840 28256 47844
rect 37952 47900 38016 47904
rect 37952 47844 37956 47900
rect 37956 47844 38012 47900
rect 38012 47844 38016 47900
rect 37952 47840 38016 47844
rect 38032 47900 38096 47904
rect 38032 47844 38036 47900
rect 38036 47844 38092 47900
rect 38092 47844 38096 47900
rect 38032 47840 38096 47844
rect 38112 47900 38176 47904
rect 38112 47844 38116 47900
rect 38116 47844 38172 47900
rect 38172 47844 38176 47900
rect 38112 47840 38176 47844
rect 38192 47900 38256 47904
rect 38192 47844 38196 47900
rect 38196 47844 38252 47900
rect 38252 47844 38256 47900
rect 38192 47840 38256 47844
rect 47952 47900 48016 47904
rect 47952 47844 47956 47900
rect 47956 47844 48012 47900
rect 48012 47844 48016 47900
rect 47952 47840 48016 47844
rect 48032 47900 48096 47904
rect 48032 47844 48036 47900
rect 48036 47844 48092 47900
rect 48092 47844 48096 47900
rect 48032 47840 48096 47844
rect 48112 47900 48176 47904
rect 48112 47844 48116 47900
rect 48116 47844 48172 47900
rect 48172 47844 48176 47900
rect 48112 47840 48176 47844
rect 48192 47900 48256 47904
rect 48192 47844 48196 47900
rect 48196 47844 48252 47900
rect 48252 47844 48256 47900
rect 48192 47840 48256 47844
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 32952 47356 33016 47360
rect 32952 47300 32956 47356
rect 32956 47300 33012 47356
rect 33012 47300 33016 47356
rect 32952 47296 33016 47300
rect 33032 47356 33096 47360
rect 33032 47300 33036 47356
rect 33036 47300 33092 47356
rect 33092 47300 33096 47356
rect 33032 47296 33096 47300
rect 33112 47356 33176 47360
rect 33112 47300 33116 47356
rect 33116 47300 33172 47356
rect 33172 47300 33176 47356
rect 33112 47296 33176 47300
rect 33192 47356 33256 47360
rect 33192 47300 33196 47356
rect 33196 47300 33252 47356
rect 33252 47300 33256 47356
rect 33192 47296 33256 47300
rect 42952 47356 43016 47360
rect 42952 47300 42956 47356
rect 42956 47300 43012 47356
rect 43012 47300 43016 47356
rect 42952 47296 43016 47300
rect 43032 47356 43096 47360
rect 43032 47300 43036 47356
rect 43036 47300 43092 47356
rect 43092 47300 43096 47356
rect 43032 47296 43096 47300
rect 43112 47356 43176 47360
rect 43112 47300 43116 47356
rect 43116 47300 43172 47356
rect 43172 47300 43176 47356
rect 43112 47296 43176 47300
rect 43192 47356 43256 47360
rect 43192 47300 43196 47356
rect 43196 47300 43252 47356
rect 43252 47300 43256 47356
rect 43192 47296 43256 47300
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 27952 46812 28016 46816
rect 27952 46756 27956 46812
rect 27956 46756 28012 46812
rect 28012 46756 28016 46812
rect 27952 46752 28016 46756
rect 28032 46812 28096 46816
rect 28032 46756 28036 46812
rect 28036 46756 28092 46812
rect 28092 46756 28096 46812
rect 28032 46752 28096 46756
rect 28112 46812 28176 46816
rect 28112 46756 28116 46812
rect 28116 46756 28172 46812
rect 28172 46756 28176 46812
rect 28112 46752 28176 46756
rect 28192 46812 28256 46816
rect 28192 46756 28196 46812
rect 28196 46756 28252 46812
rect 28252 46756 28256 46812
rect 28192 46752 28256 46756
rect 37952 46812 38016 46816
rect 37952 46756 37956 46812
rect 37956 46756 38012 46812
rect 38012 46756 38016 46812
rect 37952 46752 38016 46756
rect 38032 46812 38096 46816
rect 38032 46756 38036 46812
rect 38036 46756 38092 46812
rect 38092 46756 38096 46812
rect 38032 46752 38096 46756
rect 38112 46812 38176 46816
rect 38112 46756 38116 46812
rect 38116 46756 38172 46812
rect 38172 46756 38176 46812
rect 38112 46752 38176 46756
rect 38192 46812 38256 46816
rect 38192 46756 38196 46812
rect 38196 46756 38252 46812
rect 38252 46756 38256 46812
rect 38192 46752 38256 46756
rect 47952 46812 48016 46816
rect 47952 46756 47956 46812
rect 47956 46756 48012 46812
rect 48012 46756 48016 46812
rect 47952 46752 48016 46756
rect 48032 46812 48096 46816
rect 48032 46756 48036 46812
rect 48036 46756 48092 46812
rect 48092 46756 48096 46812
rect 48032 46752 48096 46756
rect 48112 46812 48176 46816
rect 48112 46756 48116 46812
rect 48116 46756 48172 46812
rect 48172 46756 48176 46812
rect 48112 46752 48176 46756
rect 48192 46812 48256 46816
rect 48192 46756 48196 46812
rect 48196 46756 48252 46812
rect 48252 46756 48256 46812
rect 48192 46752 48256 46756
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 32952 46268 33016 46272
rect 32952 46212 32956 46268
rect 32956 46212 33012 46268
rect 33012 46212 33016 46268
rect 32952 46208 33016 46212
rect 33032 46268 33096 46272
rect 33032 46212 33036 46268
rect 33036 46212 33092 46268
rect 33092 46212 33096 46268
rect 33032 46208 33096 46212
rect 33112 46268 33176 46272
rect 33112 46212 33116 46268
rect 33116 46212 33172 46268
rect 33172 46212 33176 46268
rect 33112 46208 33176 46212
rect 33192 46268 33256 46272
rect 33192 46212 33196 46268
rect 33196 46212 33252 46268
rect 33252 46212 33256 46268
rect 33192 46208 33256 46212
rect 42952 46268 43016 46272
rect 42952 46212 42956 46268
rect 42956 46212 43012 46268
rect 43012 46212 43016 46268
rect 42952 46208 43016 46212
rect 43032 46268 43096 46272
rect 43032 46212 43036 46268
rect 43036 46212 43092 46268
rect 43092 46212 43096 46268
rect 43032 46208 43096 46212
rect 43112 46268 43176 46272
rect 43112 46212 43116 46268
rect 43116 46212 43172 46268
rect 43172 46212 43176 46268
rect 43112 46208 43176 46212
rect 43192 46268 43256 46272
rect 43192 46212 43196 46268
rect 43196 46212 43252 46268
rect 43252 46212 43256 46268
rect 43192 46208 43256 46212
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 27952 45724 28016 45728
rect 27952 45668 27956 45724
rect 27956 45668 28012 45724
rect 28012 45668 28016 45724
rect 27952 45664 28016 45668
rect 28032 45724 28096 45728
rect 28032 45668 28036 45724
rect 28036 45668 28092 45724
rect 28092 45668 28096 45724
rect 28032 45664 28096 45668
rect 28112 45724 28176 45728
rect 28112 45668 28116 45724
rect 28116 45668 28172 45724
rect 28172 45668 28176 45724
rect 28112 45664 28176 45668
rect 28192 45724 28256 45728
rect 28192 45668 28196 45724
rect 28196 45668 28252 45724
rect 28252 45668 28256 45724
rect 28192 45664 28256 45668
rect 37952 45724 38016 45728
rect 37952 45668 37956 45724
rect 37956 45668 38012 45724
rect 38012 45668 38016 45724
rect 37952 45664 38016 45668
rect 38032 45724 38096 45728
rect 38032 45668 38036 45724
rect 38036 45668 38092 45724
rect 38092 45668 38096 45724
rect 38032 45664 38096 45668
rect 38112 45724 38176 45728
rect 38112 45668 38116 45724
rect 38116 45668 38172 45724
rect 38172 45668 38176 45724
rect 38112 45664 38176 45668
rect 38192 45724 38256 45728
rect 38192 45668 38196 45724
rect 38196 45668 38252 45724
rect 38252 45668 38256 45724
rect 38192 45664 38256 45668
rect 47952 45724 48016 45728
rect 47952 45668 47956 45724
rect 47956 45668 48012 45724
rect 48012 45668 48016 45724
rect 47952 45664 48016 45668
rect 48032 45724 48096 45728
rect 48032 45668 48036 45724
rect 48036 45668 48092 45724
rect 48092 45668 48096 45724
rect 48032 45664 48096 45668
rect 48112 45724 48176 45728
rect 48112 45668 48116 45724
rect 48116 45668 48172 45724
rect 48172 45668 48176 45724
rect 48112 45664 48176 45668
rect 48192 45724 48256 45728
rect 48192 45668 48196 45724
rect 48196 45668 48252 45724
rect 48252 45668 48256 45724
rect 48192 45664 48256 45668
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 32952 45180 33016 45184
rect 32952 45124 32956 45180
rect 32956 45124 33012 45180
rect 33012 45124 33016 45180
rect 32952 45120 33016 45124
rect 33032 45180 33096 45184
rect 33032 45124 33036 45180
rect 33036 45124 33092 45180
rect 33092 45124 33096 45180
rect 33032 45120 33096 45124
rect 33112 45180 33176 45184
rect 33112 45124 33116 45180
rect 33116 45124 33172 45180
rect 33172 45124 33176 45180
rect 33112 45120 33176 45124
rect 33192 45180 33256 45184
rect 33192 45124 33196 45180
rect 33196 45124 33252 45180
rect 33252 45124 33256 45180
rect 33192 45120 33256 45124
rect 42952 45180 43016 45184
rect 42952 45124 42956 45180
rect 42956 45124 43012 45180
rect 43012 45124 43016 45180
rect 42952 45120 43016 45124
rect 43032 45180 43096 45184
rect 43032 45124 43036 45180
rect 43036 45124 43092 45180
rect 43092 45124 43096 45180
rect 43032 45120 43096 45124
rect 43112 45180 43176 45184
rect 43112 45124 43116 45180
rect 43116 45124 43172 45180
rect 43172 45124 43176 45180
rect 43112 45120 43176 45124
rect 43192 45180 43256 45184
rect 43192 45124 43196 45180
rect 43196 45124 43252 45180
rect 43252 45124 43256 45180
rect 43192 45120 43256 45124
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 27952 44636 28016 44640
rect 27952 44580 27956 44636
rect 27956 44580 28012 44636
rect 28012 44580 28016 44636
rect 27952 44576 28016 44580
rect 28032 44636 28096 44640
rect 28032 44580 28036 44636
rect 28036 44580 28092 44636
rect 28092 44580 28096 44636
rect 28032 44576 28096 44580
rect 28112 44636 28176 44640
rect 28112 44580 28116 44636
rect 28116 44580 28172 44636
rect 28172 44580 28176 44636
rect 28112 44576 28176 44580
rect 28192 44636 28256 44640
rect 28192 44580 28196 44636
rect 28196 44580 28252 44636
rect 28252 44580 28256 44636
rect 28192 44576 28256 44580
rect 37952 44636 38016 44640
rect 37952 44580 37956 44636
rect 37956 44580 38012 44636
rect 38012 44580 38016 44636
rect 37952 44576 38016 44580
rect 38032 44636 38096 44640
rect 38032 44580 38036 44636
rect 38036 44580 38092 44636
rect 38092 44580 38096 44636
rect 38032 44576 38096 44580
rect 38112 44636 38176 44640
rect 38112 44580 38116 44636
rect 38116 44580 38172 44636
rect 38172 44580 38176 44636
rect 38112 44576 38176 44580
rect 38192 44636 38256 44640
rect 38192 44580 38196 44636
rect 38196 44580 38252 44636
rect 38252 44580 38256 44636
rect 38192 44576 38256 44580
rect 47952 44636 48016 44640
rect 47952 44580 47956 44636
rect 47956 44580 48012 44636
rect 48012 44580 48016 44636
rect 47952 44576 48016 44580
rect 48032 44636 48096 44640
rect 48032 44580 48036 44636
rect 48036 44580 48092 44636
rect 48092 44580 48096 44636
rect 48032 44576 48096 44580
rect 48112 44636 48176 44640
rect 48112 44580 48116 44636
rect 48116 44580 48172 44636
rect 48172 44580 48176 44636
rect 48112 44576 48176 44580
rect 48192 44636 48256 44640
rect 48192 44580 48196 44636
rect 48196 44580 48252 44636
rect 48252 44580 48256 44636
rect 48192 44576 48256 44580
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 32952 44092 33016 44096
rect 32952 44036 32956 44092
rect 32956 44036 33012 44092
rect 33012 44036 33016 44092
rect 32952 44032 33016 44036
rect 33032 44092 33096 44096
rect 33032 44036 33036 44092
rect 33036 44036 33092 44092
rect 33092 44036 33096 44092
rect 33032 44032 33096 44036
rect 33112 44092 33176 44096
rect 33112 44036 33116 44092
rect 33116 44036 33172 44092
rect 33172 44036 33176 44092
rect 33112 44032 33176 44036
rect 33192 44092 33256 44096
rect 33192 44036 33196 44092
rect 33196 44036 33252 44092
rect 33252 44036 33256 44092
rect 33192 44032 33256 44036
rect 42952 44092 43016 44096
rect 42952 44036 42956 44092
rect 42956 44036 43012 44092
rect 43012 44036 43016 44092
rect 42952 44032 43016 44036
rect 43032 44092 43096 44096
rect 43032 44036 43036 44092
rect 43036 44036 43092 44092
rect 43092 44036 43096 44092
rect 43032 44032 43096 44036
rect 43112 44092 43176 44096
rect 43112 44036 43116 44092
rect 43116 44036 43172 44092
rect 43172 44036 43176 44092
rect 43112 44032 43176 44036
rect 43192 44092 43256 44096
rect 43192 44036 43196 44092
rect 43196 44036 43252 44092
rect 43252 44036 43256 44092
rect 43192 44032 43256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 27952 43548 28016 43552
rect 27952 43492 27956 43548
rect 27956 43492 28012 43548
rect 28012 43492 28016 43548
rect 27952 43488 28016 43492
rect 28032 43548 28096 43552
rect 28032 43492 28036 43548
rect 28036 43492 28092 43548
rect 28092 43492 28096 43548
rect 28032 43488 28096 43492
rect 28112 43548 28176 43552
rect 28112 43492 28116 43548
rect 28116 43492 28172 43548
rect 28172 43492 28176 43548
rect 28112 43488 28176 43492
rect 28192 43548 28256 43552
rect 28192 43492 28196 43548
rect 28196 43492 28252 43548
rect 28252 43492 28256 43548
rect 28192 43488 28256 43492
rect 37952 43548 38016 43552
rect 37952 43492 37956 43548
rect 37956 43492 38012 43548
rect 38012 43492 38016 43548
rect 37952 43488 38016 43492
rect 38032 43548 38096 43552
rect 38032 43492 38036 43548
rect 38036 43492 38092 43548
rect 38092 43492 38096 43548
rect 38032 43488 38096 43492
rect 38112 43548 38176 43552
rect 38112 43492 38116 43548
rect 38116 43492 38172 43548
rect 38172 43492 38176 43548
rect 38112 43488 38176 43492
rect 38192 43548 38256 43552
rect 38192 43492 38196 43548
rect 38196 43492 38252 43548
rect 38252 43492 38256 43548
rect 38192 43488 38256 43492
rect 47952 43548 48016 43552
rect 47952 43492 47956 43548
rect 47956 43492 48012 43548
rect 48012 43492 48016 43548
rect 47952 43488 48016 43492
rect 48032 43548 48096 43552
rect 48032 43492 48036 43548
rect 48036 43492 48092 43548
rect 48092 43492 48096 43548
rect 48032 43488 48096 43492
rect 48112 43548 48176 43552
rect 48112 43492 48116 43548
rect 48116 43492 48172 43548
rect 48172 43492 48176 43548
rect 48112 43488 48176 43492
rect 48192 43548 48256 43552
rect 48192 43492 48196 43548
rect 48196 43492 48252 43548
rect 48252 43492 48256 43548
rect 48192 43488 48256 43492
rect 9260 43208 9324 43212
rect 9260 43152 9274 43208
rect 9274 43152 9324 43208
rect 9260 43148 9324 43152
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 32952 43004 33016 43008
rect 32952 42948 32956 43004
rect 32956 42948 33012 43004
rect 33012 42948 33016 43004
rect 32952 42944 33016 42948
rect 33032 43004 33096 43008
rect 33032 42948 33036 43004
rect 33036 42948 33092 43004
rect 33092 42948 33096 43004
rect 33032 42944 33096 42948
rect 33112 43004 33176 43008
rect 33112 42948 33116 43004
rect 33116 42948 33172 43004
rect 33172 42948 33176 43004
rect 33112 42944 33176 42948
rect 33192 43004 33256 43008
rect 33192 42948 33196 43004
rect 33196 42948 33252 43004
rect 33252 42948 33256 43004
rect 33192 42944 33256 42948
rect 42952 43004 43016 43008
rect 42952 42948 42956 43004
rect 42956 42948 43012 43004
rect 43012 42948 43016 43004
rect 42952 42944 43016 42948
rect 43032 43004 43096 43008
rect 43032 42948 43036 43004
rect 43036 42948 43092 43004
rect 43092 42948 43096 43004
rect 43032 42944 43096 42948
rect 43112 43004 43176 43008
rect 43112 42948 43116 43004
rect 43116 42948 43172 43004
rect 43172 42948 43176 43004
rect 43112 42944 43176 42948
rect 43192 43004 43256 43008
rect 43192 42948 43196 43004
rect 43196 42948 43252 43004
rect 43252 42948 43256 43004
rect 43192 42944 43256 42948
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 27952 42460 28016 42464
rect 27952 42404 27956 42460
rect 27956 42404 28012 42460
rect 28012 42404 28016 42460
rect 27952 42400 28016 42404
rect 28032 42460 28096 42464
rect 28032 42404 28036 42460
rect 28036 42404 28092 42460
rect 28092 42404 28096 42460
rect 28032 42400 28096 42404
rect 28112 42460 28176 42464
rect 28112 42404 28116 42460
rect 28116 42404 28172 42460
rect 28172 42404 28176 42460
rect 28112 42400 28176 42404
rect 28192 42460 28256 42464
rect 28192 42404 28196 42460
rect 28196 42404 28252 42460
rect 28252 42404 28256 42460
rect 28192 42400 28256 42404
rect 37952 42460 38016 42464
rect 37952 42404 37956 42460
rect 37956 42404 38012 42460
rect 38012 42404 38016 42460
rect 37952 42400 38016 42404
rect 38032 42460 38096 42464
rect 38032 42404 38036 42460
rect 38036 42404 38092 42460
rect 38092 42404 38096 42460
rect 38032 42400 38096 42404
rect 38112 42460 38176 42464
rect 38112 42404 38116 42460
rect 38116 42404 38172 42460
rect 38172 42404 38176 42460
rect 38112 42400 38176 42404
rect 38192 42460 38256 42464
rect 38192 42404 38196 42460
rect 38196 42404 38252 42460
rect 38252 42404 38256 42460
rect 38192 42400 38256 42404
rect 47952 42460 48016 42464
rect 47952 42404 47956 42460
rect 47956 42404 48012 42460
rect 48012 42404 48016 42460
rect 47952 42400 48016 42404
rect 48032 42460 48096 42464
rect 48032 42404 48036 42460
rect 48036 42404 48092 42460
rect 48092 42404 48096 42460
rect 48032 42400 48096 42404
rect 48112 42460 48176 42464
rect 48112 42404 48116 42460
rect 48116 42404 48172 42460
rect 48172 42404 48176 42460
rect 48112 42400 48176 42404
rect 48192 42460 48256 42464
rect 48192 42404 48196 42460
rect 48196 42404 48252 42460
rect 48252 42404 48256 42460
rect 48192 42400 48256 42404
rect 18828 41984 18892 41988
rect 18828 41928 18842 41984
rect 18842 41928 18892 41984
rect 18828 41924 18892 41928
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 32952 41916 33016 41920
rect 32952 41860 32956 41916
rect 32956 41860 33012 41916
rect 33012 41860 33016 41916
rect 32952 41856 33016 41860
rect 33032 41916 33096 41920
rect 33032 41860 33036 41916
rect 33036 41860 33092 41916
rect 33092 41860 33096 41916
rect 33032 41856 33096 41860
rect 33112 41916 33176 41920
rect 33112 41860 33116 41916
rect 33116 41860 33172 41916
rect 33172 41860 33176 41916
rect 33112 41856 33176 41860
rect 33192 41916 33256 41920
rect 33192 41860 33196 41916
rect 33196 41860 33252 41916
rect 33252 41860 33256 41916
rect 33192 41856 33256 41860
rect 42952 41916 43016 41920
rect 42952 41860 42956 41916
rect 42956 41860 43012 41916
rect 43012 41860 43016 41916
rect 42952 41856 43016 41860
rect 43032 41916 43096 41920
rect 43032 41860 43036 41916
rect 43036 41860 43092 41916
rect 43092 41860 43096 41916
rect 43032 41856 43096 41860
rect 43112 41916 43176 41920
rect 43112 41860 43116 41916
rect 43116 41860 43172 41916
rect 43172 41860 43176 41916
rect 43112 41856 43176 41860
rect 43192 41916 43256 41920
rect 43192 41860 43196 41916
rect 43196 41860 43252 41916
rect 43252 41860 43256 41916
rect 43192 41856 43256 41860
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 27952 41372 28016 41376
rect 27952 41316 27956 41372
rect 27956 41316 28012 41372
rect 28012 41316 28016 41372
rect 27952 41312 28016 41316
rect 28032 41372 28096 41376
rect 28032 41316 28036 41372
rect 28036 41316 28092 41372
rect 28092 41316 28096 41372
rect 28032 41312 28096 41316
rect 28112 41372 28176 41376
rect 28112 41316 28116 41372
rect 28116 41316 28172 41372
rect 28172 41316 28176 41372
rect 28112 41312 28176 41316
rect 28192 41372 28256 41376
rect 28192 41316 28196 41372
rect 28196 41316 28252 41372
rect 28252 41316 28256 41372
rect 28192 41312 28256 41316
rect 37952 41372 38016 41376
rect 37952 41316 37956 41372
rect 37956 41316 38012 41372
rect 38012 41316 38016 41372
rect 37952 41312 38016 41316
rect 38032 41372 38096 41376
rect 38032 41316 38036 41372
rect 38036 41316 38092 41372
rect 38092 41316 38096 41372
rect 38032 41312 38096 41316
rect 38112 41372 38176 41376
rect 38112 41316 38116 41372
rect 38116 41316 38172 41372
rect 38172 41316 38176 41372
rect 38112 41312 38176 41316
rect 38192 41372 38256 41376
rect 38192 41316 38196 41372
rect 38196 41316 38252 41372
rect 38252 41316 38256 41372
rect 38192 41312 38256 41316
rect 47952 41372 48016 41376
rect 47952 41316 47956 41372
rect 47956 41316 48012 41372
rect 48012 41316 48016 41372
rect 47952 41312 48016 41316
rect 48032 41372 48096 41376
rect 48032 41316 48036 41372
rect 48036 41316 48092 41372
rect 48092 41316 48096 41372
rect 48032 41312 48096 41316
rect 48112 41372 48176 41376
rect 48112 41316 48116 41372
rect 48116 41316 48172 41372
rect 48172 41316 48176 41372
rect 48112 41312 48176 41316
rect 48192 41372 48256 41376
rect 48192 41316 48196 41372
rect 48196 41316 48252 41372
rect 48252 41316 48256 41372
rect 48192 41312 48256 41316
rect 10732 40896 10796 40900
rect 10732 40840 10746 40896
rect 10746 40840 10796 40896
rect 10732 40836 10796 40840
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 32952 40828 33016 40832
rect 32952 40772 32956 40828
rect 32956 40772 33012 40828
rect 33012 40772 33016 40828
rect 32952 40768 33016 40772
rect 33032 40828 33096 40832
rect 33032 40772 33036 40828
rect 33036 40772 33092 40828
rect 33092 40772 33096 40828
rect 33032 40768 33096 40772
rect 33112 40828 33176 40832
rect 33112 40772 33116 40828
rect 33116 40772 33172 40828
rect 33172 40772 33176 40828
rect 33112 40768 33176 40772
rect 33192 40828 33256 40832
rect 33192 40772 33196 40828
rect 33196 40772 33252 40828
rect 33252 40772 33256 40828
rect 33192 40768 33256 40772
rect 42952 40828 43016 40832
rect 42952 40772 42956 40828
rect 42956 40772 43012 40828
rect 43012 40772 43016 40828
rect 42952 40768 43016 40772
rect 43032 40828 43096 40832
rect 43032 40772 43036 40828
rect 43036 40772 43092 40828
rect 43092 40772 43096 40828
rect 43032 40768 43096 40772
rect 43112 40828 43176 40832
rect 43112 40772 43116 40828
rect 43116 40772 43172 40828
rect 43172 40772 43176 40828
rect 43112 40768 43176 40772
rect 43192 40828 43256 40832
rect 43192 40772 43196 40828
rect 43196 40772 43252 40828
rect 43252 40772 43256 40828
rect 43192 40768 43256 40772
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 27952 40284 28016 40288
rect 27952 40228 27956 40284
rect 27956 40228 28012 40284
rect 28012 40228 28016 40284
rect 27952 40224 28016 40228
rect 28032 40284 28096 40288
rect 28032 40228 28036 40284
rect 28036 40228 28092 40284
rect 28092 40228 28096 40284
rect 28032 40224 28096 40228
rect 28112 40284 28176 40288
rect 28112 40228 28116 40284
rect 28116 40228 28172 40284
rect 28172 40228 28176 40284
rect 28112 40224 28176 40228
rect 28192 40284 28256 40288
rect 28192 40228 28196 40284
rect 28196 40228 28252 40284
rect 28252 40228 28256 40284
rect 28192 40224 28256 40228
rect 37952 40284 38016 40288
rect 37952 40228 37956 40284
rect 37956 40228 38012 40284
rect 38012 40228 38016 40284
rect 37952 40224 38016 40228
rect 38032 40284 38096 40288
rect 38032 40228 38036 40284
rect 38036 40228 38092 40284
rect 38092 40228 38096 40284
rect 38032 40224 38096 40228
rect 38112 40284 38176 40288
rect 38112 40228 38116 40284
rect 38116 40228 38172 40284
rect 38172 40228 38176 40284
rect 38112 40224 38176 40228
rect 38192 40284 38256 40288
rect 38192 40228 38196 40284
rect 38196 40228 38252 40284
rect 38252 40228 38256 40284
rect 38192 40224 38256 40228
rect 47952 40284 48016 40288
rect 47952 40228 47956 40284
rect 47956 40228 48012 40284
rect 48012 40228 48016 40284
rect 47952 40224 48016 40228
rect 48032 40284 48096 40288
rect 48032 40228 48036 40284
rect 48036 40228 48092 40284
rect 48092 40228 48096 40284
rect 48032 40224 48096 40228
rect 48112 40284 48176 40288
rect 48112 40228 48116 40284
rect 48116 40228 48172 40284
rect 48172 40228 48176 40284
rect 48112 40224 48176 40228
rect 48192 40284 48256 40288
rect 48192 40228 48196 40284
rect 48196 40228 48252 40284
rect 48252 40228 48256 40284
rect 48192 40224 48256 40228
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 32952 39740 33016 39744
rect 32952 39684 32956 39740
rect 32956 39684 33012 39740
rect 33012 39684 33016 39740
rect 32952 39680 33016 39684
rect 33032 39740 33096 39744
rect 33032 39684 33036 39740
rect 33036 39684 33092 39740
rect 33092 39684 33096 39740
rect 33032 39680 33096 39684
rect 33112 39740 33176 39744
rect 33112 39684 33116 39740
rect 33116 39684 33172 39740
rect 33172 39684 33176 39740
rect 33112 39680 33176 39684
rect 33192 39740 33256 39744
rect 33192 39684 33196 39740
rect 33196 39684 33252 39740
rect 33252 39684 33256 39740
rect 33192 39680 33256 39684
rect 42952 39740 43016 39744
rect 42952 39684 42956 39740
rect 42956 39684 43012 39740
rect 43012 39684 43016 39740
rect 42952 39680 43016 39684
rect 43032 39740 43096 39744
rect 43032 39684 43036 39740
rect 43036 39684 43092 39740
rect 43092 39684 43096 39740
rect 43032 39680 43096 39684
rect 43112 39740 43176 39744
rect 43112 39684 43116 39740
rect 43116 39684 43172 39740
rect 43172 39684 43176 39740
rect 43112 39680 43176 39684
rect 43192 39740 43256 39744
rect 43192 39684 43196 39740
rect 43196 39684 43252 39740
rect 43252 39684 43256 39740
rect 43192 39680 43256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 27952 39196 28016 39200
rect 27952 39140 27956 39196
rect 27956 39140 28012 39196
rect 28012 39140 28016 39196
rect 27952 39136 28016 39140
rect 28032 39196 28096 39200
rect 28032 39140 28036 39196
rect 28036 39140 28092 39196
rect 28092 39140 28096 39196
rect 28032 39136 28096 39140
rect 28112 39196 28176 39200
rect 28112 39140 28116 39196
rect 28116 39140 28172 39196
rect 28172 39140 28176 39196
rect 28112 39136 28176 39140
rect 28192 39196 28256 39200
rect 28192 39140 28196 39196
rect 28196 39140 28252 39196
rect 28252 39140 28256 39196
rect 28192 39136 28256 39140
rect 37952 39196 38016 39200
rect 37952 39140 37956 39196
rect 37956 39140 38012 39196
rect 38012 39140 38016 39196
rect 37952 39136 38016 39140
rect 38032 39196 38096 39200
rect 38032 39140 38036 39196
rect 38036 39140 38092 39196
rect 38092 39140 38096 39196
rect 38032 39136 38096 39140
rect 38112 39196 38176 39200
rect 38112 39140 38116 39196
rect 38116 39140 38172 39196
rect 38172 39140 38176 39196
rect 38112 39136 38176 39140
rect 38192 39196 38256 39200
rect 38192 39140 38196 39196
rect 38196 39140 38252 39196
rect 38252 39140 38256 39196
rect 38192 39136 38256 39140
rect 47952 39196 48016 39200
rect 47952 39140 47956 39196
rect 47956 39140 48012 39196
rect 48012 39140 48016 39196
rect 47952 39136 48016 39140
rect 48032 39196 48096 39200
rect 48032 39140 48036 39196
rect 48036 39140 48092 39196
rect 48092 39140 48096 39196
rect 48032 39136 48096 39140
rect 48112 39196 48176 39200
rect 48112 39140 48116 39196
rect 48116 39140 48172 39196
rect 48172 39140 48176 39196
rect 48112 39136 48176 39140
rect 48192 39196 48256 39200
rect 48192 39140 48196 39196
rect 48196 39140 48252 39196
rect 48252 39140 48256 39196
rect 48192 39136 48256 39140
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 32952 38652 33016 38656
rect 32952 38596 32956 38652
rect 32956 38596 33012 38652
rect 33012 38596 33016 38652
rect 32952 38592 33016 38596
rect 33032 38652 33096 38656
rect 33032 38596 33036 38652
rect 33036 38596 33092 38652
rect 33092 38596 33096 38652
rect 33032 38592 33096 38596
rect 33112 38652 33176 38656
rect 33112 38596 33116 38652
rect 33116 38596 33172 38652
rect 33172 38596 33176 38652
rect 33112 38592 33176 38596
rect 33192 38652 33256 38656
rect 33192 38596 33196 38652
rect 33196 38596 33252 38652
rect 33252 38596 33256 38652
rect 33192 38592 33256 38596
rect 42952 38652 43016 38656
rect 42952 38596 42956 38652
rect 42956 38596 43012 38652
rect 43012 38596 43016 38652
rect 42952 38592 43016 38596
rect 43032 38652 43096 38656
rect 43032 38596 43036 38652
rect 43036 38596 43092 38652
rect 43092 38596 43096 38652
rect 43032 38592 43096 38596
rect 43112 38652 43176 38656
rect 43112 38596 43116 38652
rect 43116 38596 43172 38652
rect 43172 38596 43176 38652
rect 43112 38592 43176 38596
rect 43192 38652 43256 38656
rect 43192 38596 43196 38652
rect 43196 38596 43252 38652
rect 43252 38596 43256 38652
rect 43192 38592 43256 38596
rect 10916 38176 10980 38180
rect 10916 38120 10930 38176
rect 10930 38120 10980 38176
rect 10916 38116 10980 38120
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 27952 38108 28016 38112
rect 27952 38052 27956 38108
rect 27956 38052 28012 38108
rect 28012 38052 28016 38108
rect 27952 38048 28016 38052
rect 28032 38108 28096 38112
rect 28032 38052 28036 38108
rect 28036 38052 28092 38108
rect 28092 38052 28096 38108
rect 28032 38048 28096 38052
rect 28112 38108 28176 38112
rect 28112 38052 28116 38108
rect 28116 38052 28172 38108
rect 28172 38052 28176 38108
rect 28112 38048 28176 38052
rect 28192 38108 28256 38112
rect 28192 38052 28196 38108
rect 28196 38052 28252 38108
rect 28252 38052 28256 38108
rect 28192 38048 28256 38052
rect 37952 38108 38016 38112
rect 37952 38052 37956 38108
rect 37956 38052 38012 38108
rect 38012 38052 38016 38108
rect 37952 38048 38016 38052
rect 38032 38108 38096 38112
rect 38032 38052 38036 38108
rect 38036 38052 38092 38108
rect 38092 38052 38096 38108
rect 38032 38048 38096 38052
rect 38112 38108 38176 38112
rect 38112 38052 38116 38108
rect 38116 38052 38172 38108
rect 38172 38052 38176 38108
rect 38112 38048 38176 38052
rect 38192 38108 38256 38112
rect 38192 38052 38196 38108
rect 38196 38052 38252 38108
rect 38252 38052 38256 38108
rect 38192 38048 38256 38052
rect 47952 38108 48016 38112
rect 47952 38052 47956 38108
rect 47956 38052 48012 38108
rect 48012 38052 48016 38108
rect 47952 38048 48016 38052
rect 48032 38108 48096 38112
rect 48032 38052 48036 38108
rect 48036 38052 48092 38108
rect 48092 38052 48096 38108
rect 48032 38048 48096 38052
rect 48112 38108 48176 38112
rect 48112 38052 48116 38108
rect 48116 38052 48172 38108
rect 48172 38052 48176 38108
rect 48112 38048 48176 38052
rect 48192 38108 48256 38112
rect 48192 38052 48196 38108
rect 48196 38052 48252 38108
rect 48252 38052 48256 38108
rect 48192 38048 48256 38052
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 32952 37564 33016 37568
rect 32952 37508 32956 37564
rect 32956 37508 33012 37564
rect 33012 37508 33016 37564
rect 32952 37504 33016 37508
rect 33032 37564 33096 37568
rect 33032 37508 33036 37564
rect 33036 37508 33092 37564
rect 33092 37508 33096 37564
rect 33032 37504 33096 37508
rect 33112 37564 33176 37568
rect 33112 37508 33116 37564
rect 33116 37508 33172 37564
rect 33172 37508 33176 37564
rect 33112 37504 33176 37508
rect 33192 37564 33256 37568
rect 33192 37508 33196 37564
rect 33196 37508 33252 37564
rect 33252 37508 33256 37564
rect 33192 37504 33256 37508
rect 42952 37564 43016 37568
rect 42952 37508 42956 37564
rect 42956 37508 43012 37564
rect 43012 37508 43016 37564
rect 42952 37504 43016 37508
rect 43032 37564 43096 37568
rect 43032 37508 43036 37564
rect 43036 37508 43092 37564
rect 43092 37508 43096 37564
rect 43032 37504 43096 37508
rect 43112 37564 43176 37568
rect 43112 37508 43116 37564
rect 43116 37508 43172 37564
rect 43172 37508 43176 37564
rect 43112 37504 43176 37508
rect 43192 37564 43256 37568
rect 43192 37508 43196 37564
rect 43196 37508 43252 37564
rect 43252 37508 43256 37564
rect 43192 37504 43256 37508
rect 11100 37224 11164 37228
rect 11100 37168 11114 37224
rect 11114 37168 11164 37224
rect 11100 37164 11164 37168
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 27952 37020 28016 37024
rect 27952 36964 27956 37020
rect 27956 36964 28012 37020
rect 28012 36964 28016 37020
rect 27952 36960 28016 36964
rect 28032 37020 28096 37024
rect 28032 36964 28036 37020
rect 28036 36964 28092 37020
rect 28092 36964 28096 37020
rect 28032 36960 28096 36964
rect 28112 37020 28176 37024
rect 28112 36964 28116 37020
rect 28116 36964 28172 37020
rect 28172 36964 28176 37020
rect 28112 36960 28176 36964
rect 28192 37020 28256 37024
rect 28192 36964 28196 37020
rect 28196 36964 28252 37020
rect 28252 36964 28256 37020
rect 28192 36960 28256 36964
rect 37952 37020 38016 37024
rect 37952 36964 37956 37020
rect 37956 36964 38012 37020
rect 38012 36964 38016 37020
rect 37952 36960 38016 36964
rect 38032 37020 38096 37024
rect 38032 36964 38036 37020
rect 38036 36964 38092 37020
rect 38092 36964 38096 37020
rect 38032 36960 38096 36964
rect 38112 37020 38176 37024
rect 38112 36964 38116 37020
rect 38116 36964 38172 37020
rect 38172 36964 38176 37020
rect 38112 36960 38176 36964
rect 38192 37020 38256 37024
rect 38192 36964 38196 37020
rect 38196 36964 38252 37020
rect 38252 36964 38256 37020
rect 38192 36960 38256 36964
rect 47952 37020 48016 37024
rect 47952 36964 47956 37020
rect 47956 36964 48012 37020
rect 48012 36964 48016 37020
rect 47952 36960 48016 36964
rect 48032 37020 48096 37024
rect 48032 36964 48036 37020
rect 48036 36964 48092 37020
rect 48092 36964 48096 37020
rect 48032 36960 48096 36964
rect 48112 37020 48176 37024
rect 48112 36964 48116 37020
rect 48116 36964 48172 37020
rect 48172 36964 48176 37020
rect 48112 36960 48176 36964
rect 48192 37020 48256 37024
rect 48192 36964 48196 37020
rect 48196 36964 48252 37020
rect 48252 36964 48256 37020
rect 48192 36960 48256 36964
rect 9260 36892 9324 36956
rect 7236 36620 7300 36684
rect 9444 36620 9508 36684
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 32952 36476 33016 36480
rect 32952 36420 32956 36476
rect 32956 36420 33012 36476
rect 33012 36420 33016 36476
rect 32952 36416 33016 36420
rect 33032 36476 33096 36480
rect 33032 36420 33036 36476
rect 33036 36420 33092 36476
rect 33092 36420 33096 36476
rect 33032 36416 33096 36420
rect 33112 36476 33176 36480
rect 33112 36420 33116 36476
rect 33116 36420 33172 36476
rect 33172 36420 33176 36476
rect 33112 36416 33176 36420
rect 33192 36476 33256 36480
rect 33192 36420 33196 36476
rect 33196 36420 33252 36476
rect 33252 36420 33256 36476
rect 33192 36416 33256 36420
rect 42952 36476 43016 36480
rect 42952 36420 42956 36476
rect 42956 36420 43012 36476
rect 43012 36420 43016 36476
rect 42952 36416 43016 36420
rect 43032 36476 43096 36480
rect 43032 36420 43036 36476
rect 43036 36420 43092 36476
rect 43092 36420 43096 36476
rect 43032 36416 43096 36420
rect 43112 36476 43176 36480
rect 43112 36420 43116 36476
rect 43116 36420 43172 36476
rect 43172 36420 43176 36476
rect 43112 36416 43176 36420
rect 43192 36476 43256 36480
rect 43192 36420 43196 36476
rect 43196 36420 43252 36476
rect 43252 36420 43256 36476
rect 43192 36416 43256 36420
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 27952 35932 28016 35936
rect 27952 35876 27956 35932
rect 27956 35876 28012 35932
rect 28012 35876 28016 35932
rect 27952 35872 28016 35876
rect 28032 35932 28096 35936
rect 28032 35876 28036 35932
rect 28036 35876 28092 35932
rect 28092 35876 28096 35932
rect 28032 35872 28096 35876
rect 28112 35932 28176 35936
rect 28112 35876 28116 35932
rect 28116 35876 28172 35932
rect 28172 35876 28176 35932
rect 28112 35872 28176 35876
rect 28192 35932 28256 35936
rect 28192 35876 28196 35932
rect 28196 35876 28252 35932
rect 28252 35876 28256 35932
rect 28192 35872 28256 35876
rect 37952 35932 38016 35936
rect 37952 35876 37956 35932
rect 37956 35876 38012 35932
rect 38012 35876 38016 35932
rect 37952 35872 38016 35876
rect 38032 35932 38096 35936
rect 38032 35876 38036 35932
rect 38036 35876 38092 35932
rect 38092 35876 38096 35932
rect 38032 35872 38096 35876
rect 38112 35932 38176 35936
rect 38112 35876 38116 35932
rect 38116 35876 38172 35932
rect 38172 35876 38176 35932
rect 38112 35872 38176 35876
rect 38192 35932 38256 35936
rect 38192 35876 38196 35932
rect 38196 35876 38252 35932
rect 38252 35876 38256 35932
rect 38192 35872 38256 35876
rect 47952 35932 48016 35936
rect 47952 35876 47956 35932
rect 47956 35876 48012 35932
rect 48012 35876 48016 35932
rect 47952 35872 48016 35876
rect 48032 35932 48096 35936
rect 48032 35876 48036 35932
rect 48036 35876 48092 35932
rect 48092 35876 48096 35932
rect 48032 35872 48096 35876
rect 48112 35932 48176 35936
rect 48112 35876 48116 35932
rect 48116 35876 48172 35932
rect 48172 35876 48176 35932
rect 48112 35872 48176 35876
rect 48192 35932 48256 35936
rect 48192 35876 48196 35932
rect 48196 35876 48252 35932
rect 48252 35876 48256 35932
rect 48192 35872 48256 35876
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 32952 35388 33016 35392
rect 32952 35332 32956 35388
rect 32956 35332 33012 35388
rect 33012 35332 33016 35388
rect 32952 35328 33016 35332
rect 33032 35388 33096 35392
rect 33032 35332 33036 35388
rect 33036 35332 33092 35388
rect 33092 35332 33096 35388
rect 33032 35328 33096 35332
rect 33112 35388 33176 35392
rect 33112 35332 33116 35388
rect 33116 35332 33172 35388
rect 33172 35332 33176 35388
rect 33112 35328 33176 35332
rect 33192 35388 33256 35392
rect 33192 35332 33196 35388
rect 33196 35332 33252 35388
rect 33252 35332 33256 35388
rect 33192 35328 33256 35332
rect 42952 35388 43016 35392
rect 42952 35332 42956 35388
rect 42956 35332 43012 35388
rect 43012 35332 43016 35388
rect 42952 35328 43016 35332
rect 43032 35388 43096 35392
rect 43032 35332 43036 35388
rect 43036 35332 43092 35388
rect 43092 35332 43096 35388
rect 43032 35328 43096 35332
rect 43112 35388 43176 35392
rect 43112 35332 43116 35388
rect 43116 35332 43172 35388
rect 43172 35332 43176 35388
rect 43112 35328 43176 35332
rect 43192 35388 43256 35392
rect 43192 35332 43196 35388
rect 43196 35332 43252 35388
rect 43252 35332 43256 35388
rect 43192 35328 43256 35332
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 27952 34844 28016 34848
rect 27952 34788 27956 34844
rect 27956 34788 28012 34844
rect 28012 34788 28016 34844
rect 27952 34784 28016 34788
rect 28032 34844 28096 34848
rect 28032 34788 28036 34844
rect 28036 34788 28092 34844
rect 28092 34788 28096 34844
rect 28032 34784 28096 34788
rect 28112 34844 28176 34848
rect 28112 34788 28116 34844
rect 28116 34788 28172 34844
rect 28172 34788 28176 34844
rect 28112 34784 28176 34788
rect 28192 34844 28256 34848
rect 28192 34788 28196 34844
rect 28196 34788 28252 34844
rect 28252 34788 28256 34844
rect 28192 34784 28256 34788
rect 37952 34844 38016 34848
rect 37952 34788 37956 34844
rect 37956 34788 38012 34844
rect 38012 34788 38016 34844
rect 37952 34784 38016 34788
rect 38032 34844 38096 34848
rect 38032 34788 38036 34844
rect 38036 34788 38092 34844
rect 38092 34788 38096 34844
rect 38032 34784 38096 34788
rect 38112 34844 38176 34848
rect 38112 34788 38116 34844
rect 38116 34788 38172 34844
rect 38172 34788 38176 34844
rect 38112 34784 38176 34788
rect 38192 34844 38256 34848
rect 38192 34788 38196 34844
rect 38196 34788 38252 34844
rect 38252 34788 38256 34844
rect 38192 34784 38256 34788
rect 47952 34844 48016 34848
rect 47952 34788 47956 34844
rect 47956 34788 48012 34844
rect 48012 34788 48016 34844
rect 47952 34784 48016 34788
rect 48032 34844 48096 34848
rect 48032 34788 48036 34844
rect 48036 34788 48092 34844
rect 48092 34788 48096 34844
rect 48032 34784 48096 34788
rect 48112 34844 48176 34848
rect 48112 34788 48116 34844
rect 48116 34788 48172 34844
rect 48172 34788 48176 34844
rect 48112 34784 48176 34788
rect 48192 34844 48256 34848
rect 48192 34788 48196 34844
rect 48196 34788 48252 34844
rect 48252 34788 48256 34844
rect 48192 34784 48256 34788
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 32952 34300 33016 34304
rect 32952 34244 32956 34300
rect 32956 34244 33012 34300
rect 33012 34244 33016 34300
rect 32952 34240 33016 34244
rect 33032 34300 33096 34304
rect 33032 34244 33036 34300
rect 33036 34244 33092 34300
rect 33092 34244 33096 34300
rect 33032 34240 33096 34244
rect 33112 34300 33176 34304
rect 33112 34244 33116 34300
rect 33116 34244 33172 34300
rect 33172 34244 33176 34300
rect 33112 34240 33176 34244
rect 33192 34300 33256 34304
rect 33192 34244 33196 34300
rect 33196 34244 33252 34300
rect 33252 34244 33256 34300
rect 33192 34240 33256 34244
rect 42952 34300 43016 34304
rect 42952 34244 42956 34300
rect 42956 34244 43012 34300
rect 43012 34244 43016 34300
rect 42952 34240 43016 34244
rect 43032 34300 43096 34304
rect 43032 34244 43036 34300
rect 43036 34244 43092 34300
rect 43092 34244 43096 34300
rect 43032 34240 43096 34244
rect 43112 34300 43176 34304
rect 43112 34244 43116 34300
rect 43116 34244 43172 34300
rect 43172 34244 43176 34300
rect 43112 34240 43176 34244
rect 43192 34300 43256 34304
rect 43192 34244 43196 34300
rect 43196 34244 43252 34300
rect 43252 34244 43256 34300
rect 43192 34240 43256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 27952 33756 28016 33760
rect 27952 33700 27956 33756
rect 27956 33700 28012 33756
rect 28012 33700 28016 33756
rect 27952 33696 28016 33700
rect 28032 33756 28096 33760
rect 28032 33700 28036 33756
rect 28036 33700 28092 33756
rect 28092 33700 28096 33756
rect 28032 33696 28096 33700
rect 28112 33756 28176 33760
rect 28112 33700 28116 33756
rect 28116 33700 28172 33756
rect 28172 33700 28176 33756
rect 28112 33696 28176 33700
rect 28192 33756 28256 33760
rect 28192 33700 28196 33756
rect 28196 33700 28252 33756
rect 28252 33700 28256 33756
rect 28192 33696 28256 33700
rect 37952 33756 38016 33760
rect 37952 33700 37956 33756
rect 37956 33700 38012 33756
rect 38012 33700 38016 33756
rect 37952 33696 38016 33700
rect 38032 33756 38096 33760
rect 38032 33700 38036 33756
rect 38036 33700 38092 33756
rect 38092 33700 38096 33756
rect 38032 33696 38096 33700
rect 38112 33756 38176 33760
rect 38112 33700 38116 33756
rect 38116 33700 38172 33756
rect 38172 33700 38176 33756
rect 38112 33696 38176 33700
rect 38192 33756 38256 33760
rect 38192 33700 38196 33756
rect 38196 33700 38252 33756
rect 38252 33700 38256 33756
rect 38192 33696 38256 33700
rect 47952 33756 48016 33760
rect 47952 33700 47956 33756
rect 47956 33700 48012 33756
rect 48012 33700 48016 33756
rect 47952 33696 48016 33700
rect 48032 33756 48096 33760
rect 48032 33700 48036 33756
rect 48036 33700 48092 33756
rect 48092 33700 48096 33756
rect 48032 33696 48096 33700
rect 48112 33756 48176 33760
rect 48112 33700 48116 33756
rect 48116 33700 48172 33756
rect 48172 33700 48176 33756
rect 48112 33696 48176 33700
rect 48192 33756 48256 33760
rect 48192 33700 48196 33756
rect 48196 33700 48252 33756
rect 48252 33700 48256 33756
rect 48192 33696 48256 33700
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 32952 33212 33016 33216
rect 32952 33156 32956 33212
rect 32956 33156 33012 33212
rect 33012 33156 33016 33212
rect 32952 33152 33016 33156
rect 33032 33212 33096 33216
rect 33032 33156 33036 33212
rect 33036 33156 33092 33212
rect 33092 33156 33096 33212
rect 33032 33152 33096 33156
rect 33112 33212 33176 33216
rect 33112 33156 33116 33212
rect 33116 33156 33172 33212
rect 33172 33156 33176 33212
rect 33112 33152 33176 33156
rect 33192 33212 33256 33216
rect 33192 33156 33196 33212
rect 33196 33156 33252 33212
rect 33252 33156 33256 33212
rect 33192 33152 33256 33156
rect 42952 33212 43016 33216
rect 42952 33156 42956 33212
rect 42956 33156 43012 33212
rect 43012 33156 43016 33212
rect 42952 33152 43016 33156
rect 43032 33212 43096 33216
rect 43032 33156 43036 33212
rect 43036 33156 43092 33212
rect 43092 33156 43096 33212
rect 43032 33152 43096 33156
rect 43112 33212 43176 33216
rect 43112 33156 43116 33212
rect 43116 33156 43172 33212
rect 43172 33156 43176 33212
rect 43112 33152 43176 33156
rect 43192 33212 43256 33216
rect 43192 33156 43196 33212
rect 43196 33156 43252 33212
rect 43252 33156 43256 33212
rect 43192 33152 43256 33156
rect 10732 33144 10796 33148
rect 10732 33088 10746 33144
rect 10746 33088 10796 33144
rect 10732 33084 10796 33088
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 27952 32668 28016 32672
rect 27952 32612 27956 32668
rect 27956 32612 28012 32668
rect 28012 32612 28016 32668
rect 27952 32608 28016 32612
rect 28032 32668 28096 32672
rect 28032 32612 28036 32668
rect 28036 32612 28092 32668
rect 28092 32612 28096 32668
rect 28032 32608 28096 32612
rect 28112 32668 28176 32672
rect 28112 32612 28116 32668
rect 28116 32612 28172 32668
rect 28172 32612 28176 32668
rect 28112 32608 28176 32612
rect 28192 32668 28256 32672
rect 28192 32612 28196 32668
rect 28196 32612 28252 32668
rect 28252 32612 28256 32668
rect 28192 32608 28256 32612
rect 37952 32668 38016 32672
rect 37952 32612 37956 32668
rect 37956 32612 38012 32668
rect 38012 32612 38016 32668
rect 37952 32608 38016 32612
rect 38032 32668 38096 32672
rect 38032 32612 38036 32668
rect 38036 32612 38092 32668
rect 38092 32612 38096 32668
rect 38032 32608 38096 32612
rect 38112 32668 38176 32672
rect 38112 32612 38116 32668
rect 38116 32612 38172 32668
rect 38172 32612 38176 32668
rect 38112 32608 38176 32612
rect 38192 32668 38256 32672
rect 38192 32612 38196 32668
rect 38196 32612 38252 32668
rect 38252 32612 38256 32668
rect 38192 32608 38256 32612
rect 47952 32668 48016 32672
rect 47952 32612 47956 32668
rect 47956 32612 48012 32668
rect 48012 32612 48016 32668
rect 47952 32608 48016 32612
rect 48032 32668 48096 32672
rect 48032 32612 48036 32668
rect 48036 32612 48092 32668
rect 48092 32612 48096 32668
rect 48032 32608 48096 32612
rect 48112 32668 48176 32672
rect 48112 32612 48116 32668
rect 48116 32612 48172 32668
rect 48172 32612 48176 32668
rect 48112 32608 48176 32612
rect 48192 32668 48256 32672
rect 48192 32612 48196 32668
rect 48196 32612 48252 32668
rect 48252 32612 48256 32668
rect 48192 32608 48256 32612
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 32952 32124 33016 32128
rect 32952 32068 32956 32124
rect 32956 32068 33012 32124
rect 33012 32068 33016 32124
rect 32952 32064 33016 32068
rect 33032 32124 33096 32128
rect 33032 32068 33036 32124
rect 33036 32068 33092 32124
rect 33092 32068 33096 32124
rect 33032 32064 33096 32068
rect 33112 32124 33176 32128
rect 33112 32068 33116 32124
rect 33116 32068 33172 32124
rect 33172 32068 33176 32124
rect 33112 32064 33176 32068
rect 33192 32124 33256 32128
rect 33192 32068 33196 32124
rect 33196 32068 33252 32124
rect 33252 32068 33256 32124
rect 33192 32064 33256 32068
rect 42952 32124 43016 32128
rect 42952 32068 42956 32124
rect 42956 32068 43012 32124
rect 43012 32068 43016 32124
rect 42952 32064 43016 32068
rect 43032 32124 43096 32128
rect 43032 32068 43036 32124
rect 43036 32068 43092 32124
rect 43092 32068 43096 32124
rect 43032 32064 43096 32068
rect 43112 32124 43176 32128
rect 43112 32068 43116 32124
rect 43116 32068 43172 32124
rect 43172 32068 43176 32124
rect 43112 32064 43176 32068
rect 43192 32124 43256 32128
rect 43192 32068 43196 32124
rect 43196 32068 43252 32124
rect 43252 32068 43256 32124
rect 43192 32064 43256 32068
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 27952 31580 28016 31584
rect 27952 31524 27956 31580
rect 27956 31524 28012 31580
rect 28012 31524 28016 31580
rect 27952 31520 28016 31524
rect 28032 31580 28096 31584
rect 28032 31524 28036 31580
rect 28036 31524 28092 31580
rect 28092 31524 28096 31580
rect 28032 31520 28096 31524
rect 28112 31580 28176 31584
rect 28112 31524 28116 31580
rect 28116 31524 28172 31580
rect 28172 31524 28176 31580
rect 28112 31520 28176 31524
rect 28192 31580 28256 31584
rect 28192 31524 28196 31580
rect 28196 31524 28252 31580
rect 28252 31524 28256 31580
rect 28192 31520 28256 31524
rect 37952 31580 38016 31584
rect 37952 31524 37956 31580
rect 37956 31524 38012 31580
rect 38012 31524 38016 31580
rect 37952 31520 38016 31524
rect 38032 31580 38096 31584
rect 38032 31524 38036 31580
rect 38036 31524 38092 31580
rect 38092 31524 38096 31580
rect 38032 31520 38096 31524
rect 38112 31580 38176 31584
rect 38112 31524 38116 31580
rect 38116 31524 38172 31580
rect 38172 31524 38176 31580
rect 38112 31520 38176 31524
rect 38192 31580 38256 31584
rect 38192 31524 38196 31580
rect 38196 31524 38252 31580
rect 38252 31524 38256 31580
rect 38192 31520 38256 31524
rect 47952 31580 48016 31584
rect 47952 31524 47956 31580
rect 47956 31524 48012 31580
rect 48012 31524 48016 31580
rect 47952 31520 48016 31524
rect 48032 31580 48096 31584
rect 48032 31524 48036 31580
rect 48036 31524 48092 31580
rect 48092 31524 48096 31580
rect 48032 31520 48096 31524
rect 48112 31580 48176 31584
rect 48112 31524 48116 31580
rect 48116 31524 48172 31580
rect 48172 31524 48176 31580
rect 48112 31520 48176 31524
rect 48192 31580 48256 31584
rect 48192 31524 48196 31580
rect 48196 31524 48252 31580
rect 48252 31524 48256 31580
rect 48192 31520 48256 31524
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 32952 31036 33016 31040
rect 32952 30980 32956 31036
rect 32956 30980 33012 31036
rect 33012 30980 33016 31036
rect 32952 30976 33016 30980
rect 33032 31036 33096 31040
rect 33032 30980 33036 31036
rect 33036 30980 33092 31036
rect 33092 30980 33096 31036
rect 33032 30976 33096 30980
rect 33112 31036 33176 31040
rect 33112 30980 33116 31036
rect 33116 30980 33172 31036
rect 33172 30980 33176 31036
rect 33112 30976 33176 30980
rect 33192 31036 33256 31040
rect 33192 30980 33196 31036
rect 33196 30980 33252 31036
rect 33252 30980 33256 31036
rect 33192 30976 33256 30980
rect 42952 31036 43016 31040
rect 42952 30980 42956 31036
rect 42956 30980 43012 31036
rect 43012 30980 43016 31036
rect 42952 30976 43016 30980
rect 43032 31036 43096 31040
rect 43032 30980 43036 31036
rect 43036 30980 43092 31036
rect 43092 30980 43096 31036
rect 43032 30976 43096 30980
rect 43112 31036 43176 31040
rect 43112 30980 43116 31036
rect 43116 30980 43172 31036
rect 43172 30980 43176 31036
rect 43112 30976 43176 30980
rect 43192 31036 43256 31040
rect 43192 30980 43196 31036
rect 43196 30980 43252 31036
rect 43252 30980 43256 31036
rect 43192 30976 43256 30980
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 27952 30492 28016 30496
rect 27952 30436 27956 30492
rect 27956 30436 28012 30492
rect 28012 30436 28016 30492
rect 27952 30432 28016 30436
rect 28032 30492 28096 30496
rect 28032 30436 28036 30492
rect 28036 30436 28092 30492
rect 28092 30436 28096 30492
rect 28032 30432 28096 30436
rect 28112 30492 28176 30496
rect 28112 30436 28116 30492
rect 28116 30436 28172 30492
rect 28172 30436 28176 30492
rect 28112 30432 28176 30436
rect 28192 30492 28256 30496
rect 28192 30436 28196 30492
rect 28196 30436 28252 30492
rect 28252 30436 28256 30492
rect 28192 30432 28256 30436
rect 37952 30492 38016 30496
rect 37952 30436 37956 30492
rect 37956 30436 38012 30492
rect 38012 30436 38016 30492
rect 37952 30432 38016 30436
rect 38032 30492 38096 30496
rect 38032 30436 38036 30492
rect 38036 30436 38092 30492
rect 38092 30436 38096 30492
rect 38032 30432 38096 30436
rect 38112 30492 38176 30496
rect 38112 30436 38116 30492
rect 38116 30436 38172 30492
rect 38172 30436 38176 30492
rect 38112 30432 38176 30436
rect 38192 30492 38256 30496
rect 38192 30436 38196 30492
rect 38196 30436 38252 30492
rect 38252 30436 38256 30492
rect 38192 30432 38256 30436
rect 47952 30492 48016 30496
rect 47952 30436 47956 30492
rect 47956 30436 48012 30492
rect 48012 30436 48016 30492
rect 47952 30432 48016 30436
rect 48032 30492 48096 30496
rect 48032 30436 48036 30492
rect 48036 30436 48092 30492
rect 48092 30436 48096 30492
rect 48032 30432 48096 30436
rect 48112 30492 48176 30496
rect 48112 30436 48116 30492
rect 48116 30436 48172 30492
rect 48172 30436 48176 30492
rect 48112 30432 48176 30436
rect 48192 30492 48256 30496
rect 48192 30436 48196 30492
rect 48196 30436 48252 30492
rect 48252 30436 48256 30492
rect 48192 30432 48256 30436
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 32952 29948 33016 29952
rect 32952 29892 32956 29948
rect 32956 29892 33012 29948
rect 33012 29892 33016 29948
rect 32952 29888 33016 29892
rect 33032 29948 33096 29952
rect 33032 29892 33036 29948
rect 33036 29892 33092 29948
rect 33092 29892 33096 29948
rect 33032 29888 33096 29892
rect 33112 29948 33176 29952
rect 33112 29892 33116 29948
rect 33116 29892 33172 29948
rect 33172 29892 33176 29948
rect 33112 29888 33176 29892
rect 33192 29948 33256 29952
rect 33192 29892 33196 29948
rect 33196 29892 33252 29948
rect 33252 29892 33256 29948
rect 33192 29888 33256 29892
rect 42952 29948 43016 29952
rect 42952 29892 42956 29948
rect 42956 29892 43012 29948
rect 43012 29892 43016 29948
rect 42952 29888 43016 29892
rect 43032 29948 43096 29952
rect 43032 29892 43036 29948
rect 43036 29892 43092 29948
rect 43092 29892 43096 29948
rect 43032 29888 43096 29892
rect 43112 29948 43176 29952
rect 43112 29892 43116 29948
rect 43116 29892 43172 29948
rect 43172 29892 43176 29948
rect 43112 29888 43176 29892
rect 43192 29948 43256 29952
rect 43192 29892 43196 29948
rect 43196 29892 43252 29948
rect 43252 29892 43256 29948
rect 43192 29888 43256 29892
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 27952 29404 28016 29408
rect 27952 29348 27956 29404
rect 27956 29348 28012 29404
rect 28012 29348 28016 29404
rect 27952 29344 28016 29348
rect 28032 29404 28096 29408
rect 28032 29348 28036 29404
rect 28036 29348 28092 29404
rect 28092 29348 28096 29404
rect 28032 29344 28096 29348
rect 28112 29404 28176 29408
rect 28112 29348 28116 29404
rect 28116 29348 28172 29404
rect 28172 29348 28176 29404
rect 28112 29344 28176 29348
rect 28192 29404 28256 29408
rect 28192 29348 28196 29404
rect 28196 29348 28252 29404
rect 28252 29348 28256 29404
rect 28192 29344 28256 29348
rect 37952 29404 38016 29408
rect 37952 29348 37956 29404
rect 37956 29348 38012 29404
rect 38012 29348 38016 29404
rect 37952 29344 38016 29348
rect 38032 29404 38096 29408
rect 38032 29348 38036 29404
rect 38036 29348 38092 29404
rect 38092 29348 38096 29404
rect 38032 29344 38096 29348
rect 38112 29404 38176 29408
rect 38112 29348 38116 29404
rect 38116 29348 38172 29404
rect 38172 29348 38176 29404
rect 38112 29344 38176 29348
rect 38192 29404 38256 29408
rect 38192 29348 38196 29404
rect 38196 29348 38252 29404
rect 38252 29348 38256 29404
rect 38192 29344 38256 29348
rect 47952 29404 48016 29408
rect 47952 29348 47956 29404
rect 47956 29348 48012 29404
rect 48012 29348 48016 29404
rect 47952 29344 48016 29348
rect 48032 29404 48096 29408
rect 48032 29348 48036 29404
rect 48036 29348 48092 29404
rect 48092 29348 48096 29404
rect 48032 29344 48096 29348
rect 48112 29404 48176 29408
rect 48112 29348 48116 29404
rect 48116 29348 48172 29404
rect 48172 29348 48176 29404
rect 48112 29344 48176 29348
rect 48192 29404 48256 29408
rect 48192 29348 48196 29404
rect 48196 29348 48252 29404
rect 48252 29348 48256 29404
rect 48192 29344 48256 29348
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 32952 28860 33016 28864
rect 32952 28804 32956 28860
rect 32956 28804 33012 28860
rect 33012 28804 33016 28860
rect 32952 28800 33016 28804
rect 33032 28860 33096 28864
rect 33032 28804 33036 28860
rect 33036 28804 33092 28860
rect 33092 28804 33096 28860
rect 33032 28800 33096 28804
rect 33112 28860 33176 28864
rect 33112 28804 33116 28860
rect 33116 28804 33172 28860
rect 33172 28804 33176 28860
rect 33112 28800 33176 28804
rect 33192 28860 33256 28864
rect 33192 28804 33196 28860
rect 33196 28804 33252 28860
rect 33252 28804 33256 28860
rect 33192 28800 33256 28804
rect 42952 28860 43016 28864
rect 42952 28804 42956 28860
rect 42956 28804 43012 28860
rect 43012 28804 43016 28860
rect 42952 28800 43016 28804
rect 43032 28860 43096 28864
rect 43032 28804 43036 28860
rect 43036 28804 43092 28860
rect 43092 28804 43096 28860
rect 43032 28800 43096 28804
rect 43112 28860 43176 28864
rect 43112 28804 43116 28860
rect 43116 28804 43172 28860
rect 43172 28804 43176 28860
rect 43112 28800 43176 28804
rect 43192 28860 43256 28864
rect 43192 28804 43196 28860
rect 43196 28804 43252 28860
rect 43252 28804 43256 28860
rect 43192 28800 43256 28804
rect 18828 28596 18892 28660
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 27952 28316 28016 28320
rect 27952 28260 27956 28316
rect 27956 28260 28012 28316
rect 28012 28260 28016 28316
rect 27952 28256 28016 28260
rect 28032 28316 28096 28320
rect 28032 28260 28036 28316
rect 28036 28260 28092 28316
rect 28092 28260 28096 28316
rect 28032 28256 28096 28260
rect 28112 28316 28176 28320
rect 28112 28260 28116 28316
rect 28116 28260 28172 28316
rect 28172 28260 28176 28316
rect 28112 28256 28176 28260
rect 28192 28316 28256 28320
rect 28192 28260 28196 28316
rect 28196 28260 28252 28316
rect 28252 28260 28256 28316
rect 28192 28256 28256 28260
rect 37952 28316 38016 28320
rect 37952 28260 37956 28316
rect 37956 28260 38012 28316
rect 38012 28260 38016 28316
rect 37952 28256 38016 28260
rect 38032 28316 38096 28320
rect 38032 28260 38036 28316
rect 38036 28260 38092 28316
rect 38092 28260 38096 28316
rect 38032 28256 38096 28260
rect 38112 28316 38176 28320
rect 38112 28260 38116 28316
rect 38116 28260 38172 28316
rect 38172 28260 38176 28316
rect 38112 28256 38176 28260
rect 38192 28316 38256 28320
rect 38192 28260 38196 28316
rect 38196 28260 38252 28316
rect 38252 28260 38256 28316
rect 38192 28256 38256 28260
rect 47952 28316 48016 28320
rect 47952 28260 47956 28316
rect 47956 28260 48012 28316
rect 48012 28260 48016 28316
rect 47952 28256 48016 28260
rect 48032 28316 48096 28320
rect 48032 28260 48036 28316
rect 48036 28260 48092 28316
rect 48092 28260 48096 28316
rect 48032 28256 48096 28260
rect 48112 28316 48176 28320
rect 48112 28260 48116 28316
rect 48116 28260 48172 28316
rect 48172 28260 48176 28316
rect 48112 28256 48176 28260
rect 48192 28316 48256 28320
rect 48192 28260 48196 28316
rect 48196 28260 48252 28316
rect 48252 28260 48256 28316
rect 48192 28256 48256 28260
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 32952 27772 33016 27776
rect 32952 27716 32956 27772
rect 32956 27716 33012 27772
rect 33012 27716 33016 27772
rect 32952 27712 33016 27716
rect 33032 27772 33096 27776
rect 33032 27716 33036 27772
rect 33036 27716 33092 27772
rect 33092 27716 33096 27772
rect 33032 27712 33096 27716
rect 33112 27772 33176 27776
rect 33112 27716 33116 27772
rect 33116 27716 33172 27772
rect 33172 27716 33176 27772
rect 33112 27712 33176 27716
rect 33192 27772 33256 27776
rect 33192 27716 33196 27772
rect 33196 27716 33252 27772
rect 33252 27716 33256 27772
rect 33192 27712 33256 27716
rect 42952 27772 43016 27776
rect 42952 27716 42956 27772
rect 42956 27716 43012 27772
rect 43012 27716 43016 27772
rect 42952 27712 43016 27716
rect 43032 27772 43096 27776
rect 43032 27716 43036 27772
rect 43036 27716 43092 27772
rect 43092 27716 43096 27772
rect 43032 27712 43096 27716
rect 43112 27772 43176 27776
rect 43112 27716 43116 27772
rect 43116 27716 43172 27772
rect 43172 27716 43176 27772
rect 43112 27712 43176 27716
rect 43192 27772 43256 27776
rect 43192 27716 43196 27772
rect 43196 27716 43252 27772
rect 43252 27716 43256 27772
rect 43192 27712 43256 27716
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 27952 27228 28016 27232
rect 27952 27172 27956 27228
rect 27956 27172 28012 27228
rect 28012 27172 28016 27228
rect 27952 27168 28016 27172
rect 28032 27228 28096 27232
rect 28032 27172 28036 27228
rect 28036 27172 28092 27228
rect 28092 27172 28096 27228
rect 28032 27168 28096 27172
rect 28112 27228 28176 27232
rect 28112 27172 28116 27228
rect 28116 27172 28172 27228
rect 28172 27172 28176 27228
rect 28112 27168 28176 27172
rect 28192 27228 28256 27232
rect 28192 27172 28196 27228
rect 28196 27172 28252 27228
rect 28252 27172 28256 27228
rect 28192 27168 28256 27172
rect 37952 27228 38016 27232
rect 37952 27172 37956 27228
rect 37956 27172 38012 27228
rect 38012 27172 38016 27228
rect 37952 27168 38016 27172
rect 38032 27228 38096 27232
rect 38032 27172 38036 27228
rect 38036 27172 38092 27228
rect 38092 27172 38096 27228
rect 38032 27168 38096 27172
rect 38112 27228 38176 27232
rect 38112 27172 38116 27228
rect 38116 27172 38172 27228
rect 38172 27172 38176 27228
rect 38112 27168 38176 27172
rect 38192 27228 38256 27232
rect 38192 27172 38196 27228
rect 38196 27172 38252 27228
rect 38252 27172 38256 27228
rect 38192 27168 38256 27172
rect 47952 27228 48016 27232
rect 47952 27172 47956 27228
rect 47956 27172 48012 27228
rect 48012 27172 48016 27228
rect 47952 27168 48016 27172
rect 48032 27228 48096 27232
rect 48032 27172 48036 27228
rect 48036 27172 48092 27228
rect 48092 27172 48096 27228
rect 48032 27168 48096 27172
rect 48112 27228 48176 27232
rect 48112 27172 48116 27228
rect 48116 27172 48172 27228
rect 48172 27172 48176 27228
rect 48112 27168 48176 27172
rect 48192 27228 48256 27232
rect 48192 27172 48196 27228
rect 48196 27172 48252 27228
rect 48252 27172 48256 27228
rect 48192 27168 48256 27172
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 32952 26684 33016 26688
rect 32952 26628 32956 26684
rect 32956 26628 33012 26684
rect 33012 26628 33016 26684
rect 32952 26624 33016 26628
rect 33032 26684 33096 26688
rect 33032 26628 33036 26684
rect 33036 26628 33092 26684
rect 33092 26628 33096 26684
rect 33032 26624 33096 26628
rect 33112 26684 33176 26688
rect 33112 26628 33116 26684
rect 33116 26628 33172 26684
rect 33172 26628 33176 26684
rect 33112 26624 33176 26628
rect 33192 26684 33256 26688
rect 33192 26628 33196 26684
rect 33196 26628 33252 26684
rect 33252 26628 33256 26684
rect 33192 26624 33256 26628
rect 42952 26684 43016 26688
rect 42952 26628 42956 26684
rect 42956 26628 43012 26684
rect 43012 26628 43016 26684
rect 42952 26624 43016 26628
rect 43032 26684 43096 26688
rect 43032 26628 43036 26684
rect 43036 26628 43092 26684
rect 43092 26628 43096 26684
rect 43032 26624 43096 26628
rect 43112 26684 43176 26688
rect 43112 26628 43116 26684
rect 43116 26628 43172 26684
rect 43172 26628 43176 26684
rect 43112 26624 43176 26628
rect 43192 26684 43256 26688
rect 43192 26628 43196 26684
rect 43196 26628 43252 26684
rect 43252 26628 43256 26684
rect 43192 26624 43256 26628
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 27952 26140 28016 26144
rect 27952 26084 27956 26140
rect 27956 26084 28012 26140
rect 28012 26084 28016 26140
rect 27952 26080 28016 26084
rect 28032 26140 28096 26144
rect 28032 26084 28036 26140
rect 28036 26084 28092 26140
rect 28092 26084 28096 26140
rect 28032 26080 28096 26084
rect 28112 26140 28176 26144
rect 28112 26084 28116 26140
rect 28116 26084 28172 26140
rect 28172 26084 28176 26140
rect 28112 26080 28176 26084
rect 28192 26140 28256 26144
rect 28192 26084 28196 26140
rect 28196 26084 28252 26140
rect 28252 26084 28256 26140
rect 28192 26080 28256 26084
rect 37952 26140 38016 26144
rect 37952 26084 37956 26140
rect 37956 26084 38012 26140
rect 38012 26084 38016 26140
rect 37952 26080 38016 26084
rect 38032 26140 38096 26144
rect 38032 26084 38036 26140
rect 38036 26084 38092 26140
rect 38092 26084 38096 26140
rect 38032 26080 38096 26084
rect 38112 26140 38176 26144
rect 38112 26084 38116 26140
rect 38116 26084 38172 26140
rect 38172 26084 38176 26140
rect 38112 26080 38176 26084
rect 38192 26140 38256 26144
rect 38192 26084 38196 26140
rect 38196 26084 38252 26140
rect 38252 26084 38256 26140
rect 38192 26080 38256 26084
rect 47952 26140 48016 26144
rect 47952 26084 47956 26140
rect 47956 26084 48012 26140
rect 48012 26084 48016 26140
rect 47952 26080 48016 26084
rect 48032 26140 48096 26144
rect 48032 26084 48036 26140
rect 48036 26084 48092 26140
rect 48092 26084 48096 26140
rect 48032 26080 48096 26084
rect 48112 26140 48176 26144
rect 48112 26084 48116 26140
rect 48116 26084 48172 26140
rect 48172 26084 48176 26140
rect 48112 26080 48176 26084
rect 48192 26140 48256 26144
rect 48192 26084 48196 26140
rect 48196 26084 48252 26140
rect 48252 26084 48256 26140
rect 48192 26080 48256 26084
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 32952 25596 33016 25600
rect 32952 25540 32956 25596
rect 32956 25540 33012 25596
rect 33012 25540 33016 25596
rect 32952 25536 33016 25540
rect 33032 25596 33096 25600
rect 33032 25540 33036 25596
rect 33036 25540 33092 25596
rect 33092 25540 33096 25596
rect 33032 25536 33096 25540
rect 33112 25596 33176 25600
rect 33112 25540 33116 25596
rect 33116 25540 33172 25596
rect 33172 25540 33176 25596
rect 33112 25536 33176 25540
rect 33192 25596 33256 25600
rect 33192 25540 33196 25596
rect 33196 25540 33252 25596
rect 33252 25540 33256 25596
rect 33192 25536 33256 25540
rect 42952 25596 43016 25600
rect 42952 25540 42956 25596
rect 42956 25540 43012 25596
rect 43012 25540 43016 25596
rect 42952 25536 43016 25540
rect 43032 25596 43096 25600
rect 43032 25540 43036 25596
rect 43036 25540 43092 25596
rect 43092 25540 43096 25596
rect 43032 25536 43096 25540
rect 43112 25596 43176 25600
rect 43112 25540 43116 25596
rect 43116 25540 43172 25596
rect 43172 25540 43176 25596
rect 43112 25536 43176 25540
rect 43192 25596 43256 25600
rect 43192 25540 43196 25596
rect 43196 25540 43252 25596
rect 43252 25540 43256 25596
rect 43192 25536 43256 25540
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 27952 25052 28016 25056
rect 27952 24996 27956 25052
rect 27956 24996 28012 25052
rect 28012 24996 28016 25052
rect 27952 24992 28016 24996
rect 28032 25052 28096 25056
rect 28032 24996 28036 25052
rect 28036 24996 28092 25052
rect 28092 24996 28096 25052
rect 28032 24992 28096 24996
rect 28112 25052 28176 25056
rect 28112 24996 28116 25052
rect 28116 24996 28172 25052
rect 28172 24996 28176 25052
rect 28112 24992 28176 24996
rect 28192 25052 28256 25056
rect 28192 24996 28196 25052
rect 28196 24996 28252 25052
rect 28252 24996 28256 25052
rect 28192 24992 28256 24996
rect 37952 25052 38016 25056
rect 37952 24996 37956 25052
rect 37956 24996 38012 25052
rect 38012 24996 38016 25052
rect 37952 24992 38016 24996
rect 38032 25052 38096 25056
rect 38032 24996 38036 25052
rect 38036 24996 38092 25052
rect 38092 24996 38096 25052
rect 38032 24992 38096 24996
rect 38112 25052 38176 25056
rect 38112 24996 38116 25052
rect 38116 24996 38172 25052
rect 38172 24996 38176 25052
rect 38112 24992 38176 24996
rect 38192 25052 38256 25056
rect 38192 24996 38196 25052
rect 38196 24996 38252 25052
rect 38252 24996 38256 25052
rect 38192 24992 38256 24996
rect 47952 25052 48016 25056
rect 47952 24996 47956 25052
rect 47956 24996 48012 25052
rect 48012 24996 48016 25052
rect 47952 24992 48016 24996
rect 48032 25052 48096 25056
rect 48032 24996 48036 25052
rect 48036 24996 48092 25052
rect 48092 24996 48096 25052
rect 48032 24992 48096 24996
rect 48112 25052 48176 25056
rect 48112 24996 48116 25052
rect 48116 24996 48172 25052
rect 48172 24996 48176 25052
rect 48112 24992 48176 24996
rect 48192 25052 48256 25056
rect 48192 24996 48196 25052
rect 48196 24996 48252 25052
rect 48252 24996 48256 25052
rect 48192 24992 48256 24996
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 7236 20300 7300 20364
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 9444 17716 9508 17780
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 10916 17036 10980 17100
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 11099 54092 11165 54093
rect 11099 54028 11100 54092
rect 11164 54028 11165 54092
rect 11099 54027 11165 54028
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 9259 43212 9325 43213
rect 9259 43148 9260 43212
rect 9324 43148 9325 43212
rect 9259 43147 9325 43148
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7235 36684 7301 36685
rect 7235 36620 7236 36684
rect 7300 36620 7301 36684
rect 7235 36619 7301 36620
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 7238 20365 7298 36619
rect 7944 35936 8264 36960
rect 9262 36957 9322 43147
rect 10731 40900 10797 40901
rect 10731 40836 10732 40900
rect 10796 40836 10797 40900
rect 10731 40835 10797 40836
rect 9259 36956 9325 36957
rect 9259 36892 9260 36956
rect 9324 36892 9325 36956
rect 9259 36891 9325 36892
rect 9443 36684 9509 36685
rect 9443 36620 9444 36684
rect 9508 36620 9509 36684
rect 9443 36619 9509 36620
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7235 20364 7301 20365
rect 7235 20300 7236 20364
rect 7300 20300 7301 20364
rect 7235 20299 7301 20300
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 9446 17781 9506 36619
rect 10734 33149 10794 40835
rect 10915 38180 10981 38181
rect 10915 38116 10916 38180
rect 10980 38116 10981 38180
rect 10915 38115 10981 38116
rect 10731 33148 10797 33149
rect 10731 33084 10732 33148
rect 10796 33084 10797 33148
rect 10731 33083 10797 33084
rect 9443 17780 9509 17781
rect 9443 17716 9444 17780
rect 9508 17716 9509 17780
rect 9443 17715 9509 17716
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 10918 17101 10978 38115
rect 11102 37229 11162 54027
rect 12944 53888 13264 54448
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 11099 37228 11165 37229
rect 11099 37164 11100 37228
rect 11164 37164 11165 37228
rect 11099 37163 11165 37164
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 10915 17100 10981 17101
rect 10915 17036 10916 17100
rect 10980 17036 10981 17100
rect 10915 17035 10981 17036
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 17944 53344 18264 54368
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 22944 53888 23264 54448
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 18827 41988 18893 41989
rect 18827 41924 18828 41988
rect 18892 41924 18893 41988
rect 18827 41923 18893 41924
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17944 38112 18264 39136
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 18830 28661 18890 41923
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 18827 28660 18893 28661
rect 18827 28596 18828 28660
rect 18892 28596 18893 28660
rect 18827 28595 18893 28596
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17944 27232 18264 28256
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 27944 54432 28264 54448
rect 27944 54368 27952 54432
rect 28016 54368 28032 54432
rect 28096 54368 28112 54432
rect 28176 54368 28192 54432
rect 28256 54368 28264 54432
rect 27944 53344 28264 54368
rect 27944 53280 27952 53344
rect 28016 53280 28032 53344
rect 28096 53280 28112 53344
rect 28176 53280 28192 53344
rect 28256 53280 28264 53344
rect 27944 52256 28264 53280
rect 27944 52192 27952 52256
rect 28016 52192 28032 52256
rect 28096 52192 28112 52256
rect 28176 52192 28192 52256
rect 28256 52192 28264 52256
rect 27944 51168 28264 52192
rect 27944 51104 27952 51168
rect 28016 51104 28032 51168
rect 28096 51104 28112 51168
rect 28176 51104 28192 51168
rect 28256 51104 28264 51168
rect 27944 50080 28264 51104
rect 27944 50016 27952 50080
rect 28016 50016 28032 50080
rect 28096 50016 28112 50080
rect 28176 50016 28192 50080
rect 28256 50016 28264 50080
rect 27944 48992 28264 50016
rect 27944 48928 27952 48992
rect 28016 48928 28032 48992
rect 28096 48928 28112 48992
rect 28176 48928 28192 48992
rect 28256 48928 28264 48992
rect 27944 47904 28264 48928
rect 27944 47840 27952 47904
rect 28016 47840 28032 47904
rect 28096 47840 28112 47904
rect 28176 47840 28192 47904
rect 28256 47840 28264 47904
rect 27944 46816 28264 47840
rect 27944 46752 27952 46816
rect 28016 46752 28032 46816
rect 28096 46752 28112 46816
rect 28176 46752 28192 46816
rect 28256 46752 28264 46816
rect 27944 45728 28264 46752
rect 27944 45664 27952 45728
rect 28016 45664 28032 45728
rect 28096 45664 28112 45728
rect 28176 45664 28192 45728
rect 28256 45664 28264 45728
rect 27944 44640 28264 45664
rect 27944 44576 27952 44640
rect 28016 44576 28032 44640
rect 28096 44576 28112 44640
rect 28176 44576 28192 44640
rect 28256 44576 28264 44640
rect 27944 43552 28264 44576
rect 27944 43488 27952 43552
rect 28016 43488 28032 43552
rect 28096 43488 28112 43552
rect 28176 43488 28192 43552
rect 28256 43488 28264 43552
rect 27944 42464 28264 43488
rect 27944 42400 27952 42464
rect 28016 42400 28032 42464
rect 28096 42400 28112 42464
rect 28176 42400 28192 42464
rect 28256 42400 28264 42464
rect 27944 41376 28264 42400
rect 27944 41312 27952 41376
rect 28016 41312 28032 41376
rect 28096 41312 28112 41376
rect 28176 41312 28192 41376
rect 28256 41312 28264 41376
rect 27944 40288 28264 41312
rect 27944 40224 27952 40288
rect 28016 40224 28032 40288
rect 28096 40224 28112 40288
rect 28176 40224 28192 40288
rect 28256 40224 28264 40288
rect 27944 39200 28264 40224
rect 27944 39136 27952 39200
rect 28016 39136 28032 39200
rect 28096 39136 28112 39200
rect 28176 39136 28192 39200
rect 28256 39136 28264 39200
rect 27944 38112 28264 39136
rect 27944 38048 27952 38112
rect 28016 38048 28032 38112
rect 28096 38048 28112 38112
rect 28176 38048 28192 38112
rect 28256 38048 28264 38112
rect 27944 37024 28264 38048
rect 27944 36960 27952 37024
rect 28016 36960 28032 37024
rect 28096 36960 28112 37024
rect 28176 36960 28192 37024
rect 28256 36960 28264 37024
rect 27944 35936 28264 36960
rect 27944 35872 27952 35936
rect 28016 35872 28032 35936
rect 28096 35872 28112 35936
rect 28176 35872 28192 35936
rect 28256 35872 28264 35936
rect 27944 34848 28264 35872
rect 27944 34784 27952 34848
rect 28016 34784 28032 34848
rect 28096 34784 28112 34848
rect 28176 34784 28192 34848
rect 28256 34784 28264 34848
rect 27944 33760 28264 34784
rect 27944 33696 27952 33760
rect 28016 33696 28032 33760
rect 28096 33696 28112 33760
rect 28176 33696 28192 33760
rect 28256 33696 28264 33760
rect 27944 32672 28264 33696
rect 27944 32608 27952 32672
rect 28016 32608 28032 32672
rect 28096 32608 28112 32672
rect 28176 32608 28192 32672
rect 28256 32608 28264 32672
rect 27944 31584 28264 32608
rect 27944 31520 27952 31584
rect 28016 31520 28032 31584
rect 28096 31520 28112 31584
rect 28176 31520 28192 31584
rect 28256 31520 28264 31584
rect 27944 30496 28264 31520
rect 27944 30432 27952 30496
rect 28016 30432 28032 30496
rect 28096 30432 28112 30496
rect 28176 30432 28192 30496
rect 28256 30432 28264 30496
rect 27944 29408 28264 30432
rect 27944 29344 27952 29408
rect 28016 29344 28032 29408
rect 28096 29344 28112 29408
rect 28176 29344 28192 29408
rect 28256 29344 28264 29408
rect 27944 28320 28264 29344
rect 27944 28256 27952 28320
rect 28016 28256 28032 28320
rect 28096 28256 28112 28320
rect 28176 28256 28192 28320
rect 28256 28256 28264 28320
rect 27944 27232 28264 28256
rect 27944 27168 27952 27232
rect 28016 27168 28032 27232
rect 28096 27168 28112 27232
rect 28176 27168 28192 27232
rect 28256 27168 28264 27232
rect 27944 26144 28264 27168
rect 27944 26080 27952 26144
rect 28016 26080 28032 26144
rect 28096 26080 28112 26144
rect 28176 26080 28192 26144
rect 28256 26080 28264 26144
rect 27944 25056 28264 26080
rect 27944 24992 27952 25056
rect 28016 24992 28032 25056
rect 28096 24992 28112 25056
rect 28176 24992 28192 25056
rect 28256 24992 28264 25056
rect 27944 23968 28264 24992
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27944 18528 28264 19552
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27944 17440 28264 18464
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27944 14176 28264 15200
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 53888 33264 54448
rect 32944 53824 32952 53888
rect 33016 53824 33032 53888
rect 33096 53824 33112 53888
rect 33176 53824 33192 53888
rect 33256 53824 33264 53888
rect 32944 52800 33264 53824
rect 32944 52736 32952 52800
rect 33016 52736 33032 52800
rect 33096 52736 33112 52800
rect 33176 52736 33192 52800
rect 33256 52736 33264 52800
rect 32944 51712 33264 52736
rect 32944 51648 32952 51712
rect 33016 51648 33032 51712
rect 33096 51648 33112 51712
rect 33176 51648 33192 51712
rect 33256 51648 33264 51712
rect 32944 50624 33264 51648
rect 32944 50560 32952 50624
rect 33016 50560 33032 50624
rect 33096 50560 33112 50624
rect 33176 50560 33192 50624
rect 33256 50560 33264 50624
rect 32944 49536 33264 50560
rect 32944 49472 32952 49536
rect 33016 49472 33032 49536
rect 33096 49472 33112 49536
rect 33176 49472 33192 49536
rect 33256 49472 33264 49536
rect 32944 48448 33264 49472
rect 32944 48384 32952 48448
rect 33016 48384 33032 48448
rect 33096 48384 33112 48448
rect 33176 48384 33192 48448
rect 33256 48384 33264 48448
rect 32944 47360 33264 48384
rect 32944 47296 32952 47360
rect 33016 47296 33032 47360
rect 33096 47296 33112 47360
rect 33176 47296 33192 47360
rect 33256 47296 33264 47360
rect 32944 46272 33264 47296
rect 32944 46208 32952 46272
rect 33016 46208 33032 46272
rect 33096 46208 33112 46272
rect 33176 46208 33192 46272
rect 33256 46208 33264 46272
rect 32944 45184 33264 46208
rect 32944 45120 32952 45184
rect 33016 45120 33032 45184
rect 33096 45120 33112 45184
rect 33176 45120 33192 45184
rect 33256 45120 33264 45184
rect 32944 44096 33264 45120
rect 32944 44032 32952 44096
rect 33016 44032 33032 44096
rect 33096 44032 33112 44096
rect 33176 44032 33192 44096
rect 33256 44032 33264 44096
rect 32944 43008 33264 44032
rect 32944 42944 32952 43008
rect 33016 42944 33032 43008
rect 33096 42944 33112 43008
rect 33176 42944 33192 43008
rect 33256 42944 33264 43008
rect 32944 41920 33264 42944
rect 32944 41856 32952 41920
rect 33016 41856 33032 41920
rect 33096 41856 33112 41920
rect 33176 41856 33192 41920
rect 33256 41856 33264 41920
rect 32944 40832 33264 41856
rect 32944 40768 32952 40832
rect 33016 40768 33032 40832
rect 33096 40768 33112 40832
rect 33176 40768 33192 40832
rect 33256 40768 33264 40832
rect 32944 39744 33264 40768
rect 32944 39680 32952 39744
rect 33016 39680 33032 39744
rect 33096 39680 33112 39744
rect 33176 39680 33192 39744
rect 33256 39680 33264 39744
rect 32944 38656 33264 39680
rect 32944 38592 32952 38656
rect 33016 38592 33032 38656
rect 33096 38592 33112 38656
rect 33176 38592 33192 38656
rect 33256 38592 33264 38656
rect 32944 37568 33264 38592
rect 32944 37504 32952 37568
rect 33016 37504 33032 37568
rect 33096 37504 33112 37568
rect 33176 37504 33192 37568
rect 33256 37504 33264 37568
rect 32944 36480 33264 37504
rect 32944 36416 32952 36480
rect 33016 36416 33032 36480
rect 33096 36416 33112 36480
rect 33176 36416 33192 36480
rect 33256 36416 33264 36480
rect 32944 35392 33264 36416
rect 32944 35328 32952 35392
rect 33016 35328 33032 35392
rect 33096 35328 33112 35392
rect 33176 35328 33192 35392
rect 33256 35328 33264 35392
rect 32944 34304 33264 35328
rect 32944 34240 32952 34304
rect 33016 34240 33032 34304
rect 33096 34240 33112 34304
rect 33176 34240 33192 34304
rect 33256 34240 33264 34304
rect 32944 33216 33264 34240
rect 32944 33152 32952 33216
rect 33016 33152 33032 33216
rect 33096 33152 33112 33216
rect 33176 33152 33192 33216
rect 33256 33152 33264 33216
rect 32944 32128 33264 33152
rect 32944 32064 32952 32128
rect 33016 32064 33032 32128
rect 33096 32064 33112 32128
rect 33176 32064 33192 32128
rect 33256 32064 33264 32128
rect 32944 31040 33264 32064
rect 32944 30976 32952 31040
rect 33016 30976 33032 31040
rect 33096 30976 33112 31040
rect 33176 30976 33192 31040
rect 33256 30976 33264 31040
rect 32944 29952 33264 30976
rect 32944 29888 32952 29952
rect 33016 29888 33032 29952
rect 33096 29888 33112 29952
rect 33176 29888 33192 29952
rect 33256 29888 33264 29952
rect 32944 28864 33264 29888
rect 32944 28800 32952 28864
rect 33016 28800 33032 28864
rect 33096 28800 33112 28864
rect 33176 28800 33192 28864
rect 33256 28800 33264 28864
rect 32944 27776 33264 28800
rect 32944 27712 32952 27776
rect 33016 27712 33032 27776
rect 33096 27712 33112 27776
rect 33176 27712 33192 27776
rect 33256 27712 33264 27776
rect 32944 26688 33264 27712
rect 32944 26624 32952 26688
rect 33016 26624 33032 26688
rect 33096 26624 33112 26688
rect 33176 26624 33192 26688
rect 33256 26624 33264 26688
rect 32944 25600 33264 26624
rect 32944 25536 32952 25600
rect 33016 25536 33032 25600
rect 33096 25536 33112 25600
rect 33176 25536 33192 25600
rect 33256 25536 33264 25600
rect 32944 24512 33264 25536
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 32944 19072 33264 20096
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32944 10368 33264 11392
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 54432 38264 54448
rect 37944 54368 37952 54432
rect 38016 54368 38032 54432
rect 38096 54368 38112 54432
rect 38176 54368 38192 54432
rect 38256 54368 38264 54432
rect 37944 53344 38264 54368
rect 37944 53280 37952 53344
rect 38016 53280 38032 53344
rect 38096 53280 38112 53344
rect 38176 53280 38192 53344
rect 38256 53280 38264 53344
rect 37944 52256 38264 53280
rect 37944 52192 37952 52256
rect 38016 52192 38032 52256
rect 38096 52192 38112 52256
rect 38176 52192 38192 52256
rect 38256 52192 38264 52256
rect 37944 51168 38264 52192
rect 37944 51104 37952 51168
rect 38016 51104 38032 51168
rect 38096 51104 38112 51168
rect 38176 51104 38192 51168
rect 38256 51104 38264 51168
rect 37944 50080 38264 51104
rect 37944 50016 37952 50080
rect 38016 50016 38032 50080
rect 38096 50016 38112 50080
rect 38176 50016 38192 50080
rect 38256 50016 38264 50080
rect 37944 48992 38264 50016
rect 37944 48928 37952 48992
rect 38016 48928 38032 48992
rect 38096 48928 38112 48992
rect 38176 48928 38192 48992
rect 38256 48928 38264 48992
rect 37944 47904 38264 48928
rect 37944 47840 37952 47904
rect 38016 47840 38032 47904
rect 38096 47840 38112 47904
rect 38176 47840 38192 47904
rect 38256 47840 38264 47904
rect 37944 46816 38264 47840
rect 37944 46752 37952 46816
rect 38016 46752 38032 46816
rect 38096 46752 38112 46816
rect 38176 46752 38192 46816
rect 38256 46752 38264 46816
rect 37944 45728 38264 46752
rect 37944 45664 37952 45728
rect 38016 45664 38032 45728
rect 38096 45664 38112 45728
rect 38176 45664 38192 45728
rect 38256 45664 38264 45728
rect 37944 44640 38264 45664
rect 37944 44576 37952 44640
rect 38016 44576 38032 44640
rect 38096 44576 38112 44640
rect 38176 44576 38192 44640
rect 38256 44576 38264 44640
rect 37944 43552 38264 44576
rect 37944 43488 37952 43552
rect 38016 43488 38032 43552
rect 38096 43488 38112 43552
rect 38176 43488 38192 43552
rect 38256 43488 38264 43552
rect 37944 42464 38264 43488
rect 37944 42400 37952 42464
rect 38016 42400 38032 42464
rect 38096 42400 38112 42464
rect 38176 42400 38192 42464
rect 38256 42400 38264 42464
rect 37944 41376 38264 42400
rect 37944 41312 37952 41376
rect 38016 41312 38032 41376
rect 38096 41312 38112 41376
rect 38176 41312 38192 41376
rect 38256 41312 38264 41376
rect 37944 40288 38264 41312
rect 37944 40224 37952 40288
rect 38016 40224 38032 40288
rect 38096 40224 38112 40288
rect 38176 40224 38192 40288
rect 38256 40224 38264 40288
rect 37944 39200 38264 40224
rect 37944 39136 37952 39200
rect 38016 39136 38032 39200
rect 38096 39136 38112 39200
rect 38176 39136 38192 39200
rect 38256 39136 38264 39200
rect 37944 38112 38264 39136
rect 37944 38048 37952 38112
rect 38016 38048 38032 38112
rect 38096 38048 38112 38112
rect 38176 38048 38192 38112
rect 38256 38048 38264 38112
rect 37944 37024 38264 38048
rect 37944 36960 37952 37024
rect 38016 36960 38032 37024
rect 38096 36960 38112 37024
rect 38176 36960 38192 37024
rect 38256 36960 38264 37024
rect 37944 35936 38264 36960
rect 37944 35872 37952 35936
rect 38016 35872 38032 35936
rect 38096 35872 38112 35936
rect 38176 35872 38192 35936
rect 38256 35872 38264 35936
rect 37944 34848 38264 35872
rect 37944 34784 37952 34848
rect 38016 34784 38032 34848
rect 38096 34784 38112 34848
rect 38176 34784 38192 34848
rect 38256 34784 38264 34848
rect 37944 33760 38264 34784
rect 37944 33696 37952 33760
rect 38016 33696 38032 33760
rect 38096 33696 38112 33760
rect 38176 33696 38192 33760
rect 38256 33696 38264 33760
rect 37944 32672 38264 33696
rect 37944 32608 37952 32672
rect 38016 32608 38032 32672
rect 38096 32608 38112 32672
rect 38176 32608 38192 32672
rect 38256 32608 38264 32672
rect 37944 31584 38264 32608
rect 37944 31520 37952 31584
rect 38016 31520 38032 31584
rect 38096 31520 38112 31584
rect 38176 31520 38192 31584
rect 38256 31520 38264 31584
rect 37944 30496 38264 31520
rect 37944 30432 37952 30496
rect 38016 30432 38032 30496
rect 38096 30432 38112 30496
rect 38176 30432 38192 30496
rect 38256 30432 38264 30496
rect 37944 29408 38264 30432
rect 37944 29344 37952 29408
rect 38016 29344 38032 29408
rect 38096 29344 38112 29408
rect 38176 29344 38192 29408
rect 38256 29344 38264 29408
rect 37944 28320 38264 29344
rect 37944 28256 37952 28320
rect 38016 28256 38032 28320
rect 38096 28256 38112 28320
rect 38176 28256 38192 28320
rect 38256 28256 38264 28320
rect 37944 27232 38264 28256
rect 37944 27168 37952 27232
rect 38016 27168 38032 27232
rect 38096 27168 38112 27232
rect 38176 27168 38192 27232
rect 38256 27168 38264 27232
rect 37944 26144 38264 27168
rect 37944 26080 37952 26144
rect 38016 26080 38032 26144
rect 38096 26080 38112 26144
rect 38176 26080 38192 26144
rect 38256 26080 38264 26144
rect 37944 25056 38264 26080
rect 37944 24992 37952 25056
rect 38016 24992 38032 25056
rect 38096 24992 38112 25056
rect 38176 24992 38192 25056
rect 38256 24992 38264 25056
rect 37944 23968 38264 24992
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 53888 43264 54448
rect 42944 53824 42952 53888
rect 43016 53824 43032 53888
rect 43096 53824 43112 53888
rect 43176 53824 43192 53888
rect 43256 53824 43264 53888
rect 42944 52800 43264 53824
rect 42944 52736 42952 52800
rect 43016 52736 43032 52800
rect 43096 52736 43112 52800
rect 43176 52736 43192 52800
rect 43256 52736 43264 52800
rect 42944 51712 43264 52736
rect 42944 51648 42952 51712
rect 43016 51648 43032 51712
rect 43096 51648 43112 51712
rect 43176 51648 43192 51712
rect 43256 51648 43264 51712
rect 42944 50624 43264 51648
rect 42944 50560 42952 50624
rect 43016 50560 43032 50624
rect 43096 50560 43112 50624
rect 43176 50560 43192 50624
rect 43256 50560 43264 50624
rect 42944 49536 43264 50560
rect 42944 49472 42952 49536
rect 43016 49472 43032 49536
rect 43096 49472 43112 49536
rect 43176 49472 43192 49536
rect 43256 49472 43264 49536
rect 42944 48448 43264 49472
rect 42944 48384 42952 48448
rect 43016 48384 43032 48448
rect 43096 48384 43112 48448
rect 43176 48384 43192 48448
rect 43256 48384 43264 48448
rect 42944 47360 43264 48384
rect 42944 47296 42952 47360
rect 43016 47296 43032 47360
rect 43096 47296 43112 47360
rect 43176 47296 43192 47360
rect 43256 47296 43264 47360
rect 42944 46272 43264 47296
rect 42944 46208 42952 46272
rect 43016 46208 43032 46272
rect 43096 46208 43112 46272
rect 43176 46208 43192 46272
rect 43256 46208 43264 46272
rect 42944 45184 43264 46208
rect 42944 45120 42952 45184
rect 43016 45120 43032 45184
rect 43096 45120 43112 45184
rect 43176 45120 43192 45184
rect 43256 45120 43264 45184
rect 42944 44096 43264 45120
rect 42944 44032 42952 44096
rect 43016 44032 43032 44096
rect 43096 44032 43112 44096
rect 43176 44032 43192 44096
rect 43256 44032 43264 44096
rect 42944 43008 43264 44032
rect 42944 42944 42952 43008
rect 43016 42944 43032 43008
rect 43096 42944 43112 43008
rect 43176 42944 43192 43008
rect 43256 42944 43264 43008
rect 42944 41920 43264 42944
rect 42944 41856 42952 41920
rect 43016 41856 43032 41920
rect 43096 41856 43112 41920
rect 43176 41856 43192 41920
rect 43256 41856 43264 41920
rect 42944 40832 43264 41856
rect 42944 40768 42952 40832
rect 43016 40768 43032 40832
rect 43096 40768 43112 40832
rect 43176 40768 43192 40832
rect 43256 40768 43264 40832
rect 42944 39744 43264 40768
rect 42944 39680 42952 39744
rect 43016 39680 43032 39744
rect 43096 39680 43112 39744
rect 43176 39680 43192 39744
rect 43256 39680 43264 39744
rect 42944 38656 43264 39680
rect 42944 38592 42952 38656
rect 43016 38592 43032 38656
rect 43096 38592 43112 38656
rect 43176 38592 43192 38656
rect 43256 38592 43264 38656
rect 42944 37568 43264 38592
rect 42944 37504 42952 37568
rect 43016 37504 43032 37568
rect 43096 37504 43112 37568
rect 43176 37504 43192 37568
rect 43256 37504 43264 37568
rect 42944 36480 43264 37504
rect 42944 36416 42952 36480
rect 43016 36416 43032 36480
rect 43096 36416 43112 36480
rect 43176 36416 43192 36480
rect 43256 36416 43264 36480
rect 42944 35392 43264 36416
rect 42944 35328 42952 35392
rect 43016 35328 43032 35392
rect 43096 35328 43112 35392
rect 43176 35328 43192 35392
rect 43256 35328 43264 35392
rect 42944 34304 43264 35328
rect 42944 34240 42952 34304
rect 43016 34240 43032 34304
rect 43096 34240 43112 34304
rect 43176 34240 43192 34304
rect 43256 34240 43264 34304
rect 42944 33216 43264 34240
rect 42944 33152 42952 33216
rect 43016 33152 43032 33216
rect 43096 33152 43112 33216
rect 43176 33152 43192 33216
rect 43256 33152 43264 33216
rect 42944 32128 43264 33152
rect 42944 32064 42952 32128
rect 43016 32064 43032 32128
rect 43096 32064 43112 32128
rect 43176 32064 43192 32128
rect 43256 32064 43264 32128
rect 42944 31040 43264 32064
rect 42944 30976 42952 31040
rect 43016 30976 43032 31040
rect 43096 30976 43112 31040
rect 43176 30976 43192 31040
rect 43256 30976 43264 31040
rect 42944 29952 43264 30976
rect 42944 29888 42952 29952
rect 43016 29888 43032 29952
rect 43096 29888 43112 29952
rect 43176 29888 43192 29952
rect 43256 29888 43264 29952
rect 42944 28864 43264 29888
rect 42944 28800 42952 28864
rect 43016 28800 43032 28864
rect 43096 28800 43112 28864
rect 43176 28800 43192 28864
rect 43256 28800 43264 28864
rect 42944 27776 43264 28800
rect 42944 27712 42952 27776
rect 43016 27712 43032 27776
rect 43096 27712 43112 27776
rect 43176 27712 43192 27776
rect 43256 27712 43264 27776
rect 42944 26688 43264 27712
rect 42944 26624 42952 26688
rect 43016 26624 43032 26688
rect 43096 26624 43112 26688
rect 43176 26624 43192 26688
rect 43256 26624 43264 26688
rect 42944 25600 43264 26624
rect 42944 25536 42952 25600
rect 43016 25536 43032 25600
rect 43096 25536 43112 25600
rect 43176 25536 43192 25600
rect 43256 25536 43264 25600
rect 42944 24512 43264 25536
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 54432 48264 54448
rect 47944 54368 47952 54432
rect 48016 54368 48032 54432
rect 48096 54368 48112 54432
rect 48176 54368 48192 54432
rect 48256 54368 48264 54432
rect 47944 53344 48264 54368
rect 47944 53280 47952 53344
rect 48016 53280 48032 53344
rect 48096 53280 48112 53344
rect 48176 53280 48192 53344
rect 48256 53280 48264 53344
rect 47944 52256 48264 53280
rect 47944 52192 47952 52256
rect 48016 52192 48032 52256
rect 48096 52192 48112 52256
rect 48176 52192 48192 52256
rect 48256 52192 48264 52256
rect 47944 51168 48264 52192
rect 47944 51104 47952 51168
rect 48016 51104 48032 51168
rect 48096 51104 48112 51168
rect 48176 51104 48192 51168
rect 48256 51104 48264 51168
rect 47944 50080 48264 51104
rect 47944 50016 47952 50080
rect 48016 50016 48032 50080
rect 48096 50016 48112 50080
rect 48176 50016 48192 50080
rect 48256 50016 48264 50080
rect 47944 48992 48264 50016
rect 47944 48928 47952 48992
rect 48016 48928 48032 48992
rect 48096 48928 48112 48992
rect 48176 48928 48192 48992
rect 48256 48928 48264 48992
rect 47944 47904 48264 48928
rect 47944 47840 47952 47904
rect 48016 47840 48032 47904
rect 48096 47840 48112 47904
rect 48176 47840 48192 47904
rect 48256 47840 48264 47904
rect 47944 46816 48264 47840
rect 47944 46752 47952 46816
rect 48016 46752 48032 46816
rect 48096 46752 48112 46816
rect 48176 46752 48192 46816
rect 48256 46752 48264 46816
rect 47944 45728 48264 46752
rect 47944 45664 47952 45728
rect 48016 45664 48032 45728
rect 48096 45664 48112 45728
rect 48176 45664 48192 45728
rect 48256 45664 48264 45728
rect 47944 44640 48264 45664
rect 47944 44576 47952 44640
rect 48016 44576 48032 44640
rect 48096 44576 48112 44640
rect 48176 44576 48192 44640
rect 48256 44576 48264 44640
rect 47944 43552 48264 44576
rect 47944 43488 47952 43552
rect 48016 43488 48032 43552
rect 48096 43488 48112 43552
rect 48176 43488 48192 43552
rect 48256 43488 48264 43552
rect 47944 42464 48264 43488
rect 47944 42400 47952 42464
rect 48016 42400 48032 42464
rect 48096 42400 48112 42464
rect 48176 42400 48192 42464
rect 48256 42400 48264 42464
rect 47944 41376 48264 42400
rect 47944 41312 47952 41376
rect 48016 41312 48032 41376
rect 48096 41312 48112 41376
rect 48176 41312 48192 41376
rect 48256 41312 48264 41376
rect 47944 40288 48264 41312
rect 47944 40224 47952 40288
rect 48016 40224 48032 40288
rect 48096 40224 48112 40288
rect 48176 40224 48192 40288
rect 48256 40224 48264 40288
rect 47944 39200 48264 40224
rect 47944 39136 47952 39200
rect 48016 39136 48032 39200
rect 48096 39136 48112 39200
rect 48176 39136 48192 39200
rect 48256 39136 48264 39200
rect 47944 38112 48264 39136
rect 47944 38048 47952 38112
rect 48016 38048 48032 38112
rect 48096 38048 48112 38112
rect 48176 38048 48192 38112
rect 48256 38048 48264 38112
rect 47944 37024 48264 38048
rect 47944 36960 47952 37024
rect 48016 36960 48032 37024
rect 48096 36960 48112 37024
rect 48176 36960 48192 37024
rect 48256 36960 48264 37024
rect 47944 35936 48264 36960
rect 47944 35872 47952 35936
rect 48016 35872 48032 35936
rect 48096 35872 48112 35936
rect 48176 35872 48192 35936
rect 48256 35872 48264 35936
rect 47944 34848 48264 35872
rect 47944 34784 47952 34848
rect 48016 34784 48032 34848
rect 48096 34784 48112 34848
rect 48176 34784 48192 34848
rect 48256 34784 48264 34848
rect 47944 33760 48264 34784
rect 47944 33696 47952 33760
rect 48016 33696 48032 33760
rect 48096 33696 48112 33760
rect 48176 33696 48192 33760
rect 48256 33696 48264 33760
rect 47944 32672 48264 33696
rect 47944 32608 47952 32672
rect 48016 32608 48032 32672
rect 48096 32608 48112 32672
rect 48176 32608 48192 32672
rect 48256 32608 48264 32672
rect 47944 31584 48264 32608
rect 47944 31520 47952 31584
rect 48016 31520 48032 31584
rect 48096 31520 48112 31584
rect 48176 31520 48192 31584
rect 48256 31520 48264 31584
rect 47944 30496 48264 31520
rect 47944 30432 47952 30496
rect 48016 30432 48032 30496
rect 48096 30432 48112 30496
rect 48176 30432 48192 30496
rect 48256 30432 48264 30496
rect 47944 29408 48264 30432
rect 47944 29344 47952 29408
rect 48016 29344 48032 29408
rect 48096 29344 48112 29408
rect 48176 29344 48192 29408
rect 48256 29344 48264 29408
rect 47944 28320 48264 29344
rect 47944 28256 47952 28320
rect 48016 28256 48032 28320
rect 48096 28256 48112 28320
rect 48176 28256 48192 28320
rect 48256 28256 48264 28320
rect 47944 27232 48264 28256
rect 47944 27168 47952 27232
rect 48016 27168 48032 27232
rect 48096 27168 48112 27232
rect 48176 27168 48192 27232
rect 48256 27168 48264 27232
rect 47944 26144 48264 27168
rect 47944 26080 47952 26144
rect 48016 26080 48032 26144
rect 48096 26080 48112 26144
rect 48176 26080 48192 26144
rect 48256 26080 48264 26144
rect 47944 25056 48264 26080
rect 47944 24992 47952 25056
rect 48016 24992 48032 25056
rect 48096 24992 48112 25056
rect 48176 24992 48192 25056
rect 48256 24992 48264 25056
rect 47944 23968 48264 24992
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_2  _096_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20608 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _097_
timestamp 1676037725
transform 1 0 18584 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _098_
timestamp 1676037725
transform 1 0 10856 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _099_
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _100_
timestamp 1676037725
transform 1 0 5336 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _101_
timestamp 1676037725
transform 1 0 6532 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1676037725
transform 1 0 4508 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp 1676037725
transform 1 0 6532 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _104_
timestamp 1676037725
transform 1 0 10948 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1676037725
transform 1 0 10856 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _106_
timestamp 1676037725
transform 1 0 7728 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1676037725
transform 1 0 9660 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1676037725
transform 1 0 6624 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1676037725
transform 1 0 6348 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _110_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 4600 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1676037725
transform 1 0 4140 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1676037725
transform 1 0 9016 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1676037725
transform 1 0 9200 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1676037725
transform 1 0 13432 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform 1 0 12604 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1676037725
transform 1 0 4784 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1676037725
transform 1 0 4600 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1676037725
transform 1 0 4508 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 4324 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 3588 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform 1 0 3956 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform 1 0 4324 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1676037725
transform 1 0 3956 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1676037725
transform 1 0 4968 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1676037725
transform 1 0 2392 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1676037725
transform 1 0 4692 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _128_
timestamp 1676037725
transform 1 0 4048 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform 1 0 3496 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1676037725
transform 1 0 7728 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1676037725
transform 1 0 8372 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1676037725
transform 1 0 8280 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1676037725
transform 1 0 9200 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1676037725
transform 1 0 9016 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1676037725
transform 1 0 7636 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _136_
timestamp 1676037725
transform 1 0 8372 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1676037725
transform 1 0 9660 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1676037725
transform 1 0 10304 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1676037725
transform 1 0 10856 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1676037725
transform 1 0 11684 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 11500 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 11868 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp 1676037725
transform 1 0 12144 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 1676037725
transform 1 0 12788 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _145_
timestamp 1676037725
transform 1 0 13524 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1676037725
transform 1 0 15548 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 12236 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 13340 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform 1 0 13340 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 1676037725
transform 1 0 17572 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1676037725
transform 1 0 20976 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1676037725
transform 1 0 20148 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1676037725
transform 1 0 19412 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1676037725
transform 1 0 20976 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 13156 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 14904 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 16836 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 19412 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1676037725
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1676037725
transform 1 0 20792 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform 1 0 25024 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 24932 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 25208 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 24564 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 18032 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 14536 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 18032 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 20056 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 25208 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 22540 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 17572 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 26220 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 18676 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 25760 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 24288 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 26680 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 22816 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 23736 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 27968 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1676037725
transform 1 0 12420 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1676037725
transform 1 0 23736 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1676037725
transform 1 0 20424 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1676037725
transform 1 0 28428 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1676037725
transform 1 0 22172 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1676037725
transform 1 0 18952 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1676037725
transform 1 0 25484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1676037725
transform 1 0 19780 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 16836 0 1 40256
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9660 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 9660 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 9108 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6348 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 6624 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8004 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9016 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 10856 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 11776 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9108 0 1 35904
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 8464 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 6716 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9200 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 5244 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 7544 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 10396 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 11408 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 8004 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 9200 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 9844 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 9936 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__190 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 11684 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 9292 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 10212 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16008 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 5060 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 5244 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 5244 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 9200 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10488 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 5428 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 6624 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 7820 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__191
timestamp 1676037725
transform 1 0 6992 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 7636 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 7452 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 7820 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 9384 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14260 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 5244 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 5428 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 6624 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 7544 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 12604 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 6808 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 7820 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 11132 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 16836 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__192
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 10028 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 12880 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15640 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 6348 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 5244 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 6624 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 7820 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 10212 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 7268 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 7820 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 8832 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__193
timestamp 1676037725
transform 1 0 16836 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 15088 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 5152 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 9200 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12972 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 31004 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21988 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20792 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10396 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 28888 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 25208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 24564 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 19136 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 27232 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 24288 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 25852 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 18584 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24656 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 24932 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 23552 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 30084 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 17112 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32292 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 19504 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9568 0 1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 12144 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 8004 0 -1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 11684 0 -1 42432
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 11868 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 9476 0 1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 15364 0 -1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 16928 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 17388 0 -1 45696
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 20056 0 -1 45696
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 18308 0 -1 50048
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 21988 0 -1 50048
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 20056 0 -1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 21988 0 -1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 17572 0 -1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 21988 0 -1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2116 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1676037725
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75
timestamp 1676037725
transform 1 0 8004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103
timestamp 1676037725
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1676037725
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1676037725
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149
timestamp 1676037725
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1676037725
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1676037725
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_215
timestamp 1676037725
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1676037725
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1676037725
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp 1676037725
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1676037725
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1676037725
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1676037725
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1676037725
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1676037725
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1676037725
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1676037725
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_383
timestamp 1676037725
transform 1 0 36340 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1676037725
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_405
timestamp 1676037725
transform 1 0 38364 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1676037725
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1676037725
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1676037725
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1676037725
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1676037725
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_485
timestamp 1676037725
transform 1 0 45724 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_497
timestamp 1676037725
transform 1 0 46828 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_503
timestamp 1676037725
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_517
timestamp 1676037725
transform 1 0 48668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1676037725
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1676037725
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1676037725
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1676037725
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1676037725
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1676037725
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1676037725
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1676037725
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1676037725
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1676037725
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1676037725
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1676037725
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1676037725
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1676037725
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1676037725
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1676037725
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1676037725
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1676037725
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_293
timestamp 1676037725
transform 1 0 28060 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1676037725
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1676037725
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1676037725
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1676037725
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1676037725
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1676037725
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1676037725
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1676037725
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1676037725
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1676037725
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1676037725
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1676037725
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1676037725
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_485
timestamp 1676037725
transform 1 0 45724 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_493
timestamp 1676037725
transform 1 0 46460 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_499
timestamp 1676037725
transform 1 0 47012 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1676037725
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_517
timestamp 1676037725
transform 1 0 48668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1676037725
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1676037725
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1676037725
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1676037725
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1676037725
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1676037725
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1676037725
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1676037725
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1676037725
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1676037725
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1676037725
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1676037725
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1676037725
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1676037725
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1676037725
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1676037725
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1676037725
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1676037725
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1676037725
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1676037725
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1676037725
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1676037725
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1676037725
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1676037725
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1676037725
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1676037725
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1676037725
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_517
timestamp 1676037725
transform 1 0 48668 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1676037725
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1676037725
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1676037725
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1676037725
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_9
timestamp 1676037725
transform 1 0 1932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_21
timestamp 1676037725
transform 1 0 3036 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_33
timestamp 1676037725
transform 1 0 4140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_45
timestamp 1676037725
transform 1 0 5244 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1676037725
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1676037725
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1676037725
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1676037725
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1676037725
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1676037725
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1676037725
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_517
timestamp 1676037725
transform 1 0 48668 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1676037725
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_9
timestamp 1676037725
transform 1 0 1932 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_21
timestamp 1676037725
transform 1 0 3036 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_203
timestamp 1676037725
transform 1 0 19780 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_215
timestamp 1676037725
transform 1 0 20884 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_227
timestamp 1676037725
transform 1 0 21988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_239
timestamp 1676037725
transform 1 0 23092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1676037725
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1676037725
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1676037725
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_175
timestamp 1676037725
transform 1 0 17204 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_187
timestamp 1676037725
transform 1 0 18308 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_199
timestamp 1676037725
transform 1 0 19412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_211
timestamp 1676037725
transform 1 0 20516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_257
timestamp 1676037725
transform 1 0 24748 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_264
timestamp 1676037725
transform 1 0 25392 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1676037725
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1676037725
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1676037725
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1676037725
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1676037725
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_9
timestamp 1676037725
transform 1 0 1932 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_21
timestamp 1676037725
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_149
timestamp 1676037725
transform 1 0 14812 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_154
timestamp 1676037725
transform 1 0 15272 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_166
timestamp 1676037725
transform 1 0 16376 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_178
timestamp 1676037725
transform 1 0 17480 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_190
timestamp 1676037725
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1676037725
transform 1 0 20700 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_218
timestamp 1676037725
transform 1 0 21160 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_230
timestamp 1676037725
transform 1 0 22264 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_237
timestamp 1676037725
transform 1 0 22908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp 1676037725
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1676037725
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1676037725
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1676037725
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_9
timestamp 1676037725
transform 1 0 1932 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_21
timestamp 1676037725
transform 1 0 3036 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_33
timestamp 1676037725
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1676037725
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1676037725
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1676037725
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1676037725
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1676037725
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1676037725
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1676037725
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1676037725
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1676037725
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1676037725
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1676037725
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1676037725
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1676037725
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_517
timestamp 1676037725
transform 1 0 48668 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1676037725
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_129
timestamp 1676037725
transform 1 0 12972 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1676037725
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1676037725
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1676037725
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1676037725
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1676037725
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1676037725
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1676037725
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1676037725
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1676037725
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1676037725
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1676037725
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_8
timestamp 1676037725
transform 1 0 1840 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_20
timestamp 1676037725
transform 1 0 2944 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_32
timestamp 1676037725
transform 1 0 4048 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_44
timestamp 1676037725
transform 1 0 5152 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1676037725
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1676037725
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1676037725
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1676037725
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1676037725
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1676037725
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1676037725
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1676037725
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1676037725
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1676037725
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1676037725
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1676037725
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1676037725
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1676037725
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1676037725
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1676037725
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1676037725
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1676037725
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1676037725
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1676037725
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1676037725
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_517
timestamp 1676037725
transform 1 0 48668 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1676037725
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_8
timestamp 1676037725
transform 1 0 1840 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1676037725
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_185
timestamp 1676037725
transform 1 0 18124 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_190
timestamp 1676037725
transform 1 0 18584 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1676037725
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1676037725
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1676037725
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1676037725
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1676037725
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1676037725
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1676037725
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1676037725
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1676037725
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1676037725
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1676037725
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1676037725
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1676037725
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1676037725
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1676037725
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1676037725
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1676037725
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1676037725
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1676037725
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1676037725
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1676037725
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1676037725
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1676037725
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1676037725
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1676037725
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1676037725
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1676037725
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1676037725
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1676037725
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1676037725
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1676037725
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1676037725
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1676037725
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1676037725
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1676037725
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1676037725
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_517
timestamp 1676037725
transform 1 0 48668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1676037725
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_9
timestamp 1676037725
transform 1 0 1932 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_21
timestamp 1676037725
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1676037725
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1676037725
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1676037725
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1676037725
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1676037725
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1676037725
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1676037725
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1676037725
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1676037725
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1676037725
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1676037725
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1676037725
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1676037725
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1676037725
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1676037725
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1676037725
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1676037725
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1676037725
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1676037725
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1676037725
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1676037725
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1676037725
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1676037725
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1676037725
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_9
timestamp 1676037725
transform 1 0 1932 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_21
timestamp 1676037725
transform 1 0 3036 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_33
timestamp 1676037725
transform 1 0 4140 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_45
timestamp 1676037725
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1676037725
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1676037725
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1676037725
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1676037725
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1676037725
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1676037725
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1676037725
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1676037725
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1676037725
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1676037725
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1676037725
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1676037725
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1676037725
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1676037725
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1676037725
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1676037725
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1676037725
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1676037725
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1676037725
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1676037725
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1676037725
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1676037725
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1676037725
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1676037725
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1676037725
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1676037725
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1676037725
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1676037725
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1676037725
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_517
timestamp 1676037725
transform 1 0 48668 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1676037725
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1676037725
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1676037725
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1676037725
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1676037725
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1676037725
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1676037725
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1676037725
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1676037725
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_223
timestamp 1676037725
transform 1 0 21620 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1676037725
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1676037725
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1676037725
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1676037725
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1676037725
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1676037725
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1676037725
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1676037725
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1676037725
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1676037725
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1676037725
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1676037725
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1676037725
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1676037725
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1676037725
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1676037725
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1676037725
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1676037725
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1676037725
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1676037725
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1676037725
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1676037725
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1676037725
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1676037725
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1676037725
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1676037725
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1676037725
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_9
timestamp 1676037725
transform 1 0 1932 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_21
timestamp 1676037725
transform 1 0 3036 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_33
timestamp 1676037725
transform 1 0 4140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_45
timestamp 1676037725
transform 1 0 5244 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp 1676037725
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1676037725
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1676037725
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1676037725
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1676037725
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1676037725
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1676037725
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1676037725
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1676037725
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1676037725
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1676037725
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1676037725
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1676037725
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1676037725
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1676037725
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1676037725
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1676037725
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1676037725
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1676037725
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1676037725
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1676037725
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1676037725
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1676037725
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1676037725
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1676037725
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1676037725
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1676037725
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1676037725
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_517
timestamp 1676037725
transform 1 0 48668 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1676037725
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_9
timestamp 1676037725
transform 1 0 1932 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_21
timestamp 1676037725
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1676037725
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1676037725
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1676037725
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1676037725
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1676037725
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1676037725
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1676037725
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1676037725
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1676037725
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1676037725
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1676037725
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1676037725
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1676037725
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1676037725
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1676037725
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1676037725
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1676037725
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1676037725
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1676037725
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1676037725
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1676037725
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1676037725
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1676037725
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1676037725
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1676037725
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1676037725
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_193
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_204
timestamp 1676037725
transform 1 0 19872 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_212
timestamp 1676037725
transform 1 0 20608 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1676037725
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1676037725
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1676037725
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1676037725
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1676037725
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1676037725
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1676037725
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1676037725
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1676037725
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1676037725
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1676037725
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1676037725
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1676037725
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1676037725
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1676037725
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1676037725
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1676037725
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1676037725
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1676037725
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1676037725
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1676037725
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1676037725
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1676037725
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1676037725
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1676037725
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_517
timestamp 1676037725
transform 1 0 48668 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1676037725
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_8
timestamp 1676037725
transform 1 0 1840 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1676037725
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1676037725
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1676037725
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1676037725
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1676037725
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1676037725
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1676037725
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1676037725
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_261
timestamp 1676037725
transform 1 0 25116 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_267
timestamp 1676037725
transform 1 0 25668 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_279
timestamp 1676037725
transform 1 0 26772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_291
timestamp 1676037725
transform 1 0 27876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1676037725
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1676037725
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1676037725
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1676037725
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1676037725
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1676037725
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1676037725
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1676037725
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1676037725
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1676037725
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1676037725
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1676037725
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1676037725
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1676037725
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1676037725
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1676037725
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1676037725
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1676037725
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_8
timestamp 1676037725
transform 1 0 1840 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_20
timestamp 1676037725
transform 1 0 2944 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_32
timestamp 1676037725
transform 1 0 4048 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_44
timestamp 1676037725
transform 1 0 5152 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1676037725
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1676037725
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1676037725
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1676037725
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1676037725
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1676037725
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1676037725
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1676037725
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1676037725
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_286
timestamp 1676037725
transform 1 0 27416 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_298
timestamp 1676037725
transform 1 0 28520 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_310
timestamp 1676037725
transform 1 0 29624 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_322
timestamp 1676037725
transform 1 0 30728 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1676037725
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1676037725
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1676037725
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1676037725
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1676037725
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1676037725
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1676037725
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1676037725
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1676037725
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1676037725
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1676037725
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1676037725
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1676037725
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1676037725
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1676037725
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1676037725
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_517
timestamp 1676037725
transform 1 0 48668 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1676037725
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1676037725
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1676037725
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1676037725
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1676037725
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1676037725
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1676037725
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1676037725
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_261
timestamp 1676037725
transform 1 0 25116 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1676037725
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1676037725
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1676037725
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1676037725
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1676037725
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1676037725
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1676037725
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1676037725
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1676037725
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1676037725
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1676037725
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1676037725
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1676037725
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1676037725
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1676037725
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1676037725
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1676037725
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1676037725
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1676037725
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1676037725
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1676037725
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1676037725
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1676037725
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1676037725
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1676037725
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1676037725
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1676037725
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1676037725
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1676037725
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_249
timestamp 1676037725
transform 1 0 24012 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_255
timestamp 1676037725
transform 1 0 24564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_267
timestamp 1676037725
transform 1 0 25668 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1676037725
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1676037725
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1676037725
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1676037725
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1676037725
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1676037725
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1676037725
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1676037725
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1676037725
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1676037725
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1676037725
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1676037725
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1676037725
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1676037725
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1676037725
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1676037725
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1676037725
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1676037725
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1676037725
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1676037725
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_517
timestamp 1676037725
transform 1 0 48668 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1676037725
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_9
timestamp 1676037725
transform 1 0 1932 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_21
timestamp 1676037725
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1676037725
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1676037725
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1676037725
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1676037725
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1676037725
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1676037725
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1676037725
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1676037725
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1676037725
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_265
timestamp 1676037725
transform 1 0 25484 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_276
timestamp 1676037725
transform 1 0 26496 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_288
timestamp 1676037725
transform 1 0 27600 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_300
timestamp 1676037725
transform 1 0 28704 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1676037725
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1676037725
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1676037725
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1676037725
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1676037725
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1676037725
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1676037725
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1676037725
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1676037725
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1676037725
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1676037725
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1676037725
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1676037725
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1676037725
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1676037725
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1676037725
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1676037725
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1676037725
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1676037725
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1676037725
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1676037725
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1676037725
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1676037725
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1676037725
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1676037725
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1676037725
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1676037725
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1676037725
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1676037725
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1676037725
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1676037725
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1676037725
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1676037725
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1676037725
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1676037725
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1676037725
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1676037725
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1676037725
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1676037725
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1676037725
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1676037725
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1676037725
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1676037725
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1676037725
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1676037725
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1676037725
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1676037725
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1676037725
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1676037725
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1676037725
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1676037725
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1676037725
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1676037725
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_517
timestamp 1676037725
transform 1 0 48668 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1676037725
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_9
timestamp 1676037725
transform 1 0 1932 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_21
timestamp 1676037725
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1676037725
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1676037725
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1676037725
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1676037725
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1676037725
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1676037725
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1676037725
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1676037725
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1676037725
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1676037725
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_233
timestamp 1676037725
transform 1 0 22540 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_241
timestamp 1676037725
transform 1 0 23276 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_247
timestamp 1676037725
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1676037725
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1676037725
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1676037725
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1676037725
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1676037725
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1676037725
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_321
timestamp 1676037725
transform 1 0 30636 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_346
timestamp 1676037725
transform 1 0 32936 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_358
timestamp 1676037725
transform 1 0 34040 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1676037725
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1676037725
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_401
timestamp 1676037725
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1676037725
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1676037725
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1676037725
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1676037725
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1676037725
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1676037725
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1676037725
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1676037725
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1676037725
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1676037725
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1676037725
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_9
timestamp 1676037725
transform 1 0 1932 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_21
timestamp 1676037725
transform 1 0 3036 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_33
timestamp 1676037725
transform 1 0 4140 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_45
timestamp 1676037725
transform 1 0 5244 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1676037725
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1676037725
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1676037725
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_173
timestamp 1676037725
transform 1 0 17020 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_182
timestamp 1676037725
transform 1 0 17848 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_194
timestamp 1676037725
transform 1 0 18952 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_206
timestamp 1676037725
transform 1 0 20056 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1676037725
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1676037725
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_249
timestamp 1676037725
transform 1 0 24012 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_255
timestamp 1676037725
transform 1 0 24564 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1676037725
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_293
timestamp 1676037725
transform 1 0 28060 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_301
timestamp 1676037725
transform 1 0 28796 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_323
timestamp 1676037725
transform 1 0 30820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1676037725
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1676037725
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1676037725
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1676037725
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1676037725
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1676037725
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1676037725
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1676037725
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1676037725
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1676037725
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1676037725
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1676037725
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1676037725
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1676037725
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1676037725
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_517
timestamp 1676037725
transform 1 0 48668 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1676037725
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1676037725
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1676037725
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1676037725
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1676037725
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1676037725
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1676037725
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1676037725
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_280
timestamp 1676037725
transform 1 0 26864 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_305
timestamp 1676037725
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1676037725
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1676037725
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1676037725
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1676037725
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1676037725
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1676037725
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1676037725
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1676037725
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1676037725
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1676037725
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1676037725
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1676037725
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1676037725
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1676037725
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1676037725
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1676037725
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1676037725
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1676037725
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1676037725
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_8
timestamp 1676037725
transform 1 0 1840 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_20
timestamp 1676037725
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_32
timestamp 1676037725
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_44
timestamp 1676037725
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1676037725
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1676037725
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1676037725
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1676037725
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1676037725
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1676037725
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1676037725
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1676037725
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1676037725
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1676037725
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1676037725
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1676037725
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1676037725
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1676037725
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1676037725
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1676037725
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1676037725
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1676037725
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_405
timestamp 1676037725
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_417
timestamp 1676037725
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_429
timestamp 1676037725
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1676037725
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1676037725
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1676037725
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1676037725
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1676037725
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1676037725
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1676037725
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_517
timestamp 1676037725
transform 1 0 48668 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1676037725
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_8
timestamp 1676037725
transform 1 0 1840 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_20
timestamp 1676037725
transform 1 0 2944 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1676037725
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1676037725
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1676037725
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1676037725
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1676037725
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1676037725
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1676037725
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1676037725
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1676037725
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1676037725
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1676037725
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1676037725
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1676037725
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1676037725
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1676037725
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1676037725
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1676037725
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_401
timestamp 1676037725
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1676037725
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1676037725
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1676037725
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1676037725
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_457
timestamp 1676037725
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1676037725
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1676037725
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1676037725
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1676037725
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1676037725
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1676037725
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1676037725
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1676037725
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1676037725
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1676037725
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1676037725
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1676037725
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1676037725
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1676037725
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1676037725
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1676037725
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1676037725
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1676037725
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1676037725
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1676037725
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1676037725
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1676037725
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1676037725
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1676037725
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1676037725
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1676037725
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1676037725
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1676037725
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_417
timestamp 1676037725
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_429
timestamp 1676037725
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1676037725
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1676037725
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1676037725
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1676037725
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1676037725
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1676037725
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1676037725
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_517
timestamp 1676037725
transform 1 0 48668 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1676037725
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_9
timestamp 1676037725
transform 1 0 1932 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_21
timestamp 1676037725
transform 1 0 3036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1676037725
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1676037725
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1676037725
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1676037725
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1676037725
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1676037725
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1676037725
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1676037725
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1676037725
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1676037725
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1676037725
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1676037725
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1676037725
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1676037725
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1676037725
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1676037725
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1676037725
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1676037725
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1676037725
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1676037725
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1676037725
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1676037725
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1676037725
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1676037725
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1676037725
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1676037725
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_401
timestamp 1676037725
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_413
timestamp 1676037725
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_419
timestamp 1676037725
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1676037725
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1676037725
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1676037725
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1676037725
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1676037725
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1676037725
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1676037725
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1676037725
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1676037725
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1676037725
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1676037725
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1676037725
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1676037725
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1676037725
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1676037725
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1676037725
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_161
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1676037725
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1676037725
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1676037725
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1676037725
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1676037725
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1676037725
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1676037725
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1676037725
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1676037725
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1676037725
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1676037725
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_305
timestamp 1676037725
transform 1 0 29164 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_313
timestamp 1676037725
transform 1 0 29900 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_322
timestamp 1676037725
transform 1 0 30728 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1676037725
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1676037725
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1676037725
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1676037725
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1676037725
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1676037725
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1676037725
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1676037725
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1676037725
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1676037725
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1676037725
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1676037725
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1676037725
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1676037725
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1676037725
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1676037725
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_517
timestamp 1676037725
transform 1 0 48668 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1676037725
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1676037725
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1676037725
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1676037725
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1676037725
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1676037725
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1676037725
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1676037725
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1676037725
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1676037725
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1676037725
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_146
timestamp 1676037725
transform 1 0 14536 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_161
timestamp 1676037725
transform 1 0 15916 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_173
timestamp 1676037725
transform 1 0 17020 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_185
timestamp 1676037725
transform 1 0 18124 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_193
timestamp 1676037725
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1676037725
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1676037725
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1676037725
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1676037725
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1676037725
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1676037725
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1676037725
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1676037725
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1676037725
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1676037725
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1676037725
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1676037725
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1676037725
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1676037725
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1676037725
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1676037725
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1676037725
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1676037725
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1676037725
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1676037725
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1676037725
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1676037725
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1676037725
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1676037725
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1676037725
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1676037725
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1676037725
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_525
timestamp 1676037725
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1676037725
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1676037725
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1676037725
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1676037725
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1676037725
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1676037725
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1676037725
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1676037725
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1676037725
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1676037725
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1676037725
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1676037725
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1676037725
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1676037725
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1676037725
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1676037725
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1676037725
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1676037725
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1676037725
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1676037725
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1676037725
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1676037725
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1676037725
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1676037725
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1676037725
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1676037725
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1676037725
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1676037725
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1676037725
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_405
timestamp 1676037725
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_417
timestamp 1676037725
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_429
timestamp 1676037725
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1676037725
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1676037725
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1676037725
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1676037725
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1676037725
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1676037725
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1676037725
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_517
timestamp 1676037725
transform 1 0 48668 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1676037725
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1676037725
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1676037725
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1676037725
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1676037725
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1676037725
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1676037725
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1676037725
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1676037725
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1676037725
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1676037725
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1676037725
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1676037725
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1676037725
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1676037725
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_221
timestamp 1676037725
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_233
timestamp 1676037725
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1676037725
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1676037725
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1676037725
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1676037725
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1676037725
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1676037725
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1676037725
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1676037725
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1676037725
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1676037725
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1676037725
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1676037725
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1676037725
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1676037725
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_401
timestamp 1676037725
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_413
timestamp 1676037725
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1676037725
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1676037725
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1676037725
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1676037725
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1676037725
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1676037725
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1676037725
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1676037725
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1676037725
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1676037725
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1676037725
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1676037725
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1676037725
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1676037725
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1676037725
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1676037725
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1676037725
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1676037725
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1676037725
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1676037725
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1676037725
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1676037725
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_237
timestamp 1676037725
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1676037725
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1676037725
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1676037725
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1676037725
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1676037725
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1676037725
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1676037725
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1676037725
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1676037725
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1676037725
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1676037725
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1676037725
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1676037725
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1676037725
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_405
timestamp 1676037725
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_417
timestamp 1676037725
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_429
timestamp 1676037725
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1676037725
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1676037725
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1676037725
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1676037725
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1676037725
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1676037725
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1676037725
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1676037725
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_517
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1676037725
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1676037725
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1676037725
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1676037725
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1676037725
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1676037725
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1676037725
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1676037725
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_109
timestamp 1676037725
transform 1 0 11132 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_126
timestamp 1676037725
transform 1 0 12696 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1676037725
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1676037725
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1676037725
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1676037725
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1676037725
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1676037725
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1676037725
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1676037725
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1676037725
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_277
timestamp 1676037725
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_289
timestamp 1676037725
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1676037725
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1676037725
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1676037725
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1676037725
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1676037725
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1676037725
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1676037725
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1676037725
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1676037725
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_401
timestamp 1676037725
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1676037725
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1676037725
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_433
timestamp 1676037725
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_445
timestamp 1676037725
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_457
timestamp 1676037725
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1676037725
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1676037725
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1676037725
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1676037725
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1676037725
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1676037725
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1676037725
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1676037725
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1676037725
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1676037725
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1676037725
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_128
timestamp 1676037725
transform 1 0 12880 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_135
timestamp 1676037725
transform 1 0 13524 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_147
timestamp 1676037725
transform 1 0 14628 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_159
timestamp 1676037725
transform 1 0 15732 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1676037725
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1676037725
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1676037725
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1676037725
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1676037725
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1676037725
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1676037725
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1676037725
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1676037725
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1676037725
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1676037725
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1676037725
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1676037725
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1676037725
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1676037725
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1676037725
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1676037725
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1676037725
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1676037725
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_405
timestamp 1676037725
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_417
timestamp 1676037725
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1676037725
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1676037725
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1676037725
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1676037725
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1676037725
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1676037725
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1676037725
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1676037725
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_517
timestamp 1676037725
transform 1 0 48668 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_525
timestamp 1676037725
transform 1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1676037725
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1676037725
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_110
timestamp 1676037725
transform 1 0 11224 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_118
timestamp 1676037725
transform 1 0 11960 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_124
timestamp 1676037725
transform 1 0 12512 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1676037725
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1676037725
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1676037725
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1676037725
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1676037725
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1676037725
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1676037725
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1676037725
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1676037725
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1676037725
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1676037725
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1676037725
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_277
timestamp 1676037725
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_289
timestamp 1676037725
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1676037725
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1676037725
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1676037725
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1676037725
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1676037725
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1676037725
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1676037725
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1676037725
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1676037725
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1676037725
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1676037725
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1676037725
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_433
timestamp 1676037725
transform 1 0 40940 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_445
timestamp 1676037725
transform 1 0 42044 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_457
timestamp 1676037725
transform 1 0 43148 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_469
timestamp 1676037725
transform 1 0 44252 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1676037725
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1676037725
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1676037725
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1676037725
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_525
timestamp 1676037725
transform 1 0 49404 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_9
timestamp 1676037725
transform 1 0 1932 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_21
timestamp 1676037725
transform 1 0 3036 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_33
timestamp 1676037725
transform 1 0 4140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_45
timestamp 1676037725
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1676037725
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1676037725
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1676037725
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1676037725
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1676037725
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1676037725
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1676037725
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1676037725
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1676037725
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1676037725
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1676037725
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1676037725
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1676037725
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1676037725
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1676037725
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1676037725
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1676037725
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1676037725
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1676037725
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1676037725
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1676037725
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1676037725
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_362
timestamp 1676037725
transform 1 0 34408 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_374
timestamp 1676037725
transform 1 0 35512 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_386
timestamp 1676037725
transform 1 0 36616 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1676037725
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_405
timestamp 1676037725
transform 1 0 38364 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_417
timestamp 1676037725
transform 1 0 39468 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_429
timestamp 1676037725
transform 1 0 40572 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_441
timestamp 1676037725
transform 1 0 41676 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1676037725
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1676037725
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1676037725
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1676037725
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1676037725
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1676037725
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1676037725
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1676037725
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_517
timestamp 1676037725
transform 1 0 48668 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_525
timestamp 1676037725
transform 1 0 49404 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1676037725
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1676037725
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1676037725
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1676037725
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1676037725
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_108
timestamp 1676037725
transform 1 0 11040 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_115
timestamp 1676037725
transform 1 0 11684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_127
timestamp 1676037725
transform 1 0 12788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1676037725
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1676037725
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1676037725
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1676037725
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1676037725
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1676037725
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1676037725
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1676037725
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1676037725
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1676037725
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1676037725
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1676037725
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1676037725
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1676037725
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1676037725
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1676037725
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1676037725
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1676037725
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1676037725
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1676037725
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1676037725
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1676037725
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1676037725
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1676037725
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1676037725
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1676037725
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1676037725
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1676037725
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1676037725
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1676037725
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1676037725
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1676037725
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1676037725
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1676037725
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1676037725
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1676037725
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1676037725
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_525
timestamp 1676037725
transform 1 0 49404 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1676037725
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1676037725
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1676037725
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1676037725
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1676037725
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1676037725
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1676037725
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1676037725
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1676037725
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1676037725
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1676037725
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1676037725
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1676037725
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1676037725
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1676037725
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1676037725
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1676037725
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1676037725
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1676037725
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1676037725
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1676037725
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1676037725
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1676037725
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1676037725
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1676037725
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1676037725
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1676037725
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1676037725
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1676037725
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_405
timestamp 1676037725
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_417
timestamp 1676037725
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_429
timestamp 1676037725
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1676037725
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1676037725
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1676037725
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1676037725
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1676037725
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1676037725
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1676037725
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1676037725
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1676037725
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_517
timestamp 1676037725
transform 1 0 48668 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_525
timestamp 1676037725
transform 1 0 49404 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1676037725
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1676037725
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1676037725
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1676037725
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1676037725
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1676037725
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1676037725
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1676037725
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1676037725
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1676037725
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1676037725
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1676037725
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1676037725
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1676037725
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1676037725
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1676037725
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1676037725
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1676037725
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1676037725
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1676037725
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1676037725
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1676037725
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1676037725
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1676037725
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1676037725
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1676037725
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_401
timestamp 1676037725
transform 1 0 37996 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_413
timestamp 1676037725
transform 1 0 39100 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1676037725
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_421
timestamp 1676037725
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_433
timestamp 1676037725
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_445
timestamp 1676037725
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_457
timestamp 1676037725
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1676037725
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1676037725
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1676037725
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1676037725
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1676037725
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1676037725
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_525
timestamp 1676037725
transform 1 0 49404 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_9
timestamp 1676037725
transform 1 0 1932 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_21
timestamp 1676037725
transform 1 0 3036 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_33
timestamp 1676037725
transform 1 0 4140 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_45
timestamp 1676037725
transform 1 0 5244 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1676037725
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1676037725
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1676037725
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1676037725
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1676037725
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_124
timestamp 1676037725
transform 1 0 12512 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_136
timestamp 1676037725
transform 1 0 13616 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_148
timestamp 1676037725
transform 1 0 14720 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_160
timestamp 1676037725
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1676037725
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1676037725
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1676037725
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1676037725
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1676037725
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1676037725
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1676037725
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1676037725
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1676037725
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1676037725
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1676037725
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1676037725
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1676037725
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1676037725
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1676037725
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1676037725
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1676037725
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1676037725
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1676037725
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1676037725
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1676037725
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_405
timestamp 1676037725
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_417
timestamp 1676037725
transform 1 0 39468 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_429
timestamp 1676037725
transform 1 0 40572 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_441
timestamp 1676037725
transform 1 0 41676 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1676037725
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1676037725
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1676037725
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1676037725
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1676037725
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1676037725
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1676037725
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1676037725
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_517
timestamp 1676037725
transform 1 0 48668 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_525
timestamp 1676037725
transform 1 0 49404 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1676037725
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1676037725
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1676037725
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_109
timestamp 1676037725
transform 1 0 11132 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_124
timestamp 1676037725
transform 1 0 12512 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_128
timestamp 1676037725
transform 1 0 12880 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_132
timestamp 1676037725
transform 1 0 13248 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1676037725
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1676037725
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1676037725
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1676037725
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1676037725
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1676037725
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1676037725
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1676037725
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1676037725
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1676037725
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1676037725
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1676037725
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1676037725
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1676037725
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1676037725
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1676037725
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1676037725
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1676037725
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1676037725
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1676037725
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_401
timestamp 1676037725
transform 1 0 37996 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_413
timestamp 1676037725
transform 1 0 39100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_419
timestamp 1676037725
transform 1 0 39652 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1676037725
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1676037725
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1676037725
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1676037725
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1676037725
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1676037725
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1676037725
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1676037725
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1676037725
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1676037725
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_525
timestamp 1676037725
transform 1 0 49404 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_21
timestamp 1676037725
transform 1 0 3036 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_33
timestamp 1676037725
transform 1 0 4140 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_45
timestamp 1676037725
transform 1 0 5244 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_53
timestamp 1676037725
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_81
timestamp 1676037725
transform 1 0 8556 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_89
timestamp 1676037725
transform 1 0 9292 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_99
timestamp 1676037725
transform 1 0 10212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1676037725
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_134
timestamp 1676037725
transform 1 0 13432 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_146
timestamp 1676037725
transform 1 0 14536 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_158
timestamp 1676037725
transform 1 0 15640 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1676037725
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1676037725
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1676037725
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1676037725
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1676037725
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1676037725
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1676037725
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1676037725
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1676037725
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1676037725
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1676037725
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1676037725
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1676037725
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1676037725
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1676037725
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1676037725
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1676037725
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1676037725
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1676037725
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1676037725
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1676037725
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1676037725
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1676037725
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1676037725
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1676037725
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1676037725
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1676037725
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1676037725
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1676037725
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1676037725
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1676037725
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1676037725
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1676037725
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1676037725
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_517
timestamp 1676037725
transform 1 0 48668 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_525
timestamp 1676037725
transform 1 0 49404 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_21
timestamp 1676037725
transform 1 0 3036 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1676037725
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_93
timestamp 1676037725
transform 1 0 9660 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_104
timestamp 1676037725
transform 1 0 10672 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_108
timestamp 1676037725
transform 1 0 11040 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_118
timestamp 1676037725
transform 1 0 11960 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_131
timestamp 1676037725
transform 1 0 13156 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1676037725
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1676037725
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1676037725
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1676037725
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1676037725
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1676037725
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1676037725
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1676037725
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1676037725
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1676037725
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1676037725
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1676037725
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1676037725
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1676037725
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1676037725
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1676037725
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1676037725
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1676037725
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1676037725
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1676037725
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1676037725
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1676037725
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1676037725
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1676037725
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_401
timestamp 1676037725
transform 1 0 37996 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1676037725
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1676037725
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1676037725
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1676037725
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1676037725
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1676037725
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1676037725
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1676037725
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1676037725
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1676037725
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1676037725
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1676037725
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_525
timestamp 1676037725
transform 1 0 49404 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_89
timestamp 1676037725
transform 1 0 9292 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_97
timestamp 1676037725
transform 1 0 10028 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1676037725
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1676037725
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1676037725
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1676037725
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1676037725
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1676037725
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1676037725
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1676037725
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1676037725
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1676037725
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1676037725
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1676037725
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1676037725
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1676037725
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1676037725
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1676037725
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1676037725
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1676037725
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1676037725
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1676037725
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1676037725
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1676037725
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1676037725
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1676037725
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1676037725
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1676037725
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1676037725
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_405
timestamp 1676037725
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_417
timestamp 1676037725
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_429
timestamp 1676037725
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1676037725
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1676037725
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1676037725
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1676037725
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1676037725
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1676037725
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1676037725
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1676037725
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1676037725
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_517
timestamp 1676037725
transform 1 0 48668 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_525
timestamp 1676037725
transform 1 0 49404 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_21
timestamp 1676037725
transform 1 0 3036 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_113
timestamp 1676037725
transform 1 0 11500 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_128
timestamp 1676037725
transform 1 0 12880 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_152
timestamp 1676037725
transform 1 0 15088 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_164
timestamp 1676037725
transform 1 0 16192 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_176
timestamp 1676037725
transform 1 0 17296 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_188
timestamp 1676037725
transform 1 0 18400 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1676037725
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1676037725
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1676037725
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1676037725
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1676037725
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1676037725
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1676037725
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1676037725
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1676037725
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1676037725
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1676037725
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1676037725
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1676037725
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1676037725
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1676037725
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1676037725
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1676037725
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1676037725
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1676037725
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1676037725
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1676037725
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1676037725
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1676037725
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1676037725
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1676037725
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1676037725
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1676037725
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1676037725
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1676037725
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1676037725
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1676037725
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1676037725
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_525
timestamp 1676037725
transform 1 0 49404 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_21
timestamp 1676037725
transform 1 0 3036 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_33
timestamp 1676037725
transform 1 0 4140 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_45
timestamp 1676037725
transform 1 0 5244 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_53
timestamp 1676037725
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_69
timestamp 1676037725
transform 1 0 7452 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_98
timestamp 1676037725
transform 1 0 10120 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1676037725
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_136
timestamp 1676037725
transform 1 0 13616 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_149
timestamp 1676037725
transform 1 0 14812 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_156
timestamp 1676037725
transform 1 0 15456 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1676037725
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1676037725
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1676037725
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1676037725
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1676037725
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1676037725
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1676037725
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1676037725
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1676037725
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1676037725
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1676037725
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1676037725
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1676037725
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1676037725
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1676037725
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1676037725
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1676037725
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1676037725
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1676037725
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1676037725
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1676037725
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1676037725
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1676037725
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_417
timestamp 1676037725
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_429
timestamp 1676037725
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1676037725
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1676037725
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1676037725
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1676037725
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1676037725
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1676037725
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1676037725
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1676037725
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1676037725
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_517
timestamp 1676037725
transform 1 0 48668 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_525
timestamp 1676037725
transform 1 0 49404 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1676037725
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_102
timestamp 1676037725
transform 1 0 10488 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_126
timestamp 1676037725
transform 1 0 12696 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1676037725
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_146
timestamp 1676037725
transform 1 0 14536 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_171
timestamp 1676037725
transform 1 0 16836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_183
timestamp 1676037725
transform 1 0 17940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1676037725
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1676037725
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1676037725
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1676037725
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1676037725
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1676037725
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1676037725
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1676037725
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1676037725
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1676037725
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1676037725
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1676037725
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1676037725
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1676037725
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1676037725
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1676037725
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1676037725
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1676037725
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1676037725
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1676037725
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_401
timestamp 1676037725
transform 1 0 37996 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_413
timestamp 1676037725
transform 1 0 39100 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1676037725
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1676037725
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1676037725
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1676037725
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1676037725
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1676037725
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1676037725
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1676037725
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1676037725
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1676037725
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1676037725
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_525
timestamp 1676037725
transform 1 0 49404 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_21
timestamp 1676037725
transform 1 0 3036 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_33
timestamp 1676037725
transform 1 0 4140 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1676037725
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1676037725
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1676037725
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_138
timestamp 1676037725
transform 1 0 13800 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1676037725
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_177
timestamp 1676037725
transform 1 0 17388 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_200
timestamp 1676037725
transform 1 0 19504 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_212
timestamp 1676037725
transform 1 0 20608 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1676037725
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1676037725
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1676037725
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1676037725
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1676037725
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1676037725
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1676037725
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1676037725
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1676037725
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1676037725
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1676037725
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1676037725
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1676037725
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1676037725
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1676037725
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1676037725
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1676037725
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1676037725
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1676037725
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1676037725
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1676037725
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1676037725
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1676037725
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1676037725
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1676037725
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1676037725
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1676037725
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1676037725
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1676037725
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_517
timestamp 1676037725
transform 1 0 48668 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_525
timestamp 1676037725
transform 1 0 49404 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_21
timestamp 1676037725
transform 1 0 3036 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_59
timestamp 1676037725
transform 1 0 6532 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_80
timestamp 1676037725
transform 1 0 8464 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_107
timestamp 1676037725
transform 1 0 10948 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_115
timestamp 1676037725
transform 1 0 11684 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_138
timestamp 1676037725
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_146
timestamp 1676037725
transform 1 0 14536 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_159
timestamp 1676037725
transform 1 0 15732 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_183
timestamp 1676037725
transform 1 0 17940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1676037725
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1676037725
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1676037725
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1676037725
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1676037725
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1676037725
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1676037725
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1676037725
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1676037725
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1676037725
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1676037725
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1676037725
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1676037725
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1676037725
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1676037725
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1676037725
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1676037725
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1676037725
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1676037725
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1676037725
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_401
timestamp 1676037725
transform 1 0 37996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_413
timestamp 1676037725
transform 1 0 39100 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_419
timestamp 1676037725
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1676037725
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1676037725
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1676037725
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1676037725
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1676037725
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1676037725
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1676037725
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1676037725
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1676037725
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1676037725
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_525
timestamp 1676037725
transform 1 0 49404 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1676037725
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1676037725
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1676037725
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1676037725
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1676037725
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_63
timestamp 1676037725
transform 1 0 6900 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_67
timestamp 1676037725
transform 1 0 7268 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_80
timestamp 1676037725
transform 1 0 8464 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_106
timestamp 1676037725
transform 1 0 10856 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_118
timestamp 1676037725
transform 1 0 11960 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_142
timestamp 1676037725
transform 1 0 14168 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_166
timestamp 1676037725
transform 1 0 16376 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_173
timestamp 1676037725
transform 1 0 17020 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_194
timestamp 1676037725
transform 1 0 18952 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_219
timestamp 1676037725
transform 1 0 21252 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1676037725
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1676037725
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1676037725
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1676037725
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1676037725
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1676037725
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1676037725
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1676037725
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1676037725
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1676037725
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1676037725
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1676037725
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1676037725
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1676037725
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1676037725
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1676037725
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1676037725
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1676037725
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1676037725
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1676037725
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1676037725
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1676037725
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1676037725
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1676037725
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1676037725
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1676037725
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1676037725
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1676037725
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1676037725
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1676037725
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_517
timestamp 1676037725
transform 1 0 48668 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_525
timestamp 1676037725
transform 1 0 49404 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_21
timestamp 1676037725
transform 1 0 3036 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_45
timestamp 1676037725
transform 1 0 5244 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_50
timestamp 1676037725
transform 1 0 5704 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_62
timestamp 1676037725
transform 1 0 6808 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_68
timestamp 1676037725
transform 1 0 7360 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_78
timestamp 1676037725
transform 1 0 8280 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_98
timestamp 1676037725
transform 1 0 10120 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_111
timestamp 1676037725
transform 1 0 11316 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_135
timestamp 1676037725
transform 1 0 13524 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1676037725
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_147
timestamp 1676037725
transform 1 0 14628 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_160
timestamp 1676037725
transform 1 0 15824 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_167
timestamp 1676037725
transform 1 0 16468 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_171
timestamp 1676037725
transform 1 0 16836 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_183
timestamp 1676037725
transform 1 0 17940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1676037725
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_220
timestamp 1676037725
transform 1 0 21344 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_232
timestamp 1676037725
transform 1 0 22448 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_244
timestamp 1676037725
transform 1 0 23552 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1676037725
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1676037725
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1676037725
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1676037725
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1676037725
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1676037725
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1676037725
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1676037725
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1676037725
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1676037725
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1676037725
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1676037725
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1676037725
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1676037725
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_401
timestamp 1676037725
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_413
timestamp 1676037725
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1676037725
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1676037725
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1676037725
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1676037725
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1676037725
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1676037725
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1676037725
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1676037725
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1676037725
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1676037725
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1676037725
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_525
timestamp 1676037725
transform 1 0 49404 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_21
timestamp 1676037725
transform 1 0 3036 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_33
timestamp 1676037725
transform 1 0 4140 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_45
timestamp 1676037725
transform 1 0 5244 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_53
timestamp 1676037725
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_63
timestamp 1676037725
transform 1 0 6900 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_71
timestamp 1676037725
transform 1 0 7636 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_82
timestamp 1676037725
transform 1 0 8648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_57_109
timestamp 1676037725
transform 1 0 11132 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_138
timestamp 1676037725
transform 1 0 13800 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_151
timestamp 1676037725
transform 1 0 14996 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_166
timestamp 1676037725
transform 1 0 16376 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_184
timestamp 1676037725
transform 1 0 18032 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_197
timestamp 1676037725
transform 1 0 19228 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_209
timestamp 1676037725
transform 1 0 20332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_221
timestamp 1676037725
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1676037725
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1676037725
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1676037725
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1676037725
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1676037725
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1676037725
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1676037725
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1676037725
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1676037725
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1676037725
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1676037725
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1676037725
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1676037725
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1676037725
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1676037725
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1676037725
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1676037725
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1676037725
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1676037725
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1676037725
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1676037725
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1676037725
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1676037725
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1676037725
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1676037725
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1676037725
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1676037725
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1676037725
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1676037725
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_517
timestamp 1676037725
transform 1 0 48668 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_525
timestamp 1676037725
transform 1 0 49404 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_53
timestamp 1676037725
transform 1 0 5980 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_78
timestamp 1676037725
transform 1 0 8280 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_97
timestamp 1676037725
transform 1 0 10028 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_108
timestamp 1676037725
transform 1 0 11040 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_121
timestamp 1676037725
transform 1 0 12236 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_134
timestamp 1676037725
transform 1 0 13432 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_163
timestamp 1676037725
transform 1 0 16100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1676037725
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1676037725
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_220
timestamp 1676037725
transform 1 0 21344 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_232
timestamp 1676037725
transform 1 0 22448 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_244
timestamp 1676037725
transform 1 0 23552 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1676037725
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1676037725
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1676037725
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1676037725
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1676037725
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1676037725
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1676037725
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1676037725
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1676037725
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1676037725
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1676037725
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1676037725
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1676037725
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1676037725
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1676037725
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1676037725
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1676037725
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1676037725
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1676037725
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1676037725
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1676037725
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1676037725
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1676037725
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1676037725
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1676037725
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1676037725
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1676037725
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_525
timestamp 1676037725
transform 1 0 49404 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_21
timestamp 1676037725
transform 1 0 3036 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_33
timestamp 1676037725
transform 1 0 4140 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_45
timestamp 1676037725
transform 1 0 5244 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_53
timestamp 1676037725
transform 1 0 5980 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_69
timestamp 1676037725
transform 1 0 7452 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_79
timestamp 1676037725
transform 1 0 8372 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_92
timestamp 1676037725
transform 1 0 9568 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1676037725
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_59_139
timestamp 1676037725
transform 1 0 13892 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_145
timestamp 1676037725
transform 1 0 14444 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_166
timestamp 1676037725
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_197
timestamp 1676037725
transform 1 0 19228 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_201
timestamp 1676037725
transform 1 0 19596 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_222
timestamp 1676037725
transform 1 0 21528 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1676037725
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1676037725
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1676037725
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1676037725
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1676037725
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1676037725
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1676037725
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1676037725
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1676037725
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1676037725
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1676037725
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1676037725
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1676037725
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1676037725
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1676037725
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1676037725
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1676037725
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1676037725
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1676037725
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1676037725
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1676037725
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1676037725
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1676037725
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1676037725
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1676037725
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1676037725
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1676037725
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1676037725
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1676037725
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1676037725
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_517
timestamp 1676037725
transform 1 0 48668 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_525
timestamp 1676037725
transform 1 0 49404 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_21
timestamp 1676037725
transform 1 0 3036 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_56
timestamp 1676037725
transform 1 0 6256 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_69
timestamp 1676037725
transform 1 0 7452 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_82
timestamp 1676037725
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_114
timestamp 1676037725
transform 1 0 11592 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_125
timestamp 1676037725
transform 1 0 12604 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_138
timestamp 1676037725
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_166
timestamp 1676037725
transform 1 0 16376 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_194
timestamp 1676037725
transform 1 0 18952 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_205
timestamp 1676037725
transform 1 0 19964 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_215
timestamp 1676037725
transform 1 0 20884 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_228
timestamp 1676037725
transform 1 0 22080 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_240
timestamp 1676037725
transform 1 0 23184 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1676037725
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1676037725
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1676037725
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1676037725
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1676037725
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1676037725
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1676037725
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1676037725
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1676037725
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1676037725
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1676037725
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1676037725
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1676037725
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1676037725
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1676037725
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1676037725
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1676037725
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1676037725
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1676037725
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1676037725
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1676037725
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1676037725
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1676037725
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1676037725
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1676037725
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1676037725
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1676037725
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_525
timestamp 1676037725
transform 1 0 49404 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_39
timestamp 1676037725
transform 1 0 4692 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_54
timestamp 1676037725
transform 1 0 6072 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_61
timestamp 1676037725
transform 1 0 6716 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_71
timestamp 1676037725
transform 1 0 7636 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_84
timestamp 1676037725
transform 1 0 8832 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_97
timestamp 1676037725
transform 1 0 10028 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1676037725
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_119
timestamp 1676037725
transform 1 0 12052 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_123
timestamp 1676037725
transform 1 0 12420 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_144
timestamp 1676037725
transform 1 0 14352 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_156
timestamp 1676037725
transform 1 0 15456 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_166
timestamp 1676037725
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_181
timestamp 1676037725
transform 1 0 17756 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_198
timestamp 1676037725
transform 1 0 19320 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_222
timestamp 1676037725
transform 1 0 21528 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_238
timestamp 1676037725
transform 1 0 23000 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_250
timestamp 1676037725
transform 1 0 24104 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_262
timestamp 1676037725
transform 1 0 25208 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_274
timestamp 1676037725
transform 1 0 26312 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1676037725
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1676037725
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1676037725
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1676037725
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1676037725
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1676037725
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1676037725
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1676037725
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1676037725
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1676037725
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1676037725
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1676037725
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1676037725
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1676037725
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1676037725
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1676037725
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1676037725
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1676037725
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1676037725
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1676037725
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1676037725
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1676037725
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1676037725
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1676037725
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1676037725
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_517
timestamp 1676037725
transform 1 0 48668 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_525
timestamp 1676037725
transform 1 0 49404 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_21
timestamp 1676037725
transform 1 0 3036 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_56
timestamp 1676037725
transform 1 0 6256 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_69
timestamp 1676037725
transform 1 0 7452 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_82
timestamp 1676037725
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_110
timestamp 1676037725
transform 1 0 11224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_117
timestamp 1676037725
transform 1 0 11868 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_132
timestamp 1676037725
transform 1 0 13248 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_164
timestamp 1676037725
transform 1 0 16192 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_176
timestamp 1676037725
transform 1 0 17296 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_181
timestamp 1676037725
transform 1 0 17756 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1676037725
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_205
timestamp 1676037725
transform 1 0 19964 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_227
timestamp 1676037725
transform 1 0 21988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_239
timestamp 1676037725
transform 1 0 23092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1676037725
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1676037725
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1676037725
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1676037725
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1676037725
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1676037725
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1676037725
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1676037725
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1676037725
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1676037725
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1676037725
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1676037725
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1676037725
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1676037725
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1676037725
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1676037725
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1676037725
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1676037725
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1676037725
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1676037725
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1676037725
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1676037725
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1676037725
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1676037725
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1676037725
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1676037725
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1676037725
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1676037725
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_525
timestamp 1676037725
transform 1 0 49404 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_21
timestamp 1676037725
transform 1 0 3036 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_33
timestamp 1676037725
transform 1 0 4140 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_41
timestamp 1676037725
transform 1 0 4876 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_54
timestamp 1676037725
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_84
timestamp 1676037725
transform 1 0 8832 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_97
timestamp 1676037725
transform 1 0 10028 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1676037725
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_119
timestamp 1676037725
transform 1 0 12052 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_131
timestamp 1676037725
transform 1 0 13156 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_138
timestamp 1676037725
transform 1 0 13800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_142
timestamp 1676037725
transform 1 0 14168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_152
timestamp 1676037725
transform 1 0 15088 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_165
timestamp 1676037725
transform 1 0 16284 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_190
timestamp 1676037725
transform 1 0 18584 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_214
timestamp 1676037725
transform 1 0 20792 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1676037725
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_236
timestamp 1676037725
transform 1 0 22816 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_248
timestamp 1676037725
transform 1 0 23920 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_260
timestamp 1676037725
transform 1 0 25024 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_272
timestamp 1676037725
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1676037725
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1676037725
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1676037725
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1676037725
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1676037725
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1676037725
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1676037725
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1676037725
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1676037725
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1676037725
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1676037725
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1676037725
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1676037725
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1676037725
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1676037725
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1676037725
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1676037725
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1676037725
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1676037725
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1676037725
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1676037725
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1676037725
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1676037725
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1676037725
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1676037725
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_517
timestamp 1676037725
transform 1 0 48668 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_525
timestamp 1676037725
transform 1 0 49404 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_66
timestamp 1676037725
transform 1 0 7176 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_79
timestamp 1676037725
transform 1 0 8372 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1676037725
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_91
timestamp 1676037725
transform 1 0 9476 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_103
timestamp 1676037725
transform 1 0 10580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_111
timestamp 1676037725
transform 1 0 11316 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_117
timestamp 1676037725
transform 1 0 11868 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1676037725
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_64_167
timestamp 1676037725
transform 1 0 16468 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1676037725
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_209
timestamp 1676037725
transform 1 0 20332 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_231
timestamp 1676037725
transform 1 0 22356 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_244
timestamp 1676037725
transform 1 0 23552 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1676037725
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1676037725
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1676037725
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1676037725
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1676037725
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1676037725
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1676037725
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1676037725
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1676037725
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1676037725
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1676037725
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1676037725
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1676037725
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1676037725
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1676037725
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1676037725
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1676037725
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1676037725
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1676037725
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1676037725
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1676037725
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1676037725
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1676037725
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1676037725
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1676037725
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1676037725
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1676037725
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_525
timestamp 1676037725
transform 1 0 49404 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_21
timestamp 1676037725
transform 1 0 3036 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_37
timestamp 1676037725
transform 1 0 4508 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_54
timestamp 1676037725
transform 1 0 6072 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_61
timestamp 1676037725
transform 1 0 6716 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_82
timestamp 1676037725
transform 1 0 8648 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_97
timestamp 1676037725
transform 1 0 10028 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_65_110
timestamp 1676037725
transform 1 0 11224 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_118
timestamp 1676037725
transform 1 0 11960 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_133
timestamp 1676037725
transform 1 0 13340 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_141
timestamp 1676037725
transform 1 0 14076 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_145
timestamp 1676037725
transform 1 0 14444 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_166
timestamp 1676037725
transform 1 0 16376 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_192
timestamp 1676037725
transform 1 0 18768 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_204
timestamp 1676037725
transform 1 0 19872 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1676037725
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1676037725
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_233
timestamp 1676037725
transform 1 0 22540 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_244
timestamp 1676037725
transform 1 0 23552 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_256
timestamp 1676037725
transform 1 0 24656 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_268
timestamp 1676037725
transform 1 0 25760 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1676037725
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1676037725
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1676037725
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1676037725
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1676037725
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1676037725
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1676037725
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1676037725
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1676037725
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1676037725
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1676037725
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1676037725
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1676037725
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1676037725
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1676037725
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1676037725
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1676037725
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1676037725
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1676037725
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1676037725
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1676037725
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1676037725
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1676037725
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1676037725
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1676037725
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_517
timestamp 1676037725
transform 1 0 48668 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_525
timestamp 1676037725
transform 1 0 49404 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_21
timestamp 1676037725
transform 1 0 3036 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_37
timestamp 1676037725
transform 1 0 4508 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_54
timestamp 1676037725
transform 1 0 6072 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_82
timestamp 1676037725
transform 1 0 8648 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_110
timestamp 1676037725
transform 1 0 11224 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_138
timestamp 1676037725
transform 1 0 13800 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_163
timestamp 1676037725
transform 1 0 16100 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_187
timestamp 1676037725
transform 1 0 18308 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1676037725
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_209
timestamp 1676037725
transform 1 0 20332 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_231
timestamp 1676037725
transform 1 0 22356 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_248
timestamp 1676037725
transform 1 0 23920 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1676037725
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1676037725
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1676037725
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1676037725
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1676037725
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1676037725
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1676037725
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1676037725
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1676037725
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1676037725
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1676037725
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1676037725
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1676037725
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1676037725
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1676037725
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1676037725
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1676037725
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1676037725
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1676037725
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1676037725
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1676037725
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1676037725
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1676037725
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1676037725
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1676037725
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1676037725
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1676037725
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_525
timestamp 1676037725
transform 1 0 49404 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1676037725
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1676037725
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_39
timestamp 1676037725
transform 1 0 4692 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_67_54
timestamp 1676037725
transform 1 0 6072 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_63
timestamp 1676037725
transform 1 0 6900 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_76
timestamp 1676037725
transform 1 0 8096 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_100
timestamp 1676037725
transform 1 0 10304 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_67_110
timestamp 1676037725
transform 1 0 11224 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_119
timestamp 1676037725
transform 1 0 12052 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_141
timestamp 1676037725
transform 1 0 14076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_151
timestamp 1676037725
transform 1 0 14996 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_158
timestamp 1676037725
transform 1 0 15640 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_165
timestamp 1676037725
transform 1 0 16284 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_180
timestamp 1676037725
transform 1 0 17664 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_189
timestamp 1676037725
transform 1 0 18492 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_213
timestamp 1676037725
transform 1 0 20700 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_221
timestamp 1676037725
transform 1 0 21436 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_233
timestamp 1676037725
transform 1 0 22540 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_238
timestamp 1676037725
transform 1 0 23000 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_251
timestamp 1676037725
transform 1 0 24196 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_263
timestamp 1676037725
transform 1 0 25300 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_275
timestamp 1676037725
transform 1 0 26404 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1676037725
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1676037725
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1676037725
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1676037725
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1676037725
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1676037725
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1676037725
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1676037725
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1676037725
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1676037725
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1676037725
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1676037725
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1676037725
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1676037725
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1676037725
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1676037725
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1676037725
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1676037725
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1676037725
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1676037725
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1676037725
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1676037725
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1676037725
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1676037725
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1676037725
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1676037725
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_517
timestamp 1676037725
transform 1 0 48668 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_525
timestamp 1676037725
transform 1 0 49404 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_21
timestamp 1676037725
transform 1 0 3036 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_52
timestamp 1676037725
transform 1 0 5888 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_60
timestamp 1676037725
transform 1 0 6624 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_82
timestamp 1676037725
transform 1 0 8648 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_96
timestamp 1676037725
transform 1 0 9936 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_102
timestamp 1676037725
transform 1 0 10488 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_112
timestamp 1676037725
transform 1 0 11408 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_125
timestamp 1676037725
transform 1 0 12604 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_68_158
timestamp 1676037725
transform 1 0 15640 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_164
timestamp 1676037725
transform 1 0 16192 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_168
timestamp 1676037725
transform 1 0 16560 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_181
timestamp 1676037725
transform 1 0 17756 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_194
timestamp 1676037725
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_238
timestamp 1676037725
transform 1 0 23000 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_68_249
timestamp 1676037725
transform 1 0 24012 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1676037725
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1676037725
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1676037725
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1676037725
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1676037725
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1676037725
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1676037725
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1676037725
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1676037725
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1676037725
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1676037725
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1676037725
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1676037725
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1676037725
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1676037725
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1676037725
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1676037725
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1676037725
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1676037725
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1676037725
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1676037725
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1676037725
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1676037725
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1676037725
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1676037725
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1676037725
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1676037725
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_525
timestamp 1676037725
transform 1 0 49404 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_21
timestamp 1676037725
transform 1 0 3036 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_33
timestamp 1676037725
transform 1 0 4140 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_45
timestamp 1676037725
transform 1 0 5244 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_53
timestamp 1676037725
transform 1 0 5980 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_68
timestamp 1676037725
transform 1 0 7360 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_76
timestamp 1676037725
transform 1 0 8096 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_100
timestamp 1676037725
transform 1 0 10304 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_69_110
timestamp 1676037725
transform 1 0 11224 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_135
timestamp 1676037725
transform 1 0 13524 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_143
timestamp 1676037725
transform 1 0 14260 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_148
timestamp 1676037725
transform 1 0 14720 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1676037725
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1676037725
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_177
timestamp 1676037725
transform 1 0 17388 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_190
timestamp 1676037725
transform 1 0 18584 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_222
timestamp 1676037725
transform 1 0 21528 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_238
timestamp 1676037725
transform 1 0 23000 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_69_248
timestamp 1676037725
transform 1 0 23920 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1676037725
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1676037725
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1676037725
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1676037725
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1676037725
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1676037725
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1676037725
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1676037725
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1676037725
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1676037725
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1676037725
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1676037725
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1676037725
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1676037725
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1676037725
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1676037725
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1676037725
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1676037725
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1676037725
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1676037725
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1676037725
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1676037725
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1676037725
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1676037725
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1676037725
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1676037725
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1676037725
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1676037725
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_517
timestamp 1676037725
transform 1 0 48668 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_525
timestamp 1676037725
transform 1 0 49404 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1676037725
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_65
timestamp 1676037725
transform 1 0 7084 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_69
timestamp 1676037725
transform 1 0 7452 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_82
timestamp 1676037725
transform 1 0 8648 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_70_96
timestamp 1676037725
transform 1 0 9936 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_119
timestamp 1676037725
transform 1 0 12052 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_125
timestamp 1676037725
transform 1 0 12604 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_138
timestamp 1676037725
transform 1 0 13800 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_163
timestamp 1676037725
transform 1 0 16100 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_194
timestamp 1676037725
transform 1 0 18952 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_205
timestamp 1676037725
transform 1 0 19964 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_218
timestamp 1676037725
transform 1 0 21160 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_242
timestamp 1676037725
transform 1 0 23368 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_248
timestamp 1676037725
transform 1 0 23920 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_253
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_70_264
timestamp 1676037725
transform 1 0 25392 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_270
timestamp 1676037725
transform 1 0 25944 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_282
timestamp 1676037725
transform 1 0 27048 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_294
timestamp 1676037725
transform 1 0 28152 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_306
timestamp 1676037725
transform 1 0 29256 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1676037725
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1676037725
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1676037725
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1676037725
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1676037725
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1676037725
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1676037725
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1676037725
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1676037725
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1676037725
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1676037725
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1676037725
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1676037725
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1676037725
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1676037725
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1676037725
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1676037725
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1676037725
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1676037725
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1676037725
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1676037725
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1676037725
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_525
timestamp 1676037725
transform 1 0 49404 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_21
timestamp 1676037725
transform 1 0 3036 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_33
timestamp 1676037725
transform 1 0 4140 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_45
timestamp 1676037725
transform 1 0 5244 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_53
timestamp 1676037725
transform 1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_64
timestamp 1676037725
transform 1 0 6992 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_72
timestamp 1676037725
transform 1 0 7728 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_86
timestamp 1676037725
transform 1 0 9016 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_110
timestamp 1676037725
transform 1 0 11224 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_118
timestamp 1676037725
transform 1 0 11960 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_142
timestamp 1676037725
transform 1 0 14168 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_166
timestamp 1676037725
transform 1 0 16376 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_180
timestamp 1676037725
transform 1 0 17664 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_188
timestamp 1676037725
transform 1 0 18400 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_193
timestamp 1676037725
transform 1 0 18860 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_206
timestamp 1676037725
transform 1 0 20056 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_212
timestamp 1676037725
transform 1 0 20608 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_235
timestamp 1676037725
transform 1 0 22724 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_248
timestamp 1676037725
transform 1 0 23920 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_263
timestamp 1676037725
transform 1 0 25300 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_275
timestamp 1676037725
transform 1 0 26404 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1676037725
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1676037725
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1676037725
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1676037725
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1676037725
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1676037725
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1676037725
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1676037725
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1676037725
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1676037725
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1676037725
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1676037725
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1676037725
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1676037725
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1676037725
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1676037725
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1676037725
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1676037725
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1676037725
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1676037725
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1676037725
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1676037725
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1676037725
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1676037725
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1676037725
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1676037725
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_517
timestamp 1676037725
transform 1 0 48668 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_525
timestamp 1676037725
transform 1 0 49404 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_72_21
timestamp 1676037725
transform 1 0 3036 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_37
timestamp 1676037725
transform 1 0 4508 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_42
timestamp 1676037725
transform 1 0 4968 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_54
timestamp 1676037725
transform 1 0 6072 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_72_61
timestamp 1676037725
transform 1 0 6716 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_73
timestamp 1676037725
transform 1 0 7820 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_72_82
timestamp 1676037725
transform 1 0 8648 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_121
timestamp 1676037725
transform 1 0 12236 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_138
timestamp 1676037725
transform 1 0 13800 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_152
timestamp 1676037725
transform 1 0 15088 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_176
timestamp 1676037725
transform 1 0 17296 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_180
timestamp 1676037725
transform 1 0 17664 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_205
timestamp 1676037725
transform 1 0 19964 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_208
timestamp 1676037725
transform 1 0 20240 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_225
timestamp 1676037725
transform 1 0 21804 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_236
timestamp 1676037725
transform 1 0 22816 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_240
timestamp 1676037725
transform 1 0 23184 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_72_250
timestamp 1676037725
transform 1 0 24104 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1676037725
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1676037725
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1676037725
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1676037725
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1676037725
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1676037725
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1676037725
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1676037725
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1676037725
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1676037725
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1676037725
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1676037725
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1676037725
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1676037725
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1676037725
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1676037725
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1676037725
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1676037725
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1676037725
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1676037725
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1676037725
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1676037725
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1676037725
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1676037725
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1676037725
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1676037725
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1676037725
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_525
timestamp 1676037725
transform 1 0 49404 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1676037725
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1676037725
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_39
timestamp 1676037725
transform 1 0 4692 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_44
timestamp 1676037725
transform 1 0 5152 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_81
timestamp 1676037725
transform 1 0 8556 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_103
timestamp 1676037725
transform 1 0 10580 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_110
timestamp 1676037725
transform 1 0 11224 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_126
timestamp 1676037725
transform 1 0 12696 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_139
timestamp 1676037725
transform 1 0 13892 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_145
timestamp 1676037725
transform 1 0 14444 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_166
timestamp 1676037725
transform 1 0 16376 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_178
timestamp 1676037725
transform 1 0 17480 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_185
timestamp 1676037725
transform 1 0 18124 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_193
timestamp 1676037725
transform 1 0 18860 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_199
timestamp 1676037725
transform 1 0 19412 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_209
timestamp 1676037725
transform 1 0 20332 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_222
timestamp 1676037725
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_251
timestamp 1676037725
transform 1 0 24196 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_263
timestamp 1676037725
transform 1 0 25300 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_275
timestamp 1676037725
transform 1 0 26404 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1676037725
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1676037725
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1676037725
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1676037725
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1676037725
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1676037725
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1676037725
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1676037725
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1676037725
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1676037725
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1676037725
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1676037725
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1676037725
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1676037725
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1676037725
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1676037725
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1676037725
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1676037725
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1676037725
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1676037725
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1676037725
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1676037725
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1676037725
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1676037725
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1676037725
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1676037725
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_517
timestamp 1676037725
transform 1 0 48668 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_525
timestamp 1676037725
transform 1 0 49404 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_21
timestamp 1676037725
transform 1 0 3036 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1676037725
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_53
timestamp 1676037725
transform 1 0 5980 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_82
timestamp 1676037725
transform 1 0 8648 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_85
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_90
timestamp 1676037725
transform 1 0 9384 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_114
timestamp 1676037725
transform 1 0 11592 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_138
timestamp 1676037725
transform 1 0 13800 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_74_153
timestamp 1676037725
transform 1 0 15180 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_159
timestamp 1676037725
transform 1 0 15732 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_180
timestamp 1676037725
transform 1 0 17664 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_186
timestamp 1676037725
transform 1 0 18216 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_194
timestamp 1676037725
transform 1 0 18952 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_208
timestamp 1676037725
transform 1 0 20240 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_234
timestamp 1676037725
transform 1 0 22632 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_246
timestamp 1676037725
transform 1 0 23736 0 1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1676037725
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1676037725
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1676037725
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1676037725
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1676037725
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1676037725
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1676037725
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1676037725
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1676037725
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1676037725
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1676037725
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1676037725
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1676037725
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1676037725
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1676037725
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1676037725
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1676037725
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1676037725
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1676037725
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1676037725
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1676037725
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1676037725
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1676037725
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1676037725
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1676037725
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1676037725
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1676037725
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_525
timestamp 1676037725
transform 1 0 49404 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_21
timestamp 1676037725
transform 1 0 3036 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_33
timestamp 1676037725
transform 1 0 4140 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_45
timestamp 1676037725
transform 1 0 5244 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_53
timestamp 1676037725
transform 1 0 5980 0 -1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_81
timestamp 1676037725
transform 1 0 8556 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_85
timestamp 1676037725
transform 1 0 8924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_90
timestamp 1676037725
transform 1 0 9384 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_97
timestamp 1676037725
transform 1 0 10028 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_110
timestamp 1676037725
transform 1 0 11224 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_124
timestamp 1676037725
transform 1 0 12512 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_132
timestamp 1676037725
transform 1 0 13248 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_137
timestamp 1676037725
transform 1 0 13708 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_145
timestamp 1676037725
transform 1 0 14444 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_158
timestamp 1676037725
transform 1 0 15640 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_162
timestamp 1676037725
transform 1 0 16008 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_166
timestamp 1676037725
transform 1 0 16376 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_169
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_174
timestamp 1676037725
transform 1 0 17112 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_181
timestamp 1676037725
transform 1 0 17756 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_205
timestamp 1676037725
transform 1 0 19964 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_222
timestamp 1676037725
transform 1 0 21528 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_236
timestamp 1676037725
transform 1 0 22816 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_248
timestamp 1676037725
transform 1 0 23920 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_260
timestamp 1676037725
transform 1 0 25024 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_272
timestamp 1676037725
transform 1 0 26128 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1676037725
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1676037725
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1676037725
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1676037725
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1676037725
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1676037725
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1676037725
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1676037725
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1676037725
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1676037725
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1676037725
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1676037725
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1676037725
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1676037725
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1676037725
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1676037725
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1676037725
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1676037725
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1676037725
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1676037725
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1676037725
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1676037725
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1676037725
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1676037725
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1676037725
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_517
timestamp 1676037725
transform 1 0 48668 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_525
timestamp 1676037725
transform 1 0 49404 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1676037725
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1676037725
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_45
timestamp 1676037725
transform 1 0 5244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_57
timestamp 1676037725
transform 1 0 6348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_69
timestamp 1676037725
transform 1 0 7452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_81
timestamp 1676037725
transform 1 0 8556 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_97
timestamp 1676037725
transform 1 0 10028 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_101
timestamp 1676037725
transform 1 0 10396 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_106
timestamp 1676037725
transform 1 0 10856 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_119
timestamp 1676037725
transform 1 0 12052 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_130
timestamp 1676037725
transform 1 0 13064 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_76_137
timestamp 1676037725
transform 1 0 13708 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_76_141
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_146
timestamp 1676037725
transform 1 0 14536 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_154
timestamp 1676037725
transform 1 0 15272 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_176
timestamp 1676037725
transform 1 0 17296 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_183
timestamp 1676037725
transform 1 0 17940 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_194
timestamp 1676037725
transform 1 0 18952 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_209
timestamp 1676037725
transform 1 0 20332 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_76_216
timestamp 1676037725
transform 1 0 20976 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_222
timestamp 1676037725
transform 1 0 21528 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_226
timestamp 1676037725
transform 1 0 21896 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_250
timestamp 1676037725
transform 1 0 24104 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_264
timestamp 1676037725
transform 1 0 25392 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_276
timestamp 1676037725
transform 1 0 26496 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_280
timestamp 1676037725
transform 1 0 26864 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_293
timestamp 1676037725
transform 1 0 28060 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_299
timestamp 1676037725
transform 1 0 28612 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1676037725
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1676037725
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1676037725
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1676037725
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1676037725
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1676037725
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1676037725
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1676037725
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1676037725
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1676037725
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1676037725
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1676037725
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1676037725
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1676037725
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1676037725
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1676037725
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1676037725
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1676037725
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1676037725
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1676037725
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1676037725
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1676037725
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1676037725
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_525
timestamp 1676037725
transform 1 0 49404 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_21
timestamp 1676037725
transform 1 0 3036 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_25
timestamp 1676037725
transform 1 0 3404 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_30
timestamp 1676037725
transform 1 0 3864 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_34
timestamp 1676037725
transform 1 0 4232 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1676037725
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1676037725
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1676037725
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1676037725
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_84
timestamp 1676037725
transform 1 0 8832 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_92
timestamp 1676037725
transform 1 0 9568 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_104
timestamp 1676037725
transform 1 0 10672 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_77_109
timestamp 1676037725
transform 1 0 11132 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_77_113
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_119
timestamp 1676037725
transform 1 0 12052 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_123
timestamp 1676037725
transform 1 0 12420 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_130
timestamp 1676037725
transform 1 0 13064 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_142
timestamp 1676037725
transform 1 0 14168 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_154
timestamp 1676037725
transform 1 0 15272 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_166
timestamp 1676037725
transform 1 0 16376 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_77_174
timestamp 1676037725
transform 1 0 17112 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_181
timestamp 1676037725
transform 1 0 17756 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_188
timestamp 1676037725
transform 1 0 18400 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_201
timestamp 1676037725
transform 1 0 19596 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_207
timestamp 1676037725
transform 1 0 20148 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1676037725
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1676037725
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_230
timestamp 1676037725
transform 1 0 22264 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_242
timestamp 1676037725
transform 1 0 23368 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_254
timestamp 1676037725
transform 1 0 24472 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_77_278
timestamp 1676037725
transform 1 0 26680 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1676037725
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1676037725
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1676037725
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1676037725
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1676037725
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1676037725
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1676037725
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1676037725
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1676037725
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1676037725
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1676037725
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1676037725
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1676037725
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1676037725
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1676037725
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1676037725
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1676037725
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1676037725
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1676037725
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1676037725
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1676037725
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1676037725
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1676037725
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1676037725
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1676037725
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_517
timestamp 1676037725
transform 1 0 48668 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_525
timestamp 1676037725
transform 1 0 49404 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_21
timestamp 1676037725
transform 1 0 3036 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_35
timestamp 1676037725
transform 1 0 4324 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_43
timestamp 1676037725
transform 1 0 5060 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_55
timestamp 1676037725
transform 1 0 6164 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_67
timestamp 1676037725
transform 1 0 7268 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_79
timestamp 1676037725
transform 1 0 8372 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1676037725
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_90
timestamp 1676037725
transform 1 0 9384 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_97
timestamp 1676037725
transform 1 0 10028 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_104
timestamp 1676037725
transform 1 0 10672 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_111
timestamp 1676037725
transform 1 0 11316 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_118
timestamp 1676037725
transform 1 0 11960 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_125
timestamp 1676037725
transform 1 0 12604 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_129
timestamp 1676037725
transform 1 0 12972 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1676037725
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1676037725
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_146
timestamp 1676037725
transform 1 0 14536 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_155
timestamp 1676037725
transform 1 0 15364 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_168
timestamp 1676037725
transform 1 0 16560 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_181
timestamp 1676037725
transform 1 0 17756 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_78_194
timestamp 1676037725
transform 1 0 18952 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_219
timestamp 1676037725
transform 1 0 21252 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_232
timestamp 1676037725
transform 1 0 22448 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_244
timestamp 1676037725
transform 1 0 23552 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_265
timestamp 1676037725
transform 1 0 25484 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_275
timestamp 1676037725
transform 1 0 26404 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_288
timestamp 1676037725
transform 1 0 27600 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_294
timestamp 1676037725
transform 1 0 28152 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_306
timestamp 1676037725
transform 1 0 29256 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1676037725
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1676037725
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1676037725
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1676037725
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1676037725
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1676037725
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1676037725
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1676037725
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1676037725
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1676037725
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1676037725
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1676037725
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1676037725
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1676037725
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1676037725
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1676037725
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1676037725
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1676037725
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1676037725
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1676037725
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1676037725
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1676037725
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_525
timestamp 1676037725
transform 1 0 49404 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_3
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_11
timestamp 1676037725
transform 1 0 2116 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_18
timestamp 1676037725
transform 1 0 2760 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_26
timestamp 1676037725
transform 1 0 3496 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_31
timestamp 1676037725
transform 1 0 3956 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1676037725
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1676037725
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1676037725
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_69
timestamp 1676037725
transform 1 0 7452 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_73
timestamp 1676037725
transform 1 0 7820 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_77
timestamp 1676037725
transform 1 0 8188 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_85
timestamp 1676037725
transform 1 0 8924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_89
timestamp 1676037725
transform 1 0 9292 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_101
timestamp 1676037725
transform 1 0 10396 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_109
timestamp 1676037725
transform 1 0 11132 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_118
timestamp 1676037725
transform 1 0 11960 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_127
timestamp 1676037725
transform 1 0 12788 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_139
timestamp 1676037725
transform 1 0 13892 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_146
timestamp 1676037725
transform 1 0 14536 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_153
timestamp 1676037725
transform 1 0 15180 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_166
timestamp 1676037725
transform 1 0 16376 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_188
timestamp 1676037725
transform 1 0 18400 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_192
timestamp 1676037725
transform 1 0 18768 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_202
timestamp 1676037725
transform 1 0 19688 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1676037725
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1676037725
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_79_230
timestamp 1676037725
transform 1 0 22264 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_256
timestamp 1676037725
transform 1 0 24656 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_268
timestamp 1676037725
transform 1 0 25760 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1676037725
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1676037725
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1676037725
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1676037725
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1676037725
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1676037725
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1676037725
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1676037725
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1676037725
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1676037725
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1676037725
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1676037725
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1676037725
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1676037725
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1676037725
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1676037725
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1676037725
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1676037725
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1676037725
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1676037725
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1676037725
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1676037725
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1676037725
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1676037725
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1676037725
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_517
timestamp 1676037725
transform 1 0 48668 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_525
timestamp 1676037725
transform 1 0 49404 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_21
timestamp 1676037725
transform 1 0 3036 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_35
timestamp 1676037725
transform 1 0 4324 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_47
timestamp 1676037725
transform 1 0 5428 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_59
timestamp 1676037725
transform 1 0 6532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_71
timestamp 1676037725
transform 1 0 7636 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_78
timestamp 1676037725
transform 1 0 8280 0 1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_109
timestamp 1676037725
transform 1 0 11132 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_113
timestamp 1676037725
transform 1 0 11500 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_125
timestamp 1676037725
transform 1 0 12604 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_133
timestamp 1676037725
transform 1 0 13340 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_138
timestamp 1676037725
transform 1 0 13800 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_141
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_145
timestamp 1676037725
transform 1 0 14444 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_166
timestamp 1676037725
transform 1 0 16376 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_194
timestamp 1676037725
transform 1 0 18952 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_202
timestamp 1676037725
transform 1 0 19688 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_226
timestamp 1676037725
transform 1 0 21896 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_80_250
timestamp 1676037725
transform 1 0 24104 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1676037725
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1676037725
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1676037725
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1676037725
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1676037725
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1676037725
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1676037725
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1676037725
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1676037725
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1676037725
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1676037725
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1676037725
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1676037725
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1676037725
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1676037725
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1676037725
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1676037725
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1676037725
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1676037725
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1676037725
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1676037725
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1676037725
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1676037725
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1676037725
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1676037725
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_501
timestamp 1676037725
transform 1 0 47196 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_525
timestamp 1676037725
transform 1 0 49404 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_21
timestamp 1676037725
transform 1 0 3036 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_81_29
timestamp 1676037725
transform 1 0 3772 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_81_36
timestamp 1676037725
transform 1 0 4416 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_81_46
timestamp 1676037725
transform 1 0 5336 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_54
timestamp 1676037725
transform 1 0 6072 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1676037725
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1676037725
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1676037725
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_105
timestamp 1676037725
transform 1 0 10764 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_110
timestamp 1676037725
transform 1 0 11224 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_125
timestamp 1676037725
transform 1 0 12604 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_129
timestamp 1676037725
transform 1 0 12972 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_142
timestamp 1676037725
transform 1 0 14168 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_166
timestamp 1676037725
transform 1 0 16376 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_174
timestamp 1676037725
transform 1 0 17112 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_198
timestamp 1676037725
transform 1 0 19320 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_222
timestamp 1676037725
transform 1 0 21528 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_251
timestamp 1676037725
transform 1 0 24196 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_257
timestamp 1676037725
transform 1 0 24748 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_270
timestamp 1676037725
transform 1 0 25944 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_278
timestamp 1676037725
transform 1 0 26680 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1676037725
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1676037725
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1676037725
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1676037725
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1676037725
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1676037725
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1676037725
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1676037725
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1676037725
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1676037725
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1676037725
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1676037725
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1676037725
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1676037725
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1676037725
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1676037725
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1676037725
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1676037725
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1676037725
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1676037725
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1676037725
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1676037725
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1676037725
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1676037725
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1676037725
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_81_517
timestamp 1676037725
transform 1 0 48668 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_525
timestamp 1676037725
transform 1 0 49404 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1676037725
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1676037725
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_112
timestamp 1676037725
transform 1 0 11408 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_125
timestamp 1676037725
transform 1 0 12604 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_138
timestamp 1676037725
transform 1 0 13800 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_163
timestamp 1676037725
transform 1 0 16100 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_170
timestamp 1676037725
transform 1 0 16744 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_194
timestamp 1676037725
transform 1 0 18952 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_197
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_221
timestamp 1676037725
transform 1 0 21436 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_229
timestamp 1676037725
transform 1 0 22172 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_250
timestamp 1676037725
transform 1 0 24104 0 1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1676037725
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1676037725
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1676037725
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1676037725
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1676037725
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1676037725
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1676037725
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1676037725
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1676037725
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1676037725
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1676037725
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1676037725
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1676037725
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1676037725
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1676037725
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1676037725
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1676037725
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1676037725
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1676037725
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1676037725
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1676037725
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1676037725
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1676037725
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1676037725
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1676037725
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1676037725
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1676037725
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_82_525
timestamp 1676037725
transform 1 0 49404 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_21
timestamp 1676037725
transform 1 0 3036 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_33
timestamp 1676037725
transform 1 0 4140 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_45
timestamp 1676037725
transform 1 0 5244 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_53
timestamp 1676037725
transform 1 0 5980 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_96
timestamp 1676037725
transform 1 0 9936 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_103
timestamp 1676037725
transform 1 0 10580 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_110
timestamp 1676037725
transform 1 0 11224 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_118
timestamp 1676037725
transform 1 0 11960 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_130
timestamp 1676037725
transform 1 0 13064 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_83_153
timestamp 1676037725
transform 1 0 15180 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_166
timestamp 1676037725
transform 1 0 16376 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_83_197
timestamp 1676037725
transform 1 0 19228 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_201
timestamp 1676037725
transform 1 0 19596 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_222
timestamp 1676037725
transform 1 0 21528 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_83_230
timestamp 1676037725
transform 1 0 22264 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_83_258
timestamp 1676037725
transform 1 0 24840 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_264
timestamp 1676037725
transform 1 0 25392 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_83_277
timestamp 1676037725
transform 1 0 26588 0 -1 47872
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1676037725
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1676037725
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1676037725
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1676037725
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1676037725
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1676037725
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1676037725
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1676037725
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1676037725
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1676037725
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1676037725
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1676037725
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1676037725
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1676037725
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1676037725
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1676037725
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1676037725
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1676037725
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1676037725
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1676037725
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1676037725
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1676037725
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1676037725
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1676037725
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1676037725
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_517
timestamp 1676037725
transform 1 0 48668 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_525
timestamp 1676037725
transform 1 0 49404 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_84_21
timestamp 1676037725
transform 1 0 3036 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1676037725
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1676037725
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_121
timestamp 1676037725
transform 1 0 12236 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_125
timestamp 1676037725
transform 1 0 12604 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_138
timestamp 1676037725
transform 1 0 13800 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_84_167
timestamp 1676037725
transform 1 0 16468 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_173
timestamp 1676037725
transform 1 0 17020 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_194
timestamp 1676037725
transform 1 0 18952 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_210
timestamp 1676037725
transform 1 0 20424 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_216
timestamp 1676037725
transform 1 0 20976 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_220
timestamp 1676037725
transform 1 0 21344 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_228
timestamp 1676037725
transform 1 0 22080 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_250
timestamp 1676037725
transform 1 0 24104 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_84_253
timestamp 1676037725
transform 1 0 24380 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_261
timestamp 1676037725
transform 1 0 25116 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_264
timestamp 1676037725
transform 1 0 25392 0 1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1676037725
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1676037725
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1676037725
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1676037725
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1676037725
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1676037725
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1676037725
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1676037725
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1676037725
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1676037725
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1676037725
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1676037725
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1676037725
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1676037725
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1676037725
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1676037725
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1676037725
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1676037725
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1676037725
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1676037725
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1676037725
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1676037725
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1676037725
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1676037725
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1676037725
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_513
timestamp 1676037725
transform 1 0 48300 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_84_525
timestamp 1676037725
transform 1 0 49404 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1676037725
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1676037725
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1676037725
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1676037725
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1676037725
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1676037725
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_81
timestamp 1676037725
transform 1 0 8556 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_89
timestamp 1676037725
transform 1 0 9292 0 -1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_85_95
timestamp 1676037725
transform 1 0 9844 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_107
timestamp 1676037725
transform 1 0 10948 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1676037725
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_121
timestamp 1676037725
transform 1 0 12236 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_125
timestamp 1676037725
transform 1 0 12604 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_149
timestamp 1676037725
transform 1 0 14812 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_166
timestamp 1676037725
transform 1 0 16376 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_175
timestamp 1676037725
transform 1 0 17204 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_185
timestamp 1676037725
transform 1 0 18124 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_85_202
timestamp 1676037725
transform 1 0 19688 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_206
timestamp 1676037725
transform 1 0 20056 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_210
timestamp 1676037725
transform 1 0 20424 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_85_247
timestamp 1676037725
transform 1 0 23828 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_261
timestamp 1676037725
transform 1 0 25116 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_274
timestamp 1676037725
transform 1 0 26312 0 -1 48960
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1676037725
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1676037725
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1676037725
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1676037725
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1676037725
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1676037725
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1676037725
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1676037725
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1676037725
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1676037725
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1676037725
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1676037725
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1676037725
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1676037725
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1676037725
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1676037725
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1676037725
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1676037725
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1676037725
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1676037725
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1676037725
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1676037725
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1676037725
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1676037725
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1676037725
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_517
timestamp 1676037725
transform 1 0 48668 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_525
timestamp 1676037725
transform 1 0 49404 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_86_21
timestamp 1676037725
transform 1 0 3036 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1676037725
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1676037725
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1676037725
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1676037725
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1676037725
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1676037725
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_109
timestamp 1676037725
transform 1 0 11132 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_117
timestamp 1676037725
transform 1 0 11868 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_125
timestamp 1676037725
transform 1 0 12604 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_138
timestamp 1676037725
transform 1 0 13800 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_147
timestamp 1676037725
transform 1 0 14628 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_157
timestamp 1676037725
transform 1 0 15548 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_170
timestamp 1676037725
transform 1 0 16744 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_194
timestamp 1676037725
transform 1 0 18952 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_86_203
timestamp 1676037725
transform 1 0 19780 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_86_218
timestamp 1676037725
transform 1 0 21160 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_242
timestamp 1676037725
transform 1 0 23368 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_250
timestamp 1676037725
transform 1 0 24104 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_86_262
timestamp 1676037725
transform 1 0 25208 0 1 48960
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_86_274
timestamp 1676037725
transform 1 0 26312 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_286
timestamp 1676037725
transform 1 0 27416 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_298
timestamp 1676037725
transform 1 0 28520 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_306
timestamp 1676037725
transform 1 0 29256 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1676037725
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1676037725
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1676037725
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1676037725
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1676037725
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1676037725
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1676037725
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1676037725
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1676037725
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1676037725
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1676037725
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1676037725
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1676037725
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1676037725
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1676037725
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1676037725
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1676037725
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1676037725
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1676037725
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1676037725
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1676037725
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1676037725
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_86_525
timestamp 1676037725
transform 1 0 49404 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_21
timestamp 1676037725
transform 1 0 3036 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_33
timestamp 1676037725
transform 1 0 4140 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_45
timestamp 1676037725
transform 1 0 5244 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_87_53
timestamp 1676037725
transform 1 0 5980 0 -1 50048
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1676037725
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1676037725
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1676037725
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1676037725
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1676037725
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_121
timestamp 1676037725
transform 1 0 12236 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_129
timestamp 1676037725
transform 1 0 12972 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_137
timestamp 1676037725
transform 1 0 13708 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1676037725
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1676037725
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_173
timestamp 1676037725
transform 1 0 17020 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_183
timestamp 1676037725
transform 1 0 17940 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_87_198
timestamp 1676037725
transform 1 0 19320 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_222
timestamp 1676037725
transform 1 0 21528 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_238
timestamp 1676037725
transform 1 0 23000 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_87_251
timestamp 1676037725
transform 1 0 24196 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_263
timestamp 1676037725
transform 1 0 25300 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_275
timestamp 1676037725
transform 1 0 26404 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1676037725
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1676037725
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1676037725
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1676037725
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1676037725
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1676037725
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1676037725
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1676037725
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1676037725
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1676037725
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1676037725
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1676037725
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1676037725
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1676037725
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1676037725
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1676037725
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1676037725
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1676037725
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1676037725
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1676037725
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1676037725
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1676037725
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1676037725
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1676037725
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1676037725
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1676037725
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_517
timestamp 1676037725
transform 1 0 48668 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_525
timestamp 1676037725
transform 1 0 49404 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1676037725
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1676037725
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1676037725
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1676037725
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1676037725
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1676037725
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1676037725
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1676037725
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1676037725
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_109
timestamp 1676037725
transform 1 0 11132 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_118
timestamp 1676037725
transform 1 0 11960 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_88_130
timestamp 1676037725
transform 1 0 13064 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_88_137
timestamp 1676037725
transform 1 0 13708 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_88_164
timestamp 1676037725
transform 1 0 16192 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_172
timestamp 1676037725
transform 1 0 16928 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_194
timestamp 1676037725
transform 1 0 18952 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_201
timestamp 1676037725
transform 1 0 19596 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_211
timestamp 1676037725
transform 1 0 20516 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_88_235
timestamp 1676037725
transform 1 0 22724 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_88_250
timestamp 1676037725
transform 1 0 24104 0 1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1676037725
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1676037725
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1676037725
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1676037725
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1676037725
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1676037725
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1676037725
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1676037725
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1676037725
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1676037725
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1676037725
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1676037725
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1676037725
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1676037725
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1676037725
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1676037725
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1676037725
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1676037725
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1676037725
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1676037725
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1676037725
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1676037725
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1676037725
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1676037725
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1676037725
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1676037725
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_513
timestamp 1676037725
transform 1 0 48300 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_525
timestamp 1676037725
transform 1 0 49404 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_21
timestamp 1676037725
transform 1 0 3036 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_33
timestamp 1676037725
transform 1 0 4140 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_45
timestamp 1676037725
transform 1 0 5244 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_53
timestamp 1676037725
transform 1 0 5980 0 -1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_69
timestamp 1676037725
transform 1 0 7452 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_77
timestamp 1676037725
transform 1 0 8188 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_82
timestamp 1676037725
transform 1 0 8648 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_89_89
timestamp 1676037725
transform 1 0 9292 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_101
timestamp 1676037725
transform 1 0 10396 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_109
timestamp 1676037725
transform 1 0 11132 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_119
timestamp 1676037725
transform 1 0 12052 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_123
timestamp 1676037725
transform 1 0 12420 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_130
timestamp 1676037725
transform 1 0 13064 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_138
timestamp 1676037725
transform 1 0 13800 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_166
timestamp 1676037725
transform 1 0 16376 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_89_193
timestamp 1676037725
transform 1 0 18860 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_201
timestamp 1676037725
transform 1 0 19596 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_212
timestamp 1676037725
transform 1 0 20608 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_89_219
timestamp 1676037725
transform 1 0 21252 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_237
timestamp 1676037725
transform 1 0 22908 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_247
timestamp 1676037725
transform 1 0 23828 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_259
timestamp 1676037725
transform 1 0 24932 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_271
timestamp 1676037725
transform 1 0 26036 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1676037725
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1676037725
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1676037725
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1676037725
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1676037725
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1676037725
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1676037725
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1676037725
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1676037725
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1676037725
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1676037725
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1676037725
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1676037725
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_89_393
timestamp 1676037725
transform 1 0 37260 0 -1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_416
timestamp 1676037725
transform 1 0 39376 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_428
timestamp 1676037725
transform 1 0 40480 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_440
timestamp 1676037725
transform 1 0 41584 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1676037725
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1676037725
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1676037725
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1676037725
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1676037725
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1676037725
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1676037725
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_517
timestamp 1676037725
transform 1 0 48668 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_525
timestamp 1676037725
transform 1 0 49404 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_90_21
timestamp 1676037725
transform 1 0 3036 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1676037725
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1676037725
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1676037725
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_65
timestamp 1676037725
transform 1 0 7084 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_90_74
timestamp 1676037725
transform 1 0 7912 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_90_82
timestamp 1676037725
transform 1 0 8648 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_91
timestamp 1676037725
transform 1 0 9476 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_90_103
timestamp 1676037725
transform 1 0 10580 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1676037725
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1676037725
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_133
timestamp 1676037725
transform 1 0 13340 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_138
timestamp 1676037725
transform 1 0 13800 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_147
timestamp 1676037725
transform 1 0 14628 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_151
timestamp 1676037725
transform 1 0 14996 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_159
timestamp 1676037725
transform 1 0 15732 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_180
timestamp 1676037725
transform 1 0 17664 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_90_193
timestamp 1676037725
transform 1 0 18860 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1676037725
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1676037725
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1676037725
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1676037725
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1676037725
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1676037725
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1676037725
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1676037725
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1676037725
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1676037725
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1676037725
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1676037725
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1676037725
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1676037725
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1676037725
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1676037725
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1676037725
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1676037725
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1676037725
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1676037725
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1676037725
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1676037725
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1676037725
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1676037725
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1676037725
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1676037725
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1676037725
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1676037725
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1676037725
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1676037725
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1676037725
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1676037725
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_90_525
timestamp 1676037725
transform 1 0 49404 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1676037725
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1676037725
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1676037725
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1676037725
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1676037725
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_91_69
timestamp 1676037725
transform 1 0 7452 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_91_75
timestamp 1676037725
transform 1 0 8004 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_91_83
timestamp 1676037725
transform 1 0 8740 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_91
timestamp 1676037725
transform 1 0 9476 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_96
timestamp 1676037725
transform 1 0 9936 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_91_103
timestamp 1676037725
transform 1 0 10580 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1676037725
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1676037725
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1676037725
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_149
timestamp 1676037725
transform 1 0 14812 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_91_160
timestamp 1676037725
transform 1 0 15824 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_91_174
timestamp 1676037725
transform 1 0 17112 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_178
timestamp 1676037725
transform 1 0 17480 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_182
timestamp 1676037725
transform 1 0 17848 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_190
timestamp 1676037725
transform 1 0 18584 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_196
timestamp 1676037725
transform 1 0 19136 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_208
timestamp 1676037725
transform 1 0 20240 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_220
timestamp 1676037725
transform 1 0 21344 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1676037725
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1676037725
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1676037725
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1676037725
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1676037725
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1676037725
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1676037725
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1676037725
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1676037725
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1676037725
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1676037725
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1676037725
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1676037725
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1676037725
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1676037725
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1676037725
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1676037725
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1676037725
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1676037725
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1676037725
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1676037725
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1676037725
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1676037725
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1676037725
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1676037725
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1676037725
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1676037725
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1676037725
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1676037725
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_517
timestamp 1676037725
transform 1 0 48668 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_525
timestamp 1676037725
transform 1 0 49404 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_92_22
timestamp 1676037725
transform 1 0 3128 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_33
timestamp 1676037725
transform 1 0 4140 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_50
timestamp 1676037725
transform 1 0 5704 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_78
timestamp 1676037725
transform 1 0 8280 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_89
timestamp 1676037725
transform 1 0 9292 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_106
timestamp 1676037725
transform 1 0 10856 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_134
timestamp 1676037725
transform 1 0 13432 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_92_141
timestamp 1676037725
transform 1 0 14076 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_145
timestamp 1676037725
transform 1 0 14444 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_162
timestamp 1676037725
transform 1 0 16008 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_190
timestamp 1676037725
transform 1 0 18584 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_215
timestamp 1676037725
transform 1 0 20884 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_219
timestamp 1676037725
transform 1 0 21252 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_231
timestamp 1676037725
transform 1 0 22356 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_243
timestamp 1676037725
transform 1 0 23460 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1676037725
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1676037725
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1676037725
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1676037725
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1676037725
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1676037725
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1676037725
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1676037725
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1676037725
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1676037725
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1676037725
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1676037725
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1676037725
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1676037725
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1676037725
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1676037725
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1676037725
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1676037725
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1676037725
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1676037725
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1676037725
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1676037725
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1676037725
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1676037725
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1676037725
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1676037725
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1676037725
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_513
timestamp 1676037725
transform 1 0 48300 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_525
timestamp 1676037725
transform 1 0 49404 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_11
timestamp 1676037725
transform 1 0 2116 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_29
timestamp 1676037725
transform 1 0 3772 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_37
timestamp 1676037725
transform 1 0 4508 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_54
timestamp 1676037725
transform 1 0 6072 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_85
timestamp 1676037725
transform 1 0 8924 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_93
timestamp 1676037725
transform 1 0 9660 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_110
timestamp 1676037725
transform 1 0 11224 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_141
timestamp 1676037725
transform 1 0 14076 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_93_149
timestamp 1676037725
transform 1 0 14812 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_166
timestamp 1676037725
transform 1 0 16376 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1676037725
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_197
timestamp 1676037725
transform 1 0 19228 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_201
timestamp 1676037725
transform 1 0 19596 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_93_218
timestamp 1676037725
transform 1 0 21160 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_93_225
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_230
timestamp 1676037725
transform 1 0 22264 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_242
timestamp 1676037725
transform 1 0 23368 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_254
timestamp 1676037725
transform 1 0 24472 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_266
timestamp 1676037725
transform 1 0 25576 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_278
timestamp 1676037725
transform 1 0 26680 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1676037725
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1676037725
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1676037725
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1676037725
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1676037725
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1676037725
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1676037725
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1676037725
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1676037725
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1676037725
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1676037725
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1676037725
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1676037725
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1676037725
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1676037725
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1676037725
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1676037725
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1676037725
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1676037725
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1676037725
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1676037725
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1676037725
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1676037725
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1676037725
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1676037725
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_517
timestamp 1676037725
transform 1 0 48668 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_525
timestamp 1676037725
transform 1 0 49404 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_9
timestamp 1676037725
transform 1 0 1932 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_26
timestamp 1676037725
transform 1 0 3496 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1676037725
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_41
timestamp 1676037725
transform 1 0 4876 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_45
timestamp 1676037725
transform 1 0 5244 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_62
timestamp 1676037725
transform 1 0 6808 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_82
timestamp 1676037725
transform 1 0 8648 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_97
timestamp 1676037725
transform 1 0 10028 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_101
timestamp 1676037725
transform 1 0 10396 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_118
timestamp 1676037725
transform 1 0 11960 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_138
timestamp 1676037725
transform 1 0 13800 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_153
timestamp 1676037725
transform 1 0 15180 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_157
timestamp 1676037725
transform 1 0 15548 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_174
timestamp 1676037725
transform 1 0 17112 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_194
timestamp 1676037725
transform 1 0 18952 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_209
timestamp 1676037725
transform 1 0 20332 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_215
timestamp 1676037725
transform 1 0 20884 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_232
timestamp 1676037725
transform 1 0 22448 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_239
timestamp 1676037725
transform 1 0 23092 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1676037725
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1676037725
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1676037725
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_289
timestamp 1676037725
transform 1 0 27692 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_296
timestamp 1676037725
transform 1 0 28336 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1676037725
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_321
timestamp 1676037725
transform 1 0 30636 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_327
timestamp 1676037725
transform 1 0 31188 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_331
timestamp 1676037725
transform 1 0 31556 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_338
timestamp 1676037725
transform 1 0 32200 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_350
timestamp 1676037725
transform 1 0 33304 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_94_362
timestamp 1676037725
transform 1 0 34408 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1676037725
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_377
timestamp 1676037725
transform 1 0 35788 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_383
timestamp 1676037725
transform 1 0 36340 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_387
timestamp 1676037725
transform 1 0 36708 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_94_394
timestamp 1676037725
transform 1 0 37352 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_402
timestamp 1676037725
transform 1 0 38088 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_94_409
timestamp 1676037725
transform 1 0 38732 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_417
timestamp 1676037725
transform 1 0 39468 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_421
timestamp 1676037725
transform 1 0 39836 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_425
timestamp 1676037725
transform 1 0 40204 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_429
timestamp 1676037725
transform 1 0 40572 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_441
timestamp 1676037725
transform 1 0 41676 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_453
timestamp 1676037725
transform 1 0 42780 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_94_465
timestamp 1676037725
transform 1 0 43884 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_94_472
timestamp 1676037725
transform 1 0 44528 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1676037725
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_489
timestamp 1676037725
transform 1 0 46092 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_495
timestamp 1676037725
transform 1 0 46644 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_500
timestamp 1676037725
transform 1 0 47104 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_94_508
timestamp 1676037725
transform 1 0 47840 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_513
timestamp 1676037725
transform 1 0 48300 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_94_521
timestamp 1676037725
transform 1 0 49036 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1676037725
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1676037725
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_29
timestamp 1676037725
transform 1 0 3772 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_37
timestamp 1676037725
transform 1 0 4508 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1676037725
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_65
timestamp 1676037725
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_82
timestamp 1676037725
transform 1 0 8648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_85
timestamp 1676037725
transform 1 0 8924 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_93
timestamp 1676037725
transform 1 0 9660 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_110
timestamp 1676037725
transform 1 0 11224 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_121
timestamp 1676037725
transform 1 0 12236 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_138
timestamp 1676037725
transform 1 0 13800 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_141
timestamp 1676037725
transform 1 0 14076 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_149
timestamp 1676037725
transform 1 0 14812 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_166
timestamp 1676037725
transform 1 0 16376 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_177
timestamp 1676037725
transform 1 0 17388 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_194
timestamp 1676037725
transform 1 0 18952 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_197
timestamp 1676037725
transform 1 0 19228 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_205
timestamp 1676037725
transform 1 0 19964 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_222
timestamp 1676037725
transform 1 0 21528 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_95_236
timestamp 1676037725
transform 1 0 22816 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_243
timestamp 1676037725
transform 1 0 23460 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_250
timestamp 1676037725
transform 1 0 24104 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_253
timestamp 1676037725
transform 1 0 24380 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_257
timestamp 1676037725
transform 1 0 24748 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_261
timestamp 1676037725
transform 1 0 25116 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_268
timestamp 1676037725
transform 1 0 25760 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_275
timestamp 1676037725
transform 1 0 26404 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1676037725
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_281
timestamp 1676037725
transform 1 0 26956 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_286
timestamp 1676037725
transform 1 0 27416 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_293
timestamp 1676037725
transform 1 0 28060 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_299
timestamp 1676037725
transform 1 0 28612 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_304
timestamp 1676037725
transform 1 0 29072 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_309
timestamp 1676037725
transform 1 0 29532 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_315
timestamp 1676037725
transform 1 0 30084 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_322
timestamp 1676037725
transform 1 0 30728 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1676037725
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1676037725
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_337
timestamp 1676037725
transform 1 0 32108 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_341
timestamp 1676037725
transform 1 0 32476 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_346
timestamp 1676037725
transform 1 0 32936 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_354
timestamp 1676037725
transform 1 0 33672 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_362
timestamp 1676037725
transform 1 0 34408 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_365
timestamp 1676037725
transform 1 0 34684 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_371
timestamp 1676037725
transform 1 0 35236 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_378
timestamp 1676037725
transform 1 0 35880 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1676037725
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1676037725
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_393
timestamp 1676037725
transform 1 0 37260 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_397
timestamp 1676037725
transform 1 0 37628 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_95_402
timestamp 1676037725
transform 1 0 38088 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_95_418
timestamp 1676037725
transform 1 0 39560 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_421
timestamp 1676037725
transform 1 0 39836 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_95_433
timestamp 1676037725
transform 1 0 40940 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_95_445
timestamp 1676037725
transform 1 0 42044 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_449
timestamp 1676037725
transform 1 0 42412 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_471
timestamp 1676037725
transform 1 0 44436 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_475
timestamp 1676037725
transform 1 0 44804 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_477
timestamp 1676037725
transform 1 0 44988 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_483
timestamp 1676037725
transform 1 0 45540 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_491
timestamp 1676037725
transform 1 0 46276 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_499
timestamp 1676037725
transform 1 0 47012 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1676037725
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_505
timestamp 1676037725
transform 1 0 47564 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_511
timestamp 1676037725
transform 1 0 48116 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_95_519
timestamp 1676037725
transform 1 0 48852 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 2300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 48024 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1676037725
transform 1 0 1564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1676037725
transform 1 0 1564 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 1564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1676037725
transform 1 0 1564 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1676037725
transform 1 0 1564 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1676037725
transform 1 0 1564 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1676037725
transform 1 0 1564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 1564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1676037725
transform 1 0 1564 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1676037725
transform 1 0 1564 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1676037725
transform 1 0 1564 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1676037725
transform 1 0 1564 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1676037725
transform 1 0 1564 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1676037725
transform 1 0 1564 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1676037725
transform 1 0 1564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1676037725
transform 1 0 1564 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1676037725
transform 1 0 1564 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1676037725
transform 1 0 1564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1676037725
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1676037725
transform 1 0 1564 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1676037725
transform 1 0 1564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1676037725
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1676037725
transform 1 0 1564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 1564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1676037725
transform 1 0 1564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1676037725
transform 1 0 1564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 21988 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1676037725
transform 1 0 28060 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1676037725
transform 1 0 28704 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1676037725
transform 1 0 29716 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1676037725
transform 1 0 30452 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1676037725
transform 1 0 31096 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1676037725
transform 1 0 31280 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1676037725
transform 1 0 31924 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1676037725
transform 1 0 32568 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1676037725
transform 1 0 33304 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1676037725
transform 1 0 34040 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1676037725
transform 1 0 22816 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1676037725
transform 1 0 34868 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1676037725
transform 1 0 35604 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1676037725
transform 1 0 36248 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1676037725
transform 1 0 36432 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1676037725
transform 1 0 37076 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1676037725
transform 1 0 37720 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1676037725
transform 1 0 38364 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1676037725
transform 1 0 38640 0 -1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1676037725
transform 1 0 40020 0 -1 54400
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1676037725
transform 1 0 40296 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1676037725
transform 1 0 22540 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1676037725
transform 1 0 23184 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1676037725
transform 1 0 23828 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1676037725
transform 1 0 24840 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1676037725
transform 1 0 25484 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1676037725
transform 1 0 26128 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1676037725
transform 1 0 27140 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1676037725
transform 1 0 27784 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1676037725
transform 1 0 32292 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1676037725
transform 1 0 35420 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1676037725
transform 1 0 38640 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1676037725
transform 1 0 42596 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1676037725
transform 1 0 45356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  input68
timestamp 1676037725
transform 1 0 42596 0 -1 54400
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  input69 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 45908 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input70
timestamp 1676037725
transform 1 0 46644 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1676037725
transform 1 0 46736 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1676037725
transform 1 0 47748 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input73
timestamp 1676037725
transform 1 0 48484 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1676037725
transform 1 0 48668 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1676037725
transform 1 0 44160 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1676037725
transform 1 0 45172 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input77 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 48852 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1676037725
transform 1 0 49036 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input79
timestamp 1676037725
transform 1 0 49036 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input80
timestamp 1676037725
transform 1 0 49036 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output81 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 47932 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1676037725
transform 1 0 1656 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1676037725
transform 1 0 1564 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1676037725
transform 1 0 1564 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1676037725
transform 1 0 1564 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1676037725
transform 1 0 1564 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1676037725
transform 1 0 1564 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1676037725
transform 1 0 1564 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1676037725
transform 1 0 1564 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1676037725
transform 1 0 1564 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1676037725
transform 1 0 1564 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1676037725
transform 1 0 1564 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1676037725
transform 1 0 1564 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1676037725
transform 1 0 1564 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1676037725
transform 1 0 1564 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1676037725
transform 1 0 1564 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1676037725
transform 1 0 1564 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1676037725
transform 1 0 1564 0 -1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1676037725
transform 1 0 1564 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1676037725
transform 1 0 1564 0 1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1676037725
transform 1 0 1564 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1676037725
transform 1 0 1564 0 -1 50048
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1676037725
transform 1 0 1564 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1676037725
transform 1 0 1564 0 1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1676037725
transform 1 0 1564 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1676037725
transform 1 0 1564 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1676037725
transform 1 0 1564 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1676037725
transform 1 0 1564 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1676037725
transform 1 0 1564 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1676037725
transform 1 0 1564 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1676037725
transform 1 0 1564 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1676037725
transform 1 0 1564 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1676037725
transform 1 0 2300 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1676037725
transform 1 0 7176 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1676037725
transform 1 0 9384 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1676037725
transform 1 0 9752 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1676037725
transform 1 0 9752 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1676037725
transform 1 0 10488 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1676037725
transform 1 0 11960 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 12604 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 12328 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 12328 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 14536 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 2024 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 14904 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 14904 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 15640 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 17112 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 17756 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 17480 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 17480 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 19688 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 20056 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 20976 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 2024 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 4232 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 4600 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 4600 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 5336 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 6808 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 7452 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 7176 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 6532 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 9108 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 12236 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 14904 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 19412 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 22172 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 25208 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 28796 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 49864 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 49864 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 49864 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 49864 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 49864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 49864 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 49864 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 49864 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 49864 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 49864 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 49864 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 49864 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 49864 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 49864 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 49864 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 49864 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 49864 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 49864 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 49864 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 49864 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 49864 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 49864 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 49864 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 49864 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 49864 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 49864 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 49864 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 49864 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 49864 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 49864 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 49864 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 49864 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 49864 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 49864 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 49864 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 49864 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 49864 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 49864 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 49864 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 49864 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 49864 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 49864 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 49864 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 49864 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 49864 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 49864 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 49864 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 49864 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 49864 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 49864 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 49864 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 49864 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 49864 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 49864 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 49864 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 18124 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14536 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 13340 0 -1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12972 0 -1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14536 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14628 0 1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14076 0 -1 50048
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14352 0 1 50048
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14536 0 -1 51136
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15824 0 1 51136
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17020 0 -1 51136
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 50048
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17112 0 1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17388 0 -1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17112 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17480 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19596 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20056 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 50048
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20884 0 1 50048
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21528 0 1 48960
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23000 0 -1 47872
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22264 0 1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22356 0 -1 46784
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22816 0 -1 45696
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20792 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37536 0 -1 51136
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 -1 44608
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 22356 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21528 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17112 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19504 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19320 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17664 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20148 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20332 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 18860 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 19688 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 20516 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 18952 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20516 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19688 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 17112 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 17388 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16652 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16100 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14536 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14904 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14536 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 17020 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 16928 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 16468 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14536 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14260 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14628 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14352 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12328 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11684 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12052 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12512 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 11960 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11684 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 10212 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10396 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9384 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8464 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6808 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 6808 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 6808 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 8740 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 9752 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 11960 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 12328 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14260 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14536 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15456 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 14536 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 15456 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 15824 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25760 0 1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 20240 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_1.mux_l1_in_1__194
timestamp 1676037725
transform 1 0 20700 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19504 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14076 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17296 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_3.mux_l2_in_0__153
timestamp 1676037725
transform 1 0 13524 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14720 0 1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11776 0 1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_5.mux_l2_in_0__160
timestamp 1676037725
transform 1 0 12696 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8556 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17112 0 -1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_7.mux_l1_in_1__162
timestamp 1676037725
transform 1 0 16468 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 15548 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13340 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10488 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_9.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15916 0 1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_9.mux_l2_in_0__163
timestamp 1676037725
transform 1 0 12328 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_9.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9016 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18032 0 1 51136
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_11.mux_l2_in_0__195
timestamp 1676037725
transform 1 0 14720 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9752 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19504 0 1 51136
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_13.mux_l2_in_0__196
timestamp 1676037725
transform 1 0 16836 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11684 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_15.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19780 0 -1 51136
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_15.mux_l2_in_0__197
timestamp 1676037725
transform 1 0 12328 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_15.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10396 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_17.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19688 0 1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_17.mux_l2_in_0_
timestamp 1676037725
transform 1 0 15732 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_17.mux_l2_in_0__198
timestamp 1676037725
transform 1 0 16836 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9108 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_19.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20332 0 1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_19.mux_l2_in_0__151
timestamp 1676037725
transform 1 0 16836 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_19.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16928 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10948 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18768 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_29.mux_l2_in_0__152
timestamp 1676037725
transform 1 0 18676 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12788 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_31.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23368 0 -1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_31.mux_l2_in_0__154
timestamp 1676037725
transform 1 0 19412 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_31.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13432 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_33.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23000 0 -1 51136
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_33.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_33.mux_l2_in_0__155
timestamp 1676037725
transform 1 0 21988 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12512 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_35.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 50048
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_35.mux_l2_in_0__156
timestamp 1676037725
transform 1 0 20792 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_35.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19596 0 1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13064 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25484 0 1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_45.mux_l2_in_0__157
timestamp 1676037725
transform 1 0 21988 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18860 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14260 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_47.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25484 0 -1 48960
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_47.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21620 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_47.mux_l2_in_0__158
timestamp 1676037725
transform 1 0 21988 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13432 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_49.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25760 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_49.mux_l2_in_0__159
timestamp 1676037725
transform 1 0 21620 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_49.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15364 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_51.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25116 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_51.mux_l2_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_51.mux_l2_in_0__161
timestamp 1676037725
transform 1 0 19136 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13524 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 26772 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27232 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_0.mux_l2_in_1__164
timestamp 1676037725
transform 1 0 18860 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 18032 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 21068 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23184 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23368 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21252 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_2.mux_l2_in_1__170
timestamp 1676037725
transform 1 0 13248 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12052 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 18400 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17756 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22724 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 22724 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 20056 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_4.mux_l2_in_1__181
timestamp 1676037725
transform 1 0 12236 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 11868 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 17204 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17204 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24472 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_6.mux_l2_in_1__188
timestamp 1676037725
transform 1 0 16192 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14996 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17480 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24288 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 22172 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 14904 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_8.mux_l2_in_1__189
timestamp 1676037725
transform 1 0 14260 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 16928 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18124 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 23092 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23092 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_10.mux_l2_in_1__165
timestamp 1676037725
transform 1 0 15180 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 13984 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 15548 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17664 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 17756 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_12.mux_l1_in_1__166
timestamp 1676037725
transform 1 0 14260 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 14260 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16928 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16100 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18492 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_14.mux_l1_in_1__167
timestamp 1676037725
transform 1 0 10764 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10396 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14168 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17848 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_16.mux_l1_in_1__168
timestamp 1676037725
transform 1 0 11408 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10212 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14352 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 17480 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20332 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l1_in_1_
timestamp 1676037725
transform 1 0 12972 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_18.mux_l1_in_1__169
timestamp 1676037725
transform 1 0 14352 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16928 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 15088 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15548 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 16836 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_20.mux_l2_in_0__171
timestamp 1676037725
transform 1 0 16284 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14904 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 14260 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14812 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_22.mux_l2_in_0__172
timestamp 1676037725
transform 1 0 13800 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14260 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 15456 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_24.mux_l2_in_0__173
timestamp 1676037725
transform 1 0 16008 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14168 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14260 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12328 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12420 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_26.mux_l2_in_0__174
timestamp 1676037725
transform 1 0 12328 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 12788 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 11684 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_28.mux_l2_in_0__175
timestamp 1676037725
transform 1 0 11776 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9752 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_30.mux_l2_in_0__176
timestamp 1676037725
transform 1 0 7176 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11040 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12512 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_32.mux_l2_in_0__177
timestamp 1676037725
transform 1 0 12144 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11684 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11224 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12144 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_34.mux_l2_in_0__178
timestamp 1676037725
transform 1 0 11684 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 13064 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10304 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_36.mux_l2_in_0__179
timestamp 1676037725
transform 1 0 10856 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 10396 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9660 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_38.mux_l1_in_0_
timestamp 1676037725
transform 1 0 8740 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_38.mux_l2_in_0_
timestamp 1676037725
transform 1 0 9108 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_38.mux_l2_in_0__180
timestamp 1676037725
transform 1 0 7084 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 7912 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 8004 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_40.mux_l2_in_0__182
timestamp 1676037725
transform 1 0 8372 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 7820 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 8004 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_42.mux_l1_in_0_
timestamp 1676037725
transform 1 0 13156 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_42.mux_l2_in_0__183
timestamp 1676037725
transform 1 0 12328 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_42.mux_l2_in_0_
timestamp 1676037725
transform 1 0 11224 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 9568 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19228 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_44.mux_l1_in_1__184
timestamp 1676037725
transform 1 0 11592 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 12972 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10948 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20976 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_46.mux_l1_in_1__185
timestamp 1676037725
transform 1 0 11684 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10396 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14260 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11132 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_48.mux_l1_in_1__186
timestamp 1676037725
transform 1 0 11684 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l1_in_1_
timestamp 1676037725
transform 1 0 11776 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14352 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 11684 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 19504 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l1_in_1_
timestamp 1676037725
transform 1 0 10580 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_50.mux_l1_in_1__187
timestamp 1676037725
transform 1 0 18216 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 14812 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 10948 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1676037725
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1676037725
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1676037725
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1676037725
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1676037725
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1676037725
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1676037725
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1676037725
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1676037725
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1676037725
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1676037725
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1676037725
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1676037725
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1676037725
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1676037725
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1676037725
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1676037725
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1676037725
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1676037725
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1676037725
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1676037725
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1676037725
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1676037725
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1676037725
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1676037725
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1676037725
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1676037725
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1676037725
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1676037725
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1676037725
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1676037725
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1676037725
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1676037725
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1676037725
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1676037725
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1676037725
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1676037725
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1676037725
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1676037725
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1676037725
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1676037725
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1676037725
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1676037725
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1676037725
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1676037725
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1676037725
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1676037725
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1676037725
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1676037725
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1676037725
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1676037725
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1676037725
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1676037725
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1676037725
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1676037725
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1676037725
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1676037725
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1676037725
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1676037725
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1676037725
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1676037725
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1676037725
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1676037725
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1676037725
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1676037725
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1676037725
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1676037725
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1676037725
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1676037725
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1676037725
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1676037725
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1676037725
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1676037725
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1676037725
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1676037725
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1676037725
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1676037725
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1676037725
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1676037725
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1676037725
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1676037725
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1676037725
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1676037725
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1676037725
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1676037725
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1676037725
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1676037725
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1676037725
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1676037725
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1676037725
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1676037725
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1676037725
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1676037725
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1676037725
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1676037725
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1676037725
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1676037725
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1676037725
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1676037725
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1676037725
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1676037725
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1676037725
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1676037725
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1676037725
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1676037725
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1676037725
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1676037725
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1676037725
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1676037725
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1676037725
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1676037725
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1676037725
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1676037725
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1676037725
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1676037725
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1676037725
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1676037725
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1676037725
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1676037725
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1676037725
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1676037725
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1676037725
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1676037725
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1676037725
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1676037725
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1676037725
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1676037725
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1676037725
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1676037725
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1676037725
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1676037725
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1676037725
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1676037725
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1676037725
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1676037725
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1676037725
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1676037725
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1676037725
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1676037725
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1676037725
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1676037725
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1676037725
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1676037725
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1676037725
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1676037725
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1676037725
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1676037725
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1676037725
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1676037725
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1676037725
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1676037725
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1676037725
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1676037725
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1676037725
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1676037725
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1676037725
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1676037725
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1676037725
transform 1 0 29440 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1676037725
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1676037725
transform 1 0 34592 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1676037725
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1676037725
transform 1 0 39744 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1676037725
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1676037725
transform 1 0 44896 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1676037725
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  wire1
timestamp 1676037725
transform 1 0 46644 0 -1 3264
box -38 -48 406 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 49238 56200 49294 57000 0 FreeSans 224 90 0 0 ccff_head_1
port 3 nsew signal input
flabel metal3 s 50200 45840 51000 45960 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 1582 56200 1638 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 chanx_left_in[20]
port 18 nsew signal input
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 chanx_left_in[21]
port 19 nsew signal input
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_in[22]
port 20 nsew signal input
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 chanx_left_in[23]
port 21 nsew signal input
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 chanx_left_in[24]
port 22 nsew signal input
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 chanx_left_in[25]
port 23 nsew signal input
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 chanx_left_in[26]
port 24 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_in[27]
port 25 nsew signal input
flabel metal3 s 0 25984 800 26104 0 FreeSans 480 0 0 0 chanx_left_in[28]
port 26 nsew signal input
flabel metal3 s 0 26800 800 26920 0 FreeSans 480 0 0 0 chanx_left_in[29]
port 27 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 28 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 29 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 30 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 31 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 32 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 33 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 34 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 35 nsew signal input
flabel metal3 s 0 27616 800 27736 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 36 nsew signal tristate
flabel metal3 s 0 35776 800 35896 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 37 nsew signal tristate
flabel metal3 s 0 36592 800 36712 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 38 nsew signal tristate
flabel metal3 s 0 37408 800 37528 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 39 nsew signal tristate
flabel metal3 s 0 38224 800 38344 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 40 nsew signal tristate
flabel metal3 s 0 39040 800 39160 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 41 nsew signal tristate
flabel metal3 s 0 39856 800 39976 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 42 nsew signal tristate
flabel metal3 s 0 40672 800 40792 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 43 nsew signal tristate
flabel metal3 s 0 41488 800 41608 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 44 nsew signal tristate
flabel metal3 s 0 42304 800 42424 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 45 nsew signal tristate
flabel metal3 s 0 43120 800 43240 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 46 nsew signal tristate
flabel metal3 s 0 28432 800 28552 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 47 nsew signal tristate
flabel metal3 s 0 43936 800 44056 0 FreeSans 480 0 0 0 chanx_left_out[20]
port 48 nsew signal tristate
flabel metal3 s 0 44752 800 44872 0 FreeSans 480 0 0 0 chanx_left_out[21]
port 49 nsew signal tristate
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 chanx_left_out[22]
port 50 nsew signal tristate
flabel metal3 s 0 46384 800 46504 0 FreeSans 480 0 0 0 chanx_left_out[23]
port 51 nsew signal tristate
flabel metal3 s 0 47200 800 47320 0 FreeSans 480 0 0 0 chanx_left_out[24]
port 52 nsew signal tristate
flabel metal3 s 0 48016 800 48136 0 FreeSans 480 0 0 0 chanx_left_out[25]
port 53 nsew signal tristate
flabel metal3 s 0 48832 800 48952 0 FreeSans 480 0 0 0 chanx_left_out[26]
port 54 nsew signal tristate
flabel metal3 s 0 49648 800 49768 0 FreeSans 480 0 0 0 chanx_left_out[27]
port 55 nsew signal tristate
flabel metal3 s 0 50464 800 50584 0 FreeSans 480 0 0 0 chanx_left_out[28]
port 56 nsew signal tristate
flabel metal3 s 0 51280 800 51400 0 FreeSans 480 0 0 0 chanx_left_out[29]
port 57 nsew signal tristate
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 30064 800 30184 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 30880 800 31000 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 31696 800 31816 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 32512 800 32632 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 34144 800 34264 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 34960 800 35080 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal2 s 21546 56200 21602 57000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 66 nsew signal input
flabel metal2 s 27986 56200 28042 57000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 67 nsew signal input
flabel metal2 s 28630 56200 28686 57000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 68 nsew signal input
flabel metal2 s 29274 56200 29330 57000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 69 nsew signal input
flabel metal2 s 29918 56200 29974 57000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 70 nsew signal input
flabel metal2 s 30562 56200 30618 57000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 71 nsew signal input
flabel metal2 s 31206 56200 31262 57000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 72 nsew signal input
flabel metal2 s 31850 56200 31906 57000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 73 nsew signal input
flabel metal2 s 32494 56200 32550 57000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 74 nsew signal input
flabel metal2 s 33138 56200 33194 57000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 75 nsew signal input
flabel metal2 s 33782 56200 33838 57000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 76 nsew signal input
flabel metal2 s 22190 56200 22246 57000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 77 nsew signal input
flabel metal2 s 34426 56200 34482 57000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 78 nsew signal input
flabel metal2 s 35070 56200 35126 57000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 79 nsew signal input
flabel metal2 s 35714 56200 35770 57000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 80 nsew signal input
flabel metal2 s 36358 56200 36414 57000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 81 nsew signal input
flabel metal2 s 37002 56200 37058 57000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 82 nsew signal input
flabel metal2 s 37646 56200 37702 57000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 83 nsew signal input
flabel metal2 s 38290 56200 38346 57000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 84 nsew signal input
flabel metal2 s 38934 56200 38990 57000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 85 nsew signal input
flabel metal2 s 39578 56200 39634 57000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 86 nsew signal input
flabel metal2 s 40222 56200 40278 57000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 87 nsew signal input
flabel metal2 s 22834 56200 22890 57000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 88 nsew signal input
flabel metal2 s 23478 56200 23534 57000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 89 nsew signal input
flabel metal2 s 24122 56200 24178 57000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 90 nsew signal input
flabel metal2 s 24766 56200 24822 57000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 91 nsew signal input
flabel metal2 s 25410 56200 25466 57000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 92 nsew signal input
flabel metal2 s 26054 56200 26110 57000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 93 nsew signal input
flabel metal2 s 26698 56200 26754 57000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 94 nsew signal input
flabel metal2 s 27342 56200 27398 57000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 95 nsew signal input
flabel metal2 s 2226 56200 2282 57000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 96 nsew signal tristate
flabel metal2 s 8666 56200 8722 57000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 97 nsew signal tristate
flabel metal2 s 9310 56200 9366 57000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 98 nsew signal tristate
flabel metal2 s 9954 56200 10010 57000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 99 nsew signal tristate
flabel metal2 s 10598 56200 10654 57000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 100 nsew signal tristate
flabel metal2 s 11242 56200 11298 57000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 101 nsew signal tristate
flabel metal2 s 11886 56200 11942 57000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 102 nsew signal tristate
flabel metal2 s 12530 56200 12586 57000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 103 nsew signal tristate
flabel metal2 s 13174 56200 13230 57000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 104 nsew signal tristate
flabel metal2 s 13818 56200 13874 57000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 105 nsew signal tristate
flabel metal2 s 14462 56200 14518 57000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 106 nsew signal tristate
flabel metal2 s 2870 56200 2926 57000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 107 nsew signal tristate
flabel metal2 s 15106 56200 15162 57000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 108 nsew signal tristate
flabel metal2 s 15750 56200 15806 57000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 109 nsew signal tristate
flabel metal2 s 16394 56200 16450 57000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 110 nsew signal tristate
flabel metal2 s 17038 56200 17094 57000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 111 nsew signal tristate
flabel metal2 s 17682 56200 17738 57000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 112 nsew signal tristate
flabel metal2 s 18326 56200 18382 57000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 113 nsew signal tristate
flabel metal2 s 18970 56200 19026 57000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 114 nsew signal tristate
flabel metal2 s 19614 56200 19670 57000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 115 nsew signal tristate
flabel metal2 s 20258 56200 20314 57000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 116 nsew signal tristate
flabel metal2 s 20902 56200 20958 57000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 117 nsew signal tristate
flabel metal2 s 3514 56200 3570 57000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 118 nsew signal tristate
flabel metal2 s 4158 56200 4214 57000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 119 nsew signal tristate
flabel metal2 s 4802 56200 4858 57000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 120 nsew signal tristate
flabel metal2 s 5446 56200 5502 57000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 121 nsew signal tristate
flabel metal2 s 6090 56200 6146 57000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 122 nsew signal tristate
flabel metal2 s 6734 56200 6790 57000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 123 nsew signal tristate
flabel metal2 s 7378 56200 7434 57000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 124 nsew signal tristate
flabel metal2 s 8022 56200 8078 57000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 125 nsew signal tristate
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 126 nsew signal tristate
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 127 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 128 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 129 nsew signal tristate
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 130 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 131 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 132 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 133 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 134 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 135 nsew signal tristate
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 136 nsew signal tristate
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 137 nsew signal tristate
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 isol_n
port 138 nsew signal input
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 prog_clk
port 139 nsew signal input
flabel metal2 s 42154 56200 42210 57000 0 FreeSans 224 90 0 0 prog_reset_top_in
port 140 nsew signal input
flabel metal2 s 42798 56200 42854 57000 0 FreeSans 224 90 0 0 reset_top_in
port 141 nsew signal input
flabel metal2 s 43442 56200 43498 57000 0 FreeSans 224 90 0 0 test_enable_top_in
port 142 nsew signal input
flabel metal2 s 45374 56200 45430 57000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 143 nsew signal input
flabel metal2 s 46018 56200 46074 57000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 144 nsew signal input
flabel metal2 s 46662 56200 46718 57000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 145 nsew signal input
flabel metal2 s 47306 56200 47362 57000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 146 nsew signal input
flabel metal2 s 47950 56200 48006 57000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 147 nsew signal input
flabel metal2 s 48594 56200 48650 57000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 148 nsew signal input
flabel metal2 s 44086 56200 44142 57000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 149 nsew signal input
flabel metal2 s 44730 56200 44786 57000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 150 nsew signal input
flabel metal3 s 50200 48016 51000 48136 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 151 nsew signal input
flabel metal3 s 50200 50192 51000 50312 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 152 nsew signal input
flabel metal3 s 50200 52368 51000 52488 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 153 nsew signal input
flabel metal3 s 50200 54544 51000 54664 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 154 nsew signal input
flabel metal3 s 0 52096 800 52216 0 FreeSans 480 0 0 0 top_width_0_height_0_subtile_0__pin_inpad_0_
port 155 nsew signal tristate
flabel metal3 s 0 52912 800 53032 0 FreeSans 480 0 0 0 top_width_0_height_0_subtile_1__pin_inpad_0_
port 156 nsew signal tristate
flabel metal3 s 0 53728 800 53848 0 FreeSans 480 0 0 0 top_width_0_height_0_subtile_2__pin_inpad_0_
port 157 nsew signal tristate
flabel metal3 s 0 54544 800 54664 0 FreeSans 480 0 0 0 top_width_0_height_0_subtile_3__pin_inpad_0_
port 158 nsew signal tristate
rlabel metal1 25484 54400 25484 54400 0 VGND
rlabel metal1 25484 53856 25484 53856 0 VPWR
rlabel metal1 19780 12886 19780 12886 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal2 19182 16932 19182 16932 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal2 18630 17340 18630 17340 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 15088 27302 15088 27302 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 18577 40698 18577 40698 0 cbx_8__0_.cbx_8__0_.ccff_head
rlabel metal1 11408 29818 11408 29818 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
rlabel metal2 18906 40239 18906 40239 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
rlabel metal1 9430 31688 9430 31688 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
rlabel metal1 9982 29512 9982 29512 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
rlabel metal1 9476 29070 9476 29070 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
rlabel metal1 10948 31382 10948 31382 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
rlabel metal1 7958 28662 7958 28662 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
rlabel metal1 8418 30804 8418 30804 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
rlabel metal2 13570 30702 13570 30702 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
rlabel metal1 13202 34102 13202 34102 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
rlabel metal1 11132 30634 11132 30634 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
rlabel metal2 12650 29886 12650 29886 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
rlabel metal1 13662 31382 13662 31382 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
rlabel metal2 13938 38080 13938 38080 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
rlabel metal1 9660 38386 9660 38386 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
rlabel metal1 8878 36890 8878 36890 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12098 28050 12098 28050 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 13984 26758 13984 26758 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 8418 37264 8418 37264 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8648 35666 8648 35666 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9706 35802 9706 35802 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10902 28526 10902 28526 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 9844 32878 9844 32878 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9476 32878 9476 32878 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10304 28730 10304 28730 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 10304 29274 10304 29274 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10764 27030 10764 27030 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 5934 36108 5934 36108 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 9798 29546 9798 29546 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 11960 20910 11960 20910 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 5842 35802 5842 35802 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6946 35122 6946 35122 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7682 35054 7682 35054 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 7958 28594 7958 28594 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7820 32810 7820 32810 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 7406 32878 7406 32878 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 7866 29750 7866 29750 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 7958 30702 7958 30702 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 9890 29631 9890 29631 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 6348 35666 6348 35666 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12880 28934 12880 28934 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 15502 20910 15502 20910 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 6486 35802 6486 35802 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7590 33558 7590 33558 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7912 33626 7912 33626 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 11822 28526 11822 28526 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 9844 32402 9844 32402 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 10442 32912 10442 32912 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 12282 28730 12282 28730 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 15962 39066 15962 39066 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 12880 28118 12880 28118 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 6394 37128 6394 37128 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9384 38522 9384 38522 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 13708 27438 13708 27438 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 5290 38726 5290 38726 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8142 36210 8142 36210 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 7866 35632 7866 35632 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9522 32538 9522 32538 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 5658 38046 5658 38046 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6716 36346 6716 36346 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 8878 35360 8878 35360 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 13846 38454 13846 38454 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 5198 37128 5198 37128 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 21390 11322 21390 11322 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 20470 5678 20470 5678 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 24656 6358 24656 6358 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 29279 14042 29279 14042 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 24702 17068 24702 17068 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 18170 6358 18170 6358 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 21252 12682 21252 12682 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 27255 14246 27255 14246 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 26450 20978 26450 20978 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 18032 13838 18032 13838 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal1 20102 14042 20102 14042 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel via1 24495 15130 24495 15130 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 20470 17170 20470 17170 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal1 18078 8942 18078 8942 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 24449 16558 24449 16558 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 2254 1588 2254 1588 0 ccff_head
rlabel metal1 48760 53618 48760 53618 0 ccff_head_1
rlabel metal3 49734 45900 49734 45900 0 ccff_tail
rlabel metal1 1886 52530 1886 52530 0 ccff_tail_0
rlabel metal3 820 3196 820 3196 0 chanx_left_in[0]
rlabel metal3 820 11356 820 11356 0 chanx_left_in[10]
rlabel metal3 820 12172 820 12172 0 chanx_left_in[11]
rlabel metal3 820 12988 820 12988 0 chanx_left_in[12]
rlabel metal3 820 13804 820 13804 0 chanx_left_in[13]
rlabel metal3 820 14620 820 14620 0 chanx_left_in[14]
rlabel metal3 820 15436 820 15436 0 chanx_left_in[15]
rlabel metal3 820 16252 820 16252 0 chanx_left_in[16]
rlabel metal3 820 17068 820 17068 0 chanx_left_in[17]
rlabel metal3 1234 17884 1234 17884 0 chanx_left_in[18]
rlabel metal3 820 18700 820 18700 0 chanx_left_in[19]
rlabel metal3 820 4012 820 4012 0 chanx_left_in[1]
rlabel metal3 820 19516 820 19516 0 chanx_left_in[20]
rlabel metal3 820 20332 820 20332 0 chanx_left_in[21]
rlabel metal3 820 21148 820 21148 0 chanx_left_in[22]
rlabel metal3 820 21964 820 21964 0 chanx_left_in[23]
rlabel metal3 820 22780 820 22780 0 chanx_left_in[24]
rlabel metal3 820 23596 820 23596 0 chanx_left_in[25]
rlabel metal3 820 24412 820 24412 0 chanx_left_in[26]
rlabel metal3 820 25228 820 25228 0 chanx_left_in[27]
rlabel metal3 1142 26044 1142 26044 0 chanx_left_in[28]
rlabel metal3 820 26860 820 26860 0 chanx_left_in[29]
rlabel metal3 820 4828 820 4828 0 chanx_left_in[2]
rlabel metal3 820 5644 820 5644 0 chanx_left_in[3]
rlabel metal3 820 6460 820 6460 0 chanx_left_in[4]
rlabel metal3 820 7276 820 7276 0 chanx_left_in[5]
rlabel metal3 1234 8092 1234 8092 0 chanx_left_in[6]
rlabel metal3 820 8908 820 8908 0 chanx_left_in[7]
rlabel metal3 820 9724 820 9724 0 chanx_left_in[8]
rlabel metal3 820 10540 820 10540 0 chanx_left_in[9]
rlabel metal3 1004 27676 1004 27676 0 chanx_left_out[0]
rlabel metal2 2806 35955 2806 35955 0 chanx_left_out[10]
rlabel metal3 1004 36652 1004 36652 0 chanx_left_out[11]
rlabel metal3 1004 37468 1004 37468 0 chanx_left_out[12]
rlabel metal3 1004 38284 1004 38284 0 chanx_left_out[13]
rlabel metal3 1004 39100 1004 39100 0 chanx_left_out[14]
rlabel metal3 1372 39916 1372 39916 0 chanx_left_out[15]
rlabel metal3 1004 40732 1004 40732 0 chanx_left_out[16]
rlabel metal3 1004 41548 1004 41548 0 chanx_left_out[17]
rlabel metal3 1004 42364 1004 42364 0 chanx_left_out[18]
rlabel metal3 1004 43180 1004 43180 0 chanx_left_out[19]
rlabel metal3 1004 28492 1004 28492 0 chanx_left_out[1]
rlabel metal3 1372 43996 1372 43996 0 chanx_left_out[20]
rlabel metal3 1004 44812 1004 44812 0 chanx_left_out[21]
rlabel metal3 1004 45628 1004 45628 0 chanx_left_out[22]
rlabel metal3 1004 46444 1004 46444 0 chanx_left_out[23]
rlabel metal3 1004 47260 1004 47260 0 chanx_left_out[24]
rlabel metal3 1004 48076 1004 48076 0 chanx_left_out[25]
rlabel metal3 1004 48892 1004 48892 0 chanx_left_out[26]
rlabel metal3 1004 49708 1004 49708 0 chanx_left_out[27]
rlabel metal3 1004 50524 1004 50524 0 chanx_left_out[28]
rlabel metal3 1004 51340 1004 51340 0 chanx_left_out[29]
rlabel metal3 1004 29308 1004 29308 0 chanx_left_out[2]
rlabel metal3 1004 30124 1004 30124 0 chanx_left_out[3]
rlabel metal3 1004 30940 1004 30940 0 chanx_left_out[4]
rlabel metal3 1004 31756 1004 31756 0 chanx_left_out[5]
rlabel metal3 1004 32572 1004 32572 0 chanx_left_out[6]
rlabel metal3 1004 33388 1004 33388 0 chanx_left_out[7]
rlabel metal3 1372 34204 1372 34204 0 chanx_left_out[8]
rlabel metal3 1004 35020 1004 35020 0 chanx_left_out[9]
rlabel metal2 21574 54648 21574 54648 0 chany_top_in[0]
rlabel metal1 28060 53550 28060 53550 0 chany_top_in[10]
rlabel metal1 28750 54230 28750 54230 0 chany_top_in[11]
rlabel metal1 29578 54230 29578 54230 0 chany_top_in[12]
rlabel metal1 30544 54162 30544 54162 0 chany_top_in[13]
rlabel metal1 31326 54196 31326 54196 0 chany_top_in[14]
rlabel metal1 31372 53550 31372 53550 0 chany_top_in[15]
rlabel metal1 32016 53550 32016 53550 0 chany_top_in[16]
rlabel metal1 32614 54230 32614 54230 0 chany_top_in[17]
rlabel metal1 33304 54230 33304 54230 0 chany_top_in[18]
rlabel metal1 33994 54230 33994 54230 0 chany_top_in[19]
rlabel metal1 22632 53550 22632 53550 0 chany_top_in[1]
rlabel metal1 34730 54230 34730 54230 0 chany_top_in[20]
rlabel metal1 35466 54162 35466 54162 0 chany_top_in[21]
rlabel metal1 36202 54162 36202 54162 0 chany_top_in[22]
rlabel metal1 36524 53550 36524 53550 0 chany_top_in[23]
rlabel metal1 37168 53550 37168 53550 0 chany_top_in[24]
rlabel metal1 37766 54230 37766 54230 0 chany_top_in[25]
rlabel metal1 38410 53550 38410 53550 0 chany_top_in[26]
rlabel metal1 38824 54162 38824 54162 0 chany_top_in[27]
rlabel metal1 39836 54162 39836 54162 0 chany_top_in[28]
rlabel metal1 40388 53550 40388 53550 0 chany_top_in[29]
rlabel metal1 22816 54162 22816 54162 0 chany_top_in[2]
rlabel metal1 23460 54162 23460 54162 0 chany_top_in[3]
rlabel metal1 24104 54162 24104 54162 0 chany_top_in[4]
rlabel metal1 24978 54162 24978 54162 0 chany_top_in[5]
rlabel metal1 25576 54162 25576 54162 0 chany_top_in[6]
rlabel metal1 26312 54162 26312 54162 0 chany_top_in[7]
rlabel metal1 27048 54162 27048 54162 0 chany_top_in[8]
rlabel metal1 27830 54162 27830 54162 0 chany_top_in[9]
rlabel metal1 2530 53006 2530 53006 0 chany_top_out[0]
rlabel metal1 8556 54230 8556 54230 0 chany_top_out[10]
rlabel metal1 9614 52530 9614 52530 0 chany_top_out[11]
rlabel metal2 9982 55711 9982 55711 0 chany_top_out[12]
rlabel metal1 10672 54230 10672 54230 0 chany_top_out[13]
rlabel metal2 11270 54920 11270 54920 0 chany_top_out[14]
rlabel metal1 12190 52530 12190 52530 0 chany_top_out[15]
rlabel metal2 12558 55711 12558 55711 0 chany_top_out[16]
rlabel metal2 13202 55711 13202 55711 0 chany_top_out[17]
rlabel metal1 13708 54230 13708 54230 0 chany_top_out[18]
rlabel metal1 14766 52530 14766 52530 0 chany_top_out[19]
rlabel metal2 2898 54920 2898 54920 0 chany_top_out[1]
rlabel metal1 15134 52972 15134 52972 0 chany_top_out[20]
rlabel metal1 15824 54230 15824 54230 0 chany_top_out[21]
rlabel metal2 16422 54920 16422 54920 0 chany_top_out[22]
rlabel metal1 17342 52530 17342 52530 0 chany_top_out[23]
rlabel metal1 17986 53006 17986 53006 0 chany_top_out[24]
rlabel metal2 18354 54920 18354 54920 0 chany_top_out[25]
rlabel metal1 18860 54230 18860 54230 0 chany_top_out[26]
rlabel metal1 19918 53006 19918 53006 0 chany_top_out[27]
rlabel metal1 20424 54094 20424 54094 0 chany_top_out[28]
rlabel metal1 21206 53618 21206 53618 0 chany_top_out[29]
rlabel metal1 3404 54230 3404 54230 0 chany_top_out[2]
rlabel metal1 4462 52530 4462 52530 0 chany_top_out[3]
rlabel metal1 4968 53006 4968 53006 0 chany_top_out[4]
rlabel metal2 5474 55158 5474 55158 0 chany_top_out[5]
rlabel metal2 6118 54920 6118 54920 0 chany_top_out[6]
rlabel metal2 6762 54376 6762 54376 0 chany_top_out[7]
rlabel metal2 7406 55711 7406 55711 0 chany_top_out[8]
rlabel metal2 8050 55711 8050 55711 0 chany_top_out[9]
rlabel metal2 11914 30090 11914 30090 0 clknet_0_prog_clk
rlabel metal2 9062 33762 9062 33762 0 clknet_4_0_0_prog_clk
rlabel metal2 14122 49300 14122 49300 0 clknet_4_10_0_prog_clk
rlabel metal2 37582 50286 37582 50286 0 clknet_4_11_0_prog_clk
rlabel metal1 18860 36754 18860 36754 0 clknet_4_12_0_prog_clk
rlabel metal2 24702 20944 24702 20944 0 clknet_4_13_0_prog_clk
rlabel metal1 14582 41174 14582 41174 0 clknet_4_14_0_prog_clk
rlabel metal2 19734 40290 19734 40290 0 clknet_4_15_0_prog_clk
rlabel metal1 14490 37298 14490 37298 0 clknet_4_1_0_prog_clk
rlabel metal2 8510 39202 8510 39202 0 clknet_4_2_0_prog_clk
rlabel metal1 8970 41106 8970 41106 0 clknet_4_3_0_prog_clk
rlabel metal1 10028 7922 10028 7922 0 clknet_4_4_0_prog_clk
rlabel metal1 10212 30770 10212 30770 0 clknet_4_5_0_prog_clk
rlabel metal1 14536 32402 14536 32402 0 clknet_4_6_0_prog_clk
rlabel metal1 19366 32266 19366 32266 0 clknet_4_7_0_prog_clk
rlabel metal1 15364 42670 15364 42670 0 clknet_4_8_0_prog_clk
rlabel metal1 20240 46002 20240 46002 0 clknet_4_9_0_prog_clk
rlabel metal2 5566 1622 5566 1622 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 8878 1622 8878 1622 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 12190 1622 12190 1622 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 15502 1622 15502 1622 0 gfpga_pad_io_soc_dir[3]
rlabel metal2 32062 1588 32062 1588 0 gfpga_pad_io_soc_in[0]
rlabel metal2 35374 1588 35374 1588 0 gfpga_pad_io_soc_in[1]
rlabel metal2 38686 1588 38686 1588 0 gfpga_pad_io_soc_in[2]
rlabel metal2 41998 1588 41998 1588 0 gfpga_pad_io_soc_in[3]
rlabel metal2 18814 1622 18814 1622 0 gfpga_pad_io_soc_out[0]
rlabel metal2 22126 1622 22126 1622 0 gfpga_pad_io_soc_out[1]
rlabel metal2 25438 1622 25438 1622 0 gfpga_pad_io_soc_out[2]
rlabel metal2 28750 1860 28750 1860 0 gfpga_pad_io_soc_out[3]
rlabel metal2 45310 1554 45310 1554 0 isol_n
rlabel metal1 6532 2278 6532 2278 0 net1
rlabel metal1 1932 16694 1932 16694 0 net10
rlabel metal2 3910 46818 3910 46818 0 net100
rlabel metal2 3450 47124 3450 47124 0 net101
rlabel metal2 4646 47668 4646 47668 0 net102
rlabel metal2 3358 48518 3358 48518 0 net103
rlabel metal1 3496 51374 3496 51374 0 net104
rlabel metal1 1794 29648 1794 29648 0 net105
rlabel metal2 1794 30022 1794 30022 0 net106
rlabel metal1 3680 31314 3680 31314 0 net107
rlabel metal2 5658 32538 5658 32538 0 net108
rlabel metal2 4738 34714 4738 34714 0 net109
rlabel via2 1886 17085 1886 17085 0 net11
rlabel metal2 6118 36108 6118 36108 0 net110
rlabel metal1 1794 34612 1794 34612 0 net111
rlabel metal2 4002 37468 4002 37468 0 net112
rlabel metal1 2622 53074 2622 53074 0 net113
rlabel metal1 7590 54162 7590 54162 0 net114
rlabel metal2 9706 52292 9706 52292 0 net115
rlabel metal1 10166 52122 10166 52122 0 net116
rlabel metal2 10902 52870 10902 52870 0 net117
rlabel metal1 11224 53550 11224 53550 0 net118
rlabel metal1 11914 52462 11914 52462 0 net119
rlabel metal1 5152 18394 5152 18394 0 net12
rlabel metal1 12420 53074 12420 53074 0 net120
rlabel metal1 12282 51034 12282 51034 0 net121
rlabel metal1 12696 51034 12696 51034 0 net122
rlabel metal1 14076 51578 14076 51578 0 net123
rlabel metal1 3496 53550 3496 53550 0 net124
rlabel metal2 15594 52598 15594 52598 0 net125
rlabel metal1 13800 54162 13800 54162 0 net126
rlabel metal1 14766 53550 14766 53550 0 net127
rlabel metal1 17020 52462 17020 52462 0 net128
rlabel metal1 17710 52122 17710 52122 0 net129
rlabel metal1 5014 18938 5014 18938 0 net13
rlabel metal1 19274 53550 19274 53550 0 net130
rlabel metal1 18400 52122 18400 52122 0 net131
rlabel metal1 20056 48858 20056 48858 0 net132
rlabel metal1 19918 54162 19918 54162 0 net133
rlabel metal2 21022 53108 21022 53108 0 net134
rlabel metal1 2300 54162 2300 54162 0 net135
rlabel metal1 4048 44438 4048 44438 0 net136
rlabel metal1 5290 53074 5290 53074 0 net137
rlabel metal1 4876 54162 4876 54162 0 net138
rlabel metal1 5520 53550 5520 53550 0 net139
rlabel metal1 7130 4046 7130 4046 0 net14
rlabel metal2 9246 52020 9246 52020 0 net140
rlabel metal1 8372 53074 8372 53074 0 net141
rlabel metal1 7544 51578 7544 51578 0 net142
rlabel metal1 6854 2414 6854 2414 0 net143
rlabel metal1 9338 2380 9338 2380 0 net144
rlabel metal1 13386 2414 13386 2414 0 net145
rlabel metal2 18354 3978 18354 3978 0 net146
rlabel metal1 18998 8874 18998 8874 0 net147
rlabel metal1 21666 6698 21666 6698 0 net148
rlabel metal1 23184 6698 23184 6698 0 net149
rlabel metal2 1886 20145 1886 20145 0 net15
rlabel metal2 28842 4590 28842 4590 0 net150
rlabel metal1 17204 44846 17204 44846 0 net151
rlabel metal1 19044 43962 19044 43962 0 net152
rlabel metal1 13570 46138 13570 46138 0 net153
rlabel metal1 18952 44846 18952 44846 0 net154
rlabel metal2 20746 48042 20746 48042 0 net155
rlabel metal1 20516 48110 20516 48110 0 net156
rlabel metal1 20746 45458 20746 45458 0 net157
rlabel metal2 22034 44540 22034 44540 0 net158
rlabel metal2 21850 43588 21850 43588 0 net159
rlabel metal1 4508 20434 4508 20434 0 net16
rlabel metal2 12926 46750 12926 46750 0 net160
rlabel metal1 19596 42194 19596 42194 0 net161
rlabel metal1 16008 45526 16008 45526 0 net162
rlabel metal2 13386 48314 13386 48314 0 net163
rlabel metal1 18538 41582 18538 41582 0 net164
rlabel metal1 14904 30226 14904 30226 0 net165
rlabel metal1 14582 29614 14582 29614 0 net166
rlabel metal2 10810 24378 10810 24378 0 net167
rlabel metal1 11132 25262 11132 25262 0 net168
rlabel metal1 14306 33082 14306 33082 0 net169
rlabel metal1 3358 21522 3358 21522 0 net17
rlabel metal1 12972 23698 12972 23698 0 net170
rlabel metal2 16514 40358 16514 40358 0 net171
rlabel metal2 14030 39202 14030 39202 0 net172
rlabel metal1 16238 38964 16238 38964 0 net173
rlabel metal1 12696 35258 12696 35258 0 net174
rlabel metal1 11408 35666 11408 35666 0 net175
rlabel metal1 13340 39066 13340 39066 0 net176
rlabel metal1 12236 43418 12236 43418 0 net177
rlabel metal1 12972 42330 12972 42330 0 net178
rlabel metal2 10810 43792 10810 43792 0 net179
rlabel metal1 2668 22066 2668 22066 0 net18
rlabel metal1 7866 39950 7866 39950 0 net180
rlabel metal1 12351 23086 12351 23086 0 net181
rlabel metal1 8280 40494 8280 40494 0 net182
rlabel metal2 12558 44302 12558 44302 0 net183
rlabel metal2 11822 36550 11822 36550 0 net184
rlabel metal1 11362 37842 11362 37842 0 net185
rlabel metal1 12052 39406 12052 39406 0 net186
rlabel metal1 18354 38930 18354 38930 0 net187
rlabel metal1 15916 32878 15916 32878 0 net188
rlabel metal1 14904 31790 14904 31790 0 net189
rlabel metal1 3910 23154 3910 23154 0 net19
rlabel metal2 11914 33490 11914 33490 0 net190
rlabel metal1 7636 32402 7636 32402 0 net191
rlabel metal2 16882 37842 16882 37842 0 net192
rlabel metal1 16284 40086 16284 40086 0 net193
rlabel metal2 20930 44166 20930 44166 0 net194
rlabel metal1 14168 51442 14168 51442 0 net195
rlabel metal1 16698 51782 16698 51782 0 net196
rlabel metal1 14260 47770 14260 47770 0 net197
rlabel metal1 16606 44370 16606 44370 0 net198
rlabel metal1 33212 2822 33212 2822 0 net199
rlabel metal2 47058 52122 47058 52122 0 net2
rlabel metal1 2714 23698 2714 23698 0 net20
rlabel metal1 3404 24786 3404 24786 0 net21
rlabel metal1 3450 25330 3450 25330 0 net22
rlabel metal2 2530 42466 2530 42466 0 net23
rlabel metal1 4186 27030 4186 27030 0 net24
rlabel metal1 5566 5270 5566 5270 0 net25
rlabel metal1 6670 5542 6670 5542 0 net26
rlabel metal1 4830 6834 4830 6834 0 net27
rlabel metal1 6026 7174 6026 7174 0 net28
rlabel metal1 6256 8330 6256 8330 0 net29
rlabel metal1 7222 3502 7222 3502 0 net3
rlabel metal2 1610 17034 1610 17034 0 net30
rlabel metal1 6256 9894 6256 9894 0 net31
rlabel metal1 7314 10438 7314 10438 0 net32
rlabel metal1 21666 52870 21666 52870 0 net33
rlabel metal1 13984 50966 13984 50966 0 net34
rlabel metal1 10396 38250 10396 38250 0 net35
rlabel via2 9614 36907 9614 36907 0 net36
rlabel metal1 27692 49198 27692 49198 0 net37
rlabel metal1 27508 49946 27508 49946 0 net38
rlabel metal1 27416 53686 27416 53686 0 net39
rlabel metal1 6394 11526 6394 11526 0 net4
rlabel metal1 31970 53448 31970 53448 0 net40
rlabel metal2 32798 54434 32798 54434 0 net41
rlabel metal1 20194 54130 20194 54130 0 net42
rlabel metal2 34270 47549 34270 47549 0 net43
rlabel metal2 18446 52237 18446 52237 0 net44
rlabel metal2 35098 54009 35098 54009 0 net45
rlabel metal2 33810 51544 33810 51544 0 net46
rlabel metal1 36087 54026 36087 54026 0 net47
rlabel metal1 33442 53754 33442 53754 0 net48
rlabel metal2 33534 50116 33534 50116 0 net49
rlabel metal1 6900 12070 6900 12070 0 net5
rlabel metal1 37904 53958 37904 53958 0 net50
rlabel metal2 38686 46648 38686 46648 0 net51
rlabel metal2 38962 44088 38962 44088 0 net52
rlabel metal2 40250 44156 40250 44156 0 net53
rlabel metal2 40066 50694 40066 50694 0 net54
rlabel metal1 18170 49946 18170 49946 0 net55
rlabel metal1 20654 54060 20654 54060 0 net56
rlabel metal2 18538 52666 18538 52666 0 net57
rlabel metal2 20010 52870 20010 52870 0 net58
rlabel metal1 21482 50966 21482 50966 0 net59
rlabel metal1 7176 13158 7176 13158 0 net6
rlabel metal1 24886 54298 24886 54298 0 net60
rlabel metal1 20838 49300 20838 49300 0 net61
rlabel metal2 12742 52258 12742 52258 0 net62
rlabel metal2 24978 10098 24978 10098 0 net63
rlabel metal1 31510 2346 31510 2346 0 net64
rlabel metal1 37421 2482 37421 2482 0 net65
rlabel metal1 42918 2550 42918 2550 0 net66
rlabel metal1 21804 11118 21804 11118 0 net67
rlabel metal1 23085 17238 23085 17238 0 net68
rlabel metal2 46138 47600 46138 47600 0 net69
rlabel metal1 1656 14042 1656 14042 0 net7
rlabel metal2 46874 49402 46874 49402 0 net70
rlabel metal2 46966 46886 46966 46886 0 net71
rlabel metal1 47886 53958 47886 53958 0 net72
rlabel metal2 48622 44615 48622 44615 0 net73
rlabel metal2 48898 46138 48898 46138 0 net74
rlabel metal2 44390 49096 44390 49096 0 net75
rlabel metal1 45356 53958 45356 53958 0 net76
rlabel metal2 49082 44336 49082 44336 0 net77
rlabel metal2 49266 46886 49266 46886 0 net78
rlabel metal1 49082 47770 49082 47770 0 net79
rlabel metal1 4416 14994 4416 14994 0 net8
rlabel metal1 49036 52870 49036 52870 0 net80
rlabel metal2 34362 22474 34362 22474 0 net81
rlabel metal1 2990 52462 2990 52462 0 net82
rlabel metal1 4347 28050 4347 28050 0 net83
rlabel metal2 4094 37978 4094 37978 0 net84
rlabel metal2 1794 39236 1794 39236 0 net85
rlabel metal1 2277 37842 2277 37842 0 net86
rlabel metal1 2277 38318 2277 38318 0 net87
rlabel metal2 4646 38964 4646 38964 0 net88
rlabel metal1 1794 40052 1794 40052 0 net89
rlabel metal1 4784 15606 4784 15606 0 net9
rlabel metal1 6854 41140 6854 41140 0 net90
rlabel metal1 2277 41582 2277 41582 0 net91
rlabel metal2 1610 46546 1610 46546 0 net92
rlabel metal2 5382 46512 5382 46512 0 net93
rlabel metal2 1794 28577 1794 28577 0 net94
rlabel metal1 2277 44370 2277 44370 0 net95
rlabel metal2 4370 43316 4370 43316 0 net96
rlabel metal2 3726 44336 3726 44336 0 net97
rlabel metal1 2277 46546 2277 46546 0 net98
rlabel metal2 4186 46070 4186 46070 0 net99
rlabel metal2 48622 1894 48622 1894 0 prog_clk
rlabel metal1 42412 54230 42412 54230 0 prog_reset_top_in
rlabel metal1 17480 42738 17480 42738 0 sb_8__0_.mem_left_track_1.ccff_head
rlabel metal1 20378 44710 20378 44710 0 sb_8__0_.mem_left_track_1.ccff_tail
rlabel metal1 20838 44268 20838 44268 0 sb_8__0_.mem_left_track_1.mem_out\[0\]
rlabel metal1 14168 50218 14168 50218 0 sb_8__0_.mem_left_track_11.ccff_head
rlabel metal1 16100 51306 16100 51306 0 sb_8__0_.mem_left_track_11.ccff_tail
rlabel metal1 17388 51442 17388 51442 0 sb_8__0_.mem_left_track_11.mem_out\[0\]
rlabel metal2 17434 50524 17434 50524 0 sb_8__0_.mem_left_track_13.ccff_tail
rlabel metal1 18860 51510 18860 51510 0 sb_8__0_.mem_left_track_13.mem_out\[0\]
rlabel metal1 18170 48178 18170 48178 0 sb_8__0_.mem_left_track_15.ccff_tail
rlabel metal1 18354 50150 18354 50150 0 sb_8__0_.mem_left_track_15.mem_out\[0\]
rlabel metal2 17434 47260 17434 47260 0 sb_8__0_.mem_left_track_17.ccff_tail
rlabel metal1 18952 47974 18952 47974 0 sb_8__0_.mem_left_track_17.mem_out\[0\]
rlabel metal1 18860 46342 18860 46342 0 sb_8__0_.mem_left_track_19.ccff_tail
rlabel metal1 18998 47226 18998 47226 0 sb_8__0_.mem_left_track_19.mem_out\[0\]
rlabel metal2 20010 45390 20010 45390 0 sb_8__0_.mem_left_track_29.ccff_tail
rlabel metal1 21528 47226 21528 47226 0 sb_8__0_.mem_left_track_29.mem_out\[0\]
rlabel metal1 13938 47090 13938 47090 0 sb_8__0_.mem_left_track_3.ccff_tail
rlabel metal1 18170 46138 18170 46138 0 sb_8__0_.mem_left_track_3.mem_out\[0\]
rlabel metal2 21482 46376 21482 46376 0 sb_8__0_.mem_left_track_31.ccff_tail
rlabel metal1 21666 46682 21666 46682 0 sb_8__0_.mem_left_track_31.mem_out\[0\]
rlabel metal1 20746 50218 20746 50218 0 sb_8__0_.mem_left_track_33.ccff_tail
rlabel metal2 21114 49232 21114 49232 0 sb_8__0_.mem_left_track_33.mem_out\[0\]
rlabel metal1 20286 48212 20286 48212 0 sb_8__0_.mem_left_track_35.ccff_tail
rlabel metal2 22678 50048 22678 50048 0 sb_8__0_.mem_left_track_35.mem_out\[0\]
rlabel metal1 19458 45356 19458 45356 0 sb_8__0_.mem_left_track_45.ccff_tail
rlabel metal1 25070 48246 25070 48246 0 sb_8__0_.mem_left_track_45.mem_out\[0\]
rlabel metal2 22678 45696 22678 45696 0 sb_8__0_.mem_left_track_47.ccff_tail
rlabel metal2 24794 46784 24794 46784 0 sb_8__0_.mem_left_track_47.mem_out\[0\]
rlabel via1 23598 43826 23598 43826 0 sb_8__0_.mem_left_track_49.ccff_tail
rlabel metal1 24242 46682 24242 46682 0 sb_8__0_.mem_left_track_49.mem_out\[0\]
rlabel metal1 14628 46954 14628 46954 0 sb_8__0_.mem_left_track_5.ccff_tail
rlabel metal1 15088 47566 15088 47566 0 sb_8__0_.mem_left_track_5.mem_out\[0\]
rlabel metal2 24058 45186 24058 45186 0 sb_8__0_.mem_left_track_51.mem_out\[0\]
rlabel metal2 14030 46308 14030 46308 0 sb_8__0_.mem_left_track_7.ccff_tail
rlabel metal2 16054 48450 16054 48450 0 sb_8__0_.mem_left_track_7.mem_out\[0\]
rlabel via1 16514 49283 16514 49283 0 sb_8__0_.mem_left_track_9.mem_out\[0\]
rlabel metal2 21390 42772 21390 42772 0 sb_8__0_.mem_top_track_0.ccff_tail
rlabel metal1 27554 44914 27554 44914 0 sb_8__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 18722 41684 18722 41684 0 sb_8__0_.mem_top_track_0.mem_out\[1\]
rlabel metal1 19918 36550 19918 36550 0 sb_8__0_.mem_top_track_10.ccff_head
rlabel metal1 17572 34646 17572 34646 0 sb_8__0_.mem_top_track_10.ccff_tail
rlabel metal1 20010 35768 20010 35768 0 sb_8__0_.mem_top_track_10.mem_out\[0\]
rlabel metal1 17388 34986 17388 34986 0 sb_8__0_.mem_top_track_10.mem_out\[1\]
rlabel metal1 18124 33830 18124 33830 0 sb_8__0_.mem_top_track_12.ccff_tail
rlabel metal1 16560 33898 16560 33898 0 sb_8__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 14996 33422 14996 33422 0 sb_8__0_.mem_top_track_14.ccff_tail
rlabel metal1 17802 31994 17802 31994 0 sb_8__0_.mem_top_track_14.mem_out\[0\]
rlabel metal2 14858 33524 14858 33524 0 sb_8__0_.mem_top_track_16.ccff_tail
rlabel metal1 17802 36210 17802 36210 0 sb_8__0_.mem_top_track_16.mem_out\[0\]
rlabel metal1 18032 37774 18032 37774 0 sb_8__0_.mem_top_track_18.ccff_tail
rlabel metal1 18124 37298 18124 37298 0 sb_8__0_.mem_top_track_18.mem_out\[0\]
rlabel metal2 19090 33728 19090 33728 0 sb_8__0_.mem_top_track_2.ccff_tail
rlabel metal1 21022 34408 21022 34408 0 sb_8__0_.mem_top_track_2.mem_out\[0\]
rlabel metal1 21666 34714 21666 34714 0 sb_8__0_.mem_top_track_2.mem_out\[1\]
rlabel metal1 18078 38454 18078 38454 0 sb_8__0_.mem_top_track_20.ccff_tail
rlabel metal1 16744 38250 16744 38250 0 sb_8__0_.mem_top_track_20.mem_out\[0\]
rlabel metal1 15824 38182 15824 38182 0 sb_8__0_.mem_top_track_22.ccff_tail
rlabel metal2 14858 37468 14858 37468 0 sb_8__0_.mem_top_track_22.mem_out\[0\]
rlabel metal1 15456 36346 15456 36346 0 sb_8__0_.mem_top_track_24.ccff_tail
rlabel metal2 16054 36448 16054 36448 0 sb_8__0_.mem_top_track_24.mem_out\[0\]
rlabel metal1 13984 32334 13984 32334 0 sb_8__0_.mem_top_track_26.ccff_tail
rlabel metal1 13018 32334 13018 32334 0 sb_8__0_.mem_top_track_26.mem_out\[0\]
rlabel metal2 12374 35122 12374 35122 0 sb_8__0_.mem_top_track_28.ccff_tail
rlabel metal1 12006 31892 12006 31892 0 sb_8__0_.mem_top_track_28.mem_out\[0\]
rlabel metal2 13570 36550 13570 36550 0 sb_8__0_.mem_top_track_30.ccff_tail
rlabel metal2 13570 35360 13570 35360 0 sb_8__0_.mem_top_track_30.mem_out\[0\]
rlabel metal1 11776 39950 11776 39950 0 sb_8__0_.mem_top_track_32.ccff_tail
rlabel metal2 13110 37978 13110 37978 0 sb_8__0_.mem_top_track_32.mem_out\[0\]
rlabel metal1 13662 42058 13662 42058 0 sb_8__0_.mem_top_track_34.ccff_tail
rlabel metal1 13386 39950 13386 39950 0 sb_8__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 11040 40902 11040 40902 0 sb_8__0_.mem_top_track_36.ccff_tail
rlabel metal1 12236 41446 12236 41446 0 sb_8__0_.mem_top_track_36.mem_out\[0\]
rlabel metal1 8970 38454 8970 38454 0 sb_8__0_.mem_top_track_38.ccff_tail
rlabel metal1 8004 38386 8004 38386 0 sb_8__0_.mem_top_track_38.mem_out\[0\]
rlabel metal1 18446 33422 18446 33422 0 sb_8__0_.mem_top_track_4.ccff_tail
rlabel metal1 21390 34170 21390 34170 0 sb_8__0_.mem_top_track_4.mem_out\[0\]
rlabel metal1 20884 32538 20884 32538 0 sb_8__0_.mem_top_track_4.mem_out\[1\]
rlabel metal1 8740 40562 8740 40562 0 sb_8__0_.mem_top_track_40.ccff_tail
rlabel metal2 8602 38624 8602 38624 0 sb_8__0_.mem_top_track_40.mem_out\[0\]
rlabel metal1 11684 42874 11684 42874 0 sb_8__0_.mem_top_track_42.ccff_tail
rlabel metal2 10534 40783 10534 40783 0 sb_8__0_.mem_top_track_42.mem_out\[0\]
rlabel metal1 14352 40426 14352 40426 0 sb_8__0_.mem_top_track_44.ccff_tail
rlabel metal1 15548 40902 15548 40902 0 sb_8__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 16054 41242 16054 41242 0 sb_8__0_.mem_top_track_46.ccff_tail
rlabel metal1 14536 41038 14536 41038 0 sb_8__0_.mem_top_track_46.mem_out\[0\]
rlabel metal1 15134 42738 15134 42738 0 sb_8__0_.mem_top_track_48.ccff_tail
rlabel metal2 20378 41820 20378 41820 0 sb_8__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 13570 38760 13570 38760 0 sb_8__0_.mem_top_track_50.mem_out\[0\]
rlabel metal2 20010 39576 20010 39576 0 sb_8__0_.mem_top_track_6.ccff_tail
rlabel metal2 21942 38046 21942 38046 0 sb_8__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 19228 38862 19228 38862 0 sb_8__0_.mem_top_track_6.mem_out\[1\]
rlabel metal2 21482 39100 21482 39100 0 sb_8__0_.mem_top_track_8.mem_out\[0\]
rlabel metal1 19320 36822 19320 36822 0 sb_8__0_.mem_top_track_8.mem_out\[1\]
rlabel metal1 13386 43112 13386 43112 0 sb_8__0_.mux_left_track_1.out
rlabel metal1 23966 43656 23966 43656 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19918 44098 19918 44098 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15778 43350 15778 43350 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 6118 36142 6118 36142 0 sb_8__0_.mux_left_track_11.out
rlabel metal1 17802 51238 17802 51238 0 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 9982 47124 9982 47124 0 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7820 37230 7820 37230 0 sb_8__0_.mux_left_track_13.out
rlabel metal2 19550 51149 19550 51149 0 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15226 46954 15226 46954 0 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5842 35734 5842 35734 0 sb_8__0_.mux_left_track_15.out
rlabel metal1 17802 47770 17802 47770 0 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14766 46172 14766 46172 0 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7682 42534 7682 42534 0 sb_8__0_.mux_left_track_17.out
rlabel metal1 16560 44710 16560 44710 0 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X
rlabel via1 15134 42245 15134 42245 0 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7084 36890 7084 36890 0 sb_8__0_.mux_left_track_19.out
rlabel metal1 17618 44846 17618 44846 0 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12558 41752 12558 41752 0 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5428 37842 5428 37842 0 sb_8__0_.mux_left_track_29.out
rlabel metal1 19826 44370 19826 44370 0 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13018 43792 13018 43792 0 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7314 45050 7314 45050 0 sb_8__0_.mux_left_track_3.out
rlabel metal1 13754 47022 13754 47022 0 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12742 46070 12742 46070 0 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 8234 35054 8234 35054 0 sb_8__0_.mux_left_track_31.out
rlabel metal1 18630 44982 18630 44982 0 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13800 43758 13800 43758 0 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 10902 43554 10902 43554 0 sb_8__0_.mux_left_track_33.out
rlabel metal1 19366 48620 19366 48620 0 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12742 45492 12742 45492 0 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 13110 44710 13110 44710 0 sb_8__0_.mux_left_track_35.out
rlabel metal1 20930 48042 20930 48042 0 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13846 44846 13846 44846 0 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6992 38998 6992 38998 0 sb_8__0_.mux_left_track_45.out
rlabel metal1 19412 45594 19412 45594 0 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14766 43758 14766 43758 0 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13478 43316 13478 43316 0 sb_8__0_.mux_left_track_47.out
rlabel metal1 23552 44846 23552 44846 0 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13846 43282 13846 43282 0 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13662 34680 13662 34680 0 sb_8__0_.mux_left_track_49.out
rlabel metal2 22494 45424 22494 45424 0 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 17894 42602 17894 42602 0 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5704 39066 5704 39066 0 sb_8__0_.mux_left_track_5.out
rlabel metal2 13570 48144 13570 48144 0 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 8786 45764 8786 45764 0 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8418 32402 8418 32402 0 sb_8__0_.mux_left_track_51.out
rlabel metal1 20838 42534 20838 42534 0 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18538 36550 18538 36550 0 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 5796 38318 5796 38318 0 sb_8__0_.mux_left_track_7.out
rlabel metal1 14996 46682 14996 46682 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15042 45322 15042 45322 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 11362 45084 11362 45084 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 5934 36890 5934 36890 0 sb_8__0_.mux_left_track_9.out
rlabel metal1 13662 48110 13662 48110 0 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 12650 46750 12650 46750 0 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21160 47974 21160 47974 0 sb_8__0_.mux_top_track_0.out
rlabel metal1 25944 43758 25944 43758 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 26128 43690 26128 43690 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 24610 43486 24610 43486 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19458 41786 19458 41786 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21022 43418 21022 43418 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 17756 51986 17756 51986 0 sb_8__0_.mux_top_track_10.out
rlabel metal1 22586 36890 22586 36890 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22402 37536 22402 37536 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16330 35802 16330 35802 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15042 35666 15042 35666 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 16468 35462 16468 35462 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 15870 43078 15870 43078 0 sb_8__0_.mux_top_track_12.out
rlabel metal1 17618 35802 17618 35802 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14444 33524 14444 33524 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16422 35530 16422 35530 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 16744 41990 16744 41990 0 sb_8__0_.mux_top_track_14.out
rlabel metal1 14674 33388 14674 33388 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12190 24378 12190 24378 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 15962 41820 15962 41820 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17112 43078 17112 43078 0 sb_8__0_.mux_top_track_16.out
rlabel metal1 15548 35054 15548 35054 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13800 34986 13800 34986 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15134 34918 15134 34918 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15134 51986 15134 51986 0 sb_8__0_.mux_top_track_18.out
rlabel metal1 18906 39338 18906 39338 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 15088 33286 15088 33286 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16928 43180 16928 43180 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17986 41718 17986 41718 0 sb_8__0_.mux_top_track_2.out
rlabel metal2 21758 37332 21758 37332 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21666 36924 21666 36924 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20102 33626 20102 33626 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15456 23834 15456 23834 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18492 33626 18492 33626 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 13984 51374 13984 51374 0 sb_8__0_.mux_top_track_20.out
rlabel metal1 15962 35258 15962 35258 0 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 16698 41242 16698 41242 0 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13570 45254 13570 45254 0 sb_8__0_.mux_top_track_22.out
rlabel metal1 14812 36618 14812 36618 0 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 14766 39610 14766 39610 0 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14306 44744 14306 44744 0 sb_8__0_.mux_top_track_24.out
rlabel metal2 15502 37910 15502 37910 0 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 14214 39168 14214 39168 0 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 12006 47158 12006 47158 0 sb_8__0_.mux_top_track_26.out
rlabel metal2 13386 34374 13386 34374 0 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12650 36346 12650 36346 0 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 9798 46274 9798 46274 0 sb_8__0_.mux_top_track_28.out
rlabel metal1 11638 27574 11638 27574 0 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10258 35802 10258 35802 0 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11500 45050 11500 45050 0 sb_8__0_.mux_top_track_30.out
rlabel metal1 13248 35258 13248 35258 0 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13110 39066 13110 39066 0 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 11178 46138 11178 46138 0 sb_8__0_.mux_top_track_32.out
rlabel metal2 12328 40324 12328 40324 0 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11592 43418 11592 43418 0 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10442 47770 10442 47770 0 sb_8__0_.mux_top_track_34.out
rlabel metal1 12374 39066 12374 39066 0 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11638 44880 11638 44880 0 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9798 47770 9798 47770 0 sb_8__0_.mux_top_track_36.out
rlabel metal1 12788 40698 12788 40698 0 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10166 43418 10166 43418 0 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7820 45322 7820 45322 0 sb_8__0_.mux_top_track_38.out
rlabel metal2 8786 37570 8786 37570 0 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8648 45458 8648 45458 0 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 17802 42330 17802 42330 0 sb_8__0_.mux_top_track_4.out
rlabel metal1 20976 34986 20976 34986 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20838 35054 20838 35054 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 18032 33626 18032 33626 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 14766 23290 14766 23290 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17020 33626 17020 33626 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 7958 46138 7958 46138 0 sb_8__0_.mux_top_track_40.out
rlabel metal1 7912 35802 7912 35802 0 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7820 40698 7820 40698 0 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9430 48858 9430 48858 0 sb_8__0_.mux_top_track_42.out
rlabel metal1 13294 39610 13294 39610 0 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11270 46342 11270 46342 0 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 10212 51374 10212 51374 0 sb_8__0_.mux_top_track_44.out
rlabel metal1 18630 41990 18630 41990 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10534 36890 10534 36890 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12834 41786 12834 41786 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9614 51306 9614 51306 0 sb_8__0_.mux_top_track_46.out
rlabel via2 14766 41667 14766 41667 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13984 41514 13984 41514 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14306 41854 14306 41854 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 9614 51918 9614 51918 0 sb_8__0_.mux_top_track_48.out
rlabel metal1 19642 42330 19642 42330 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 12466 39933 12466 39933 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14168 42534 14168 42534 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 8188 51986 8188 51986 0 sb_8__0_.mux_top_track_50.out
rlabel metal1 18630 42058 18630 42058 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10718 39610 10718 39610 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 14214 43418 14214 43418 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19044 51986 19044 51986 0 sb_8__0_.mux_top_track_6.out
rlabel metal1 22908 41446 22908 41446 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23460 41514 23460 41514 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20148 39270 20148 39270 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 17112 33082 17112 33082 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 18308 39610 18308 39610 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 19780 44166 19780 44166 0 sb_8__0_.mux_top_track_8.out
rlabel metal1 23644 39338 23644 39338 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23460 39406 23460 39406 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17434 36516 17434 36516 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 14950 32096 14950 32096 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 17342 36550 17342 36550 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 45402 55413 45402 55413 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
rlabel metal1 46368 54162 46368 54162 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
rlabel metal1 46736 53550 46736 53550 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
rlabel metal1 47564 54162 47564 54162 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
rlabel metal2 47978 55711 47978 55711 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
rlabel metal1 48668 53550 48668 53550 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
rlabel metal1 44160 53550 44160 53550 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
rlabel metal1 44988 54162 44988 54162 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
rlabel via2 48990 48059 48990 48059 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel via2 49082 50269 49082 50269 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
rlabel via2 49082 52445 49082 52445 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 49082 53839 49082 53839 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal3 2016 52156 2016 52156 0 top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 2154 52972 2154 52972 0 top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 1740 53788 1740 53788 0 top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 2062 54604 2062 54604 0 top_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 57000
<< end >>
