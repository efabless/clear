magic
tech sky130A
magscale 1 2
timestamp 1656242503
<< obsli1 >>
rect 1104 2159 21896 20689
<< obsm1 >>
rect 1104 2128 22434 20868
<< metal2 >>
rect 1674 22200 1730 23000
rect 2042 22200 2098 23000
rect 2410 22200 2466 23000
rect 2778 22200 2834 23000
rect 3146 22200 3202 23000
rect 3514 22200 3570 23000
rect 3882 22200 3938 23000
rect 4250 22200 4306 23000
rect 4618 22200 4674 23000
rect 4986 22200 5042 23000
rect 5354 22200 5410 23000
rect 5722 22200 5778 23000
rect 6090 22200 6146 23000
rect 6458 22200 6514 23000
rect 6826 22200 6882 23000
rect 7194 22200 7250 23000
rect 7562 22200 7618 23000
rect 7930 22200 7986 23000
rect 8298 22200 8354 23000
rect 8666 22200 8722 23000
rect 9034 22200 9090 23000
rect 9402 22200 9458 23000
rect 9770 22200 9826 23000
rect 10138 22200 10194 23000
rect 10506 22200 10562 23000
rect 10874 22200 10930 23000
rect 11242 22200 11298 23000
rect 11610 22200 11666 23000
rect 11978 22200 12034 23000
rect 12346 22200 12402 23000
rect 12714 22200 12770 23000
rect 13082 22200 13138 23000
rect 13450 22200 13506 23000
rect 13818 22200 13874 23000
rect 14186 22200 14242 23000
rect 14554 22200 14610 23000
rect 14922 22200 14978 23000
rect 15290 22200 15346 23000
rect 15658 22200 15714 23000
rect 16026 22200 16082 23000
rect 16394 22200 16450 23000
rect 16762 22200 16818 23000
rect 17130 22200 17186 23000
rect 17498 22200 17554 23000
rect 17866 22200 17922 23000
rect 18234 22200 18290 23000
rect 18602 22200 18658 23000
rect 18970 22200 19026 23000
rect 19338 22200 19394 23000
rect 19706 22200 19762 23000
rect 20074 22200 20130 23000
rect 20442 22200 20498 23000
rect 20810 22200 20866 23000
rect 21178 22200 21234 23000
rect 2226 0 2282 800
rect 6826 0 6882 800
rect 11426 0 11482 800
rect 16026 0 16082 800
rect 20626 0 20682 800
<< obsm2 >>
rect 1306 22144 1618 22250
rect 1786 22144 1986 22250
rect 2154 22144 2354 22250
rect 2522 22144 2722 22250
rect 2890 22144 3090 22250
rect 3258 22144 3458 22250
rect 3626 22144 3826 22250
rect 3994 22144 4194 22250
rect 4362 22144 4562 22250
rect 4730 22144 4930 22250
rect 5098 22144 5298 22250
rect 5466 22144 5666 22250
rect 5834 22144 6034 22250
rect 6202 22144 6402 22250
rect 6570 22144 6770 22250
rect 6938 22144 7138 22250
rect 7306 22144 7506 22250
rect 7674 22144 7874 22250
rect 8042 22144 8242 22250
rect 8410 22144 8610 22250
rect 8778 22144 8978 22250
rect 9146 22144 9346 22250
rect 9514 22144 9714 22250
rect 9882 22144 10082 22250
rect 10250 22144 10450 22250
rect 10618 22144 10818 22250
rect 10986 22144 11186 22250
rect 11354 22144 11554 22250
rect 11722 22144 11922 22250
rect 12090 22144 12290 22250
rect 12458 22144 12658 22250
rect 12826 22144 13026 22250
rect 13194 22144 13394 22250
rect 13562 22144 13762 22250
rect 13930 22144 14130 22250
rect 14298 22144 14498 22250
rect 14666 22144 14866 22250
rect 15034 22144 15234 22250
rect 15402 22144 15602 22250
rect 15770 22144 15970 22250
rect 16138 22144 16338 22250
rect 16506 22144 16706 22250
rect 16874 22144 17074 22250
rect 17242 22144 17442 22250
rect 17610 22144 17810 22250
rect 17978 22144 18178 22250
rect 18346 22144 18546 22250
rect 18714 22144 18914 22250
rect 19082 22144 19282 22250
rect 19450 22144 19650 22250
rect 19818 22144 20018 22250
rect 20186 22144 20386 22250
rect 20554 22144 20754 22250
rect 20922 22144 21122 22250
rect 21290 22144 22428 22250
rect 1306 856 22428 22144
rect 1306 734 2170 856
rect 2338 734 6770 856
rect 6938 734 11370 856
rect 11538 734 15970 856
rect 16138 734 20570 856
rect 20738 734 22428 856
<< metal3 >>
rect 0 21224 800 21344
rect 22200 21224 23000 21344
rect 0 20816 800 20936
rect 22200 20816 23000 20936
rect 0 20408 800 20528
rect 22200 20408 23000 20528
rect 0 20000 800 20120
rect 22200 20000 23000 20120
rect 0 19592 800 19712
rect 22200 19592 23000 19712
rect 0 19184 800 19304
rect 22200 19184 23000 19304
rect 0 18776 800 18896
rect 22200 18776 23000 18896
rect 0 18368 800 18488
rect 22200 18368 23000 18488
rect 0 17960 800 18080
rect 22200 17960 23000 18080
rect 0 17552 800 17672
rect 22200 17552 23000 17672
rect 0 17144 800 17264
rect 22200 17144 23000 17264
rect 0 16736 800 16856
rect 22200 16736 23000 16856
rect 0 16328 800 16448
rect 22200 16328 23000 16448
rect 0 15920 800 16040
rect 22200 15920 23000 16040
rect 0 15512 800 15632
rect 22200 15512 23000 15632
rect 0 15104 800 15224
rect 22200 15104 23000 15224
rect 0 14696 800 14816
rect 22200 14696 23000 14816
rect 0 14288 800 14408
rect 22200 14288 23000 14408
rect 0 13880 800 14000
rect 22200 13880 23000 14000
rect 0 13472 800 13592
rect 22200 13472 23000 13592
rect 0 13064 800 13184
rect 22200 13064 23000 13184
rect 0 12656 800 12776
rect 22200 12656 23000 12776
rect 0 12248 800 12368
rect 22200 12248 23000 12368
rect 0 11840 800 11960
rect 22200 11840 23000 11960
rect 0 11432 800 11552
rect 22200 11432 23000 11552
rect 0 11024 800 11144
rect 22200 11024 23000 11144
rect 0 10616 800 10736
rect 22200 10616 23000 10736
rect 0 10208 800 10328
rect 22200 10208 23000 10328
rect 0 9800 800 9920
rect 22200 9800 23000 9920
rect 0 9392 800 9512
rect 22200 9392 23000 9512
rect 0 8984 800 9104
rect 22200 8984 23000 9104
rect 0 8576 800 8696
rect 22200 8576 23000 8696
rect 0 8168 800 8288
rect 22200 8168 23000 8288
rect 0 7760 800 7880
rect 22200 7760 23000 7880
rect 0 7352 800 7472
rect 22200 7352 23000 7472
rect 0 6944 800 7064
rect 22200 6944 23000 7064
rect 0 6536 800 6656
rect 22200 6536 23000 6656
rect 0 6128 800 6248
rect 22200 6128 23000 6248
rect 0 5720 800 5840
rect 22200 5720 23000 5840
rect 0 5312 800 5432
rect 22200 5312 23000 5432
rect 0 4904 800 5024
rect 22200 4904 23000 5024
rect 0 4496 800 4616
rect 22200 4496 23000 4616
rect 0 4088 800 4208
rect 22200 4088 23000 4208
rect 0 3680 800 3800
rect 22200 3680 23000 3800
rect 0 3272 800 3392
rect 22200 3272 23000 3392
rect 0 2864 800 2984
rect 22200 2864 23000 2984
rect 0 2456 800 2576
rect 22200 2456 23000 2576
rect 0 2048 800 2168
rect 22200 2048 23000 2168
rect 0 1640 800 1760
rect 22200 1640 23000 1760
<< obsm3 >>
rect 880 21144 22120 21317
rect 800 21016 22202 21144
rect 880 20736 22120 21016
rect 800 20608 22202 20736
rect 880 20328 22120 20608
rect 800 20200 22202 20328
rect 880 19920 22120 20200
rect 800 19792 22202 19920
rect 880 19512 22120 19792
rect 800 19384 22202 19512
rect 880 19104 22120 19384
rect 800 18976 22202 19104
rect 880 18696 22120 18976
rect 800 18568 22202 18696
rect 880 18288 22120 18568
rect 800 18160 22202 18288
rect 880 17880 22120 18160
rect 800 17752 22202 17880
rect 880 17472 22120 17752
rect 800 17344 22202 17472
rect 880 17064 22120 17344
rect 800 16936 22202 17064
rect 880 16656 22120 16936
rect 800 16528 22202 16656
rect 880 16248 22120 16528
rect 800 16120 22202 16248
rect 880 15840 22120 16120
rect 800 15712 22202 15840
rect 880 15432 22120 15712
rect 800 15304 22202 15432
rect 880 15024 22120 15304
rect 800 14896 22202 15024
rect 880 14616 22120 14896
rect 800 14488 22202 14616
rect 880 14208 22120 14488
rect 800 14080 22202 14208
rect 880 13800 22120 14080
rect 800 13672 22202 13800
rect 880 13392 22120 13672
rect 800 13264 22202 13392
rect 880 12984 22120 13264
rect 800 12856 22202 12984
rect 880 12576 22120 12856
rect 800 12448 22202 12576
rect 880 12168 22120 12448
rect 800 12040 22202 12168
rect 880 11760 22120 12040
rect 800 11632 22202 11760
rect 880 11352 22120 11632
rect 800 11224 22202 11352
rect 880 10944 22120 11224
rect 800 10816 22202 10944
rect 880 10536 22120 10816
rect 800 10408 22202 10536
rect 880 10128 22120 10408
rect 800 10000 22202 10128
rect 880 9720 22120 10000
rect 800 9592 22202 9720
rect 880 9312 22120 9592
rect 800 9184 22202 9312
rect 880 8904 22120 9184
rect 800 8776 22202 8904
rect 880 8496 22120 8776
rect 800 8368 22202 8496
rect 880 8088 22120 8368
rect 800 7960 22202 8088
rect 880 7680 22120 7960
rect 800 7552 22202 7680
rect 880 7272 22120 7552
rect 800 7144 22202 7272
rect 880 6864 22120 7144
rect 800 6736 22202 6864
rect 880 6456 22120 6736
rect 800 6328 22202 6456
rect 880 6048 22120 6328
rect 800 5920 22202 6048
rect 880 5640 22120 5920
rect 800 5512 22202 5640
rect 880 5232 22120 5512
rect 800 5104 22202 5232
rect 880 4824 22120 5104
rect 800 4696 22202 4824
rect 880 4416 22120 4696
rect 800 4288 22202 4416
rect 880 4008 22120 4288
rect 800 3880 22202 4008
rect 880 3600 22120 3880
rect 800 3472 22202 3600
rect 880 3192 22120 3472
rect 800 3064 22202 3192
rect 880 2784 22120 3064
rect 800 2656 22202 2784
rect 880 2376 22120 2656
rect 800 2248 22202 2376
rect 880 1968 22120 2248
rect 800 1840 22202 1968
rect 880 1667 22120 1840
<< metal4 >>
rect 3543 2128 3863 20720
rect 6142 2128 6462 20720
rect 8741 2128 9061 20720
rect 11340 2128 11660 20720
rect 13939 2128 14259 20720
rect 16538 2128 16858 20720
rect 19137 2128 19457 20720
rect 21736 2128 22056 20720
<< obsm4 >>
rect 3943 2891 6062 20229
rect 6542 2891 8661 20229
rect 9141 2891 11260 20229
rect 11740 2891 13859 20229
rect 14339 2891 16458 20229
rect 16938 2891 19057 20229
rect 19537 2891 20549 20229
<< labels >>
rlabel metal2 s 1674 22200 1730 23000 6 SC_IN_TOP
port 1 nsew signal input
rlabel metal2 s 21178 22200 21234 23000 6 SC_OUT_TOP
port 2 nsew signal output
rlabel metal2 s 5354 22200 5410 23000 6 Test_en_N_out
port 3 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 Test_en_S_in
port 4 nsew signal input
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 5 nsew ground bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 5 nsew ground bidirectional
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 5 nsew ground bidirectional
rlabel metal4 s 21736 2128 22056 20720 6 VGND
port 5 nsew ground bidirectional
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 6 nsew power bidirectional
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 6 nsew power bidirectional
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 6 nsew power bidirectional
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 6 nsew power bidirectional
rlabel metal2 s 2226 0 2282 800 6 ccff_head
port 7 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 ccff_tail
port 8 nsew signal output
rlabel metal3 s 0 5312 800 5432 6 chanx_left_in[0]
port 9 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[10]
port 10 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 chanx_left_in[11]
port 11 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 chanx_left_in[12]
port 12 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 chanx_left_in[13]
port 13 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 chanx_left_in[14]
port 14 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 chanx_left_in[15]
port 15 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[16]
port 16 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[17]
port 17 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[18]
port 18 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 chanx_left_in[19]
port 19 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[1]
port 20 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[2]
port 21 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 chanx_left_in[3]
port 22 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 chanx_left_in[4]
port 23 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 chanx_left_in[5]
port 24 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 chanx_left_in[6]
port 25 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 chanx_left_in[7]
port 26 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[8]
port 27 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[9]
port 28 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 chanx_left_out[0]
port 29 nsew signal output
rlabel metal3 s 0 17552 800 17672 6 chanx_left_out[10]
port 30 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[11]
port 31 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[12]
port 32 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[13]
port 33 nsew signal output
rlabel metal3 s 0 19184 800 19304 6 chanx_left_out[14]
port 34 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 chanx_left_out[15]
port 35 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 chanx_left_out[16]
port 36 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 chanx_left_out[17]
port 37 nsew signal output
rlabel metal3 s 0 20816 800 20936 6 chanx_left_out[18]
port 38 nsew signal output
rlabel metal3 s 0 21224 800 21344 6 chanx_left_out[19]
port 39 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 chanx_left_out[1]
port 40 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 chanx_left_out[2]
port 41 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 chanx_left_out[3]
port 42 nsew signal output
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[4]
port 43 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[5]
port 44 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 chanx_left_out[6]
port 45 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 chanx_left_out[7]
port 46 nsew signal output
rlabel metal3 s 0 16736 800 16856 6 chanx_left_out[8]
port 47 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 chanx_left_out[9]
port 48 nsew signal output
rlabel metal3 s 22200 5312 23000 5432 6 chanx_right_in[0]
port 49 nsew signal input
rlabel metal3 s 22200 9392 23000 9512 6 chanx_right_in[10]
port 50 nsew signal input
rlabel metal3 s 22200 9800 23000 9920 6 chanx_right_in[11]
port 51 nsew signal input
rlabel metal3 s 22200 10208 23000 10328 6 chanx_right_in[12]
port 52 nsew signal input
rlabel metal3 s 22200 10616 23000 10736 6 chanx_right_in[13]
port 53 nsew signal input
rlabel metal3 s 22200 11024 23000 11144 6 chanx_right_in[14]
port 54 nsew signal input
rlabel metal3 s 22200 11432 23000 11552 6 chanx_right_in[15]
port 55 nsew signal input
rlabel metal3 s 22200 11840 23000 11960 6 chanx_right_in[16]
port 56 nsew signal input
rlabel metal3 s 22200 12248 23000 12368 6 chanx_right_in[17]
port 57 nsew signal input
rlabel metal3 s 22200 12656 23000 12776 6 chanx_right_in[18]
port 58 nsew signal input
rlabel metal3 s 22200 13064 23000 13184 6 chanx_right_in[19]
port 59 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 chanx_right_in[1]
port 60 nsew signal input
rlabel metal3 s 22200 6128 23000 6248 6 chanx_right_in[2]
port 61 nsew signal input
rlabel metal3 s 22200 6536 23000 6656 6 chanx_right_in[3]
port 62 nsew signal input
rlabel metal3 s 22200 6944 23000 7064 6 chanx_right_in[4]
port 63 nsew signal input
rlabel metal3 s 22200 7352 23000 7472 6 chanx_right_in[5]
port 64 nsew signal input
rlabel metal3 s 22200 7760 23000 7880 6 chanx_right_in[6]
port 65 nsew signal input
rlabel metal3 s 22200 8168 23000 8288 6 chanx_right_in[7]
port 66 nsew signal input
rlabel metal3 s 22200 8576 23000 8696 6 chanx_right_in[8]
port 67 nsew signal input
rlabel metal3 s 22200 8984 23000 9104 6 chanx_right_in[9]
port 68 nsew signal input
rlabel metal3 s 22200 13472 23000 13592 6 chanx_right_out[0]
port 69 nsew signal output
rlabel metal3 s 22200 17552 23000 17672 6 chanx_right_out[10]
port 70 nsew signal output
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[11]
port 71 nsew signal output
rlabel metal3 s 22200 18368 23000 18488 6 chanx_right_out[12]
port 72 nsew signal output
rlabel metal3 s 22200 18776 23000 18896 6 chanx_right_out[13]
port 73 nsew signal output
rlabel metal3 s 22200 19184 23000 19304 6 chanx_right_out[14]
port 74 nsew signal output
rlabel metal3 s 22200 19592 23000 19712 6 chanx_right_out[15]
port 75 nsew signal output
rlabel metal3 s 22200 20000 23000 20120 6 chanx_right_out[16]
port 76 nsew signal output
rlabel metal3 s 22200 20408 23000 20528 6 chanx_right_out[17]
port 77 nsew signal output
rlabel metal3 s 22200 20816 23000 20936 6 chanx_right_out[18]
port 78 nsew signal output
rlabel metal3 s 22200 21224 23000 21344 6 chanx_right_out[19]
port 79 nsew signal output
rlabel metal3 s 22200 13880 23000 14000 6 chanx_right_out[1]
port 80 nsew signal output
rlabel metal3 s 22200 14288 23000 14408 6 chanx_right_out[2]
port 81 nsew signal output
rlabel metal3 s 22200 14696 23000 14816 6 chanx_right_out[3]
port 82 nsew signal output
rlabel metal3 s 22200 15104 23000 15224 6 chanx_right_out[4]
port 83 nsew signal output
rlabel metal3 s 22200 15512 23000 15632 6 chanx_right_out[5]
port 84 nsew signal output
rlabel metal3 s 22200 15920 23000 16040 6 chanx_right_out[6]
port 85 nsew signal output
rlabel metal3 s 22200 16328 23000 16448 6 chanx_right_out[7]
port 86 nsew signal output
rlabel metal3 s 22200 16736 23000 16856 6 chanx_right_out[8]
port 87 nsew signal output
rlabel metal3 s 22200 17144 23000 17264 6 chanx_right_out[9]
port 88 nsew signal output
rlabel metal2 s 6458 22200 6514 23000 6 chany_top_in[0]
port 89 nsew signal input
rlabel metal2 s 10138 22200 10194 23000 6 chany_top_in[10]
port 90 nsew signal input
rlabel metal2 s 10506 22200 10562 23000 6 chany_top_in[11]
port 91 nsew signal input
rlabel metal2 s 10874 22200 10930 23000 6 chany_top_in[12]
port 92 nsew signal input
rlabel metal2 s 11242 22200 11298 23000 6 chany_top_in[13]
port 93 nsew signal input
rlabel metal2 s 11610 22200 11666 23000 6 chany_top_in[14]
port 94 nsew signal input
rlabel metal2 s 11978 22200 12034 23000 6 chany_top_in[15]
port 95 nsew signal input
rlabel metal2 s 12346 22200 12402 23000 6 chany_top_in[16]
port 96 nsew signal input
rlabel metal2 s 12714 22200 12770 23000 6 chany_top_in[17]
port 97 nsew signal input
rlabel metal2 s 13082 22200 13138 23000 6 chany_top_in[18]
port 98 nsew signal input
rlabel metal2 s 13450 22200 13506 23000 6 chany_top_in[19]
port 99 nsew signal input
rlabel metal2 s 6826 22200 6882 23000 6 chany_top_in[1]
port 100 nsew signal input
rlabel metal2 s 7194 22200 7250 23000 6 chany_top_in[2]
port 101 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[3]
port 102 nsew signal input
rlabel metal2 s 7930 22200 7986 23000 6 chany_top_in[4]
port 103 nsew signal input
rlabel metal2 s 8298 22200 8354 23000 6 chany_top_in[5]
port 104 nsew signal input
rlabel metal2 s 8666 22200 8722 23000 6 chany_top_in[6]
port 105 nsew signal input
rlabel metal2 s 9034 22200 9090 23000 6 chany_top_in[7]
port 106 nsew signal input
rlabel metal2 s 9402 22200 9458 23000 6 chany_top_in[8]
port 107 nsew signal input
rlabel metal2 s 9770 22200 9826 23000 6 chany_top_in[9]
port 108 nsew signal input
rlabel metal2 s 13818 22200 13874 23000 6 chany_top_out[0]
port 109 nsew signal output
rlabel metal2 s 17498 22200 17554 23000 6 chany_top_out[10]
port 110 nsew signal output
rlabel metal2 s 17866 22200 17922 23000 6 chany_top_out[11]
port 111 nsew signal output
rlabel metal2 s 18234 22200 18290 23000 6 chany_top_out[12]
port 112 nsew signal output
rlabel metal2 s 18602 22200 18658 23000 6 chany_top_out[13]
port 113 nsew signal output
rlabel metal2 s 18970 22200 19026 23000 6 chany_top_out[14]
port 114 nsew signal output
rlabel metal2 s 19338 22200 19394 23000 6 chany_top_out[15]
port 115 nsew signal output
rlabel metal2 s 19706 22200 19762 23000 6 chany_top_out[16]
port 116 nsew signal output
rlabel metal2 s 20074 22200 20130 23000 6 chany_top_out[17]
port 117 nsew signal output
rlabel metal2 s 20442 22200 20498 23000 6 chany_top_out[18]
port 118 nsew signal output
rlabel metal2 s 20810 22200 20866 23000 6 chany_top_out[19]
port 119 nsew signal output
rlabel metal2 s 14186 22200 14242 23000 6 chany_top_out[1]
port 120 nsew signal output
rlabel metal2 s 14554 22200 14610 23000 6 chany_top_out[2]
port 121 nsew signal output
rlabel metal2 s 14922 22200 14978 23000 6 chany_top_out[3]
port 122 nsew signal output
rlabel metal2 s 15290 22200 15346 23000 6 chany_top_out[4]
port 123 nsew signal output
rlabel metal2 s 15658 22200 15714 23000 6 chany_top_out[5]
port 124 nsew signal output
rlabel metal2 s 16026 22200 16082 23000 6 chany_top_out[6]
port 125 nsew signal output
rlabel metal2 s 16394 22200 16450 23000 6 chany_top_out[7]
port 126 nsew signal output
rlabel metal2 s 16762 22200 16818 23000 6 chany_top_out[8]
port 127 nsew signal output
rlabel metal2 s 17130 22200 17186 23000 6 chany_top_out[9]
port 128 nsew signal output
rlabel metal2 s 5722 22200 5778 23000 6 clk_3_N_out
port 129 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 clk_3_S_in
port 130 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 left_bottom_grid_pin_11_
port 131 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 left_bottom_grid_pin_13_
port 132 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 left_bottom_grid_pin_15_
port 133 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 left_bottom_grid_pin_17_
port 134 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 left_bottom_grid_pin_1_
port 135 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 left_bottom_grid_pin_3_
port 136 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_5_
port 137 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_7_
port 138 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 left_bottom_grid_pin_9_
port 139 nsew signal input
rlabel metal2 s 4986 22200 5042 23000 6 prog_clk_0_N_in
port 140 nsew signal input
rlabel metal2 s 6090 22200 6146 23000 6 prog_clk_3_N_out
port 141 nsew signal output
rlabel metal2 s 11426 0 11482 800 6 prog_clk_3_S_in
port 142 nsew signal input
rlabel metal3 s 22200 3680 23000 3800 6 right_bottom_grid_pin_11_
port 143 nsew signal input
rlabel metal3 s 22200 4088 23000 4208 6 right_bottom_grid_pin_13_
port 144 nsew signal input
rlabel metal3 s 22200 4496 23000 4616 6 right_bottom_grid_pin_15_
port 145 nsew signal input
rlabel metal3 s 22200 4904 23000 5024 6 right_bottom_grid_pin_17_
port 146 nsew signal input
rlabel metal3 s 22200 1640 23000 1760 6 right_bottom_grid_pin_1_
port 147 nsew signal input
rlabel metal3 s 22200 2048 23000 2168 6 right_bottom_grid_pin_3_
port 148 nsew signal input
rlabel metal3 s 22200 2456 23000 2576 6 right_bottom_grid_pin_5_
port 149 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_7_
port 150 nsew signal input
rlabel metal3 s 22200 3272 23000 3392 6 right_bottom_grid_pin_9_
port 151 nsew signal input
rlabel metal2 s 2042 22200 2098 23000 6 top_left_grid_pin_42_
port 152 nsew signal input
rlabel metal2 s 2410 22200 2466 23000 6 top_left_grid_pin_43_
port 153 nsew signal input
rlabel metal2 s 2778 22200 2834 23000 6 top_left_grid_pin_44_
port 154 nsew signal input
rlabel metal2 s 3146 22200 3202 23000 6 top_left_grid_pin_45_
port 155 nsew signal input
rlabel metal2 s 3514 22200 3570 23000 6 top_left_grid_pin_46_
port 156 nsew signal input
rlabel metal2 s 3882 22200 3938 23000 6 top_left_grid_pin_47_
port 157 nsew signal input
rlabel metal2 s 4250 22200 4306 23000 6 top_left_grid_pin_48_
port 158 nsew signal input
rlabel metal2 s 4618 22200 4674 23000 6 top_left_grid_pin_49_
port 159 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1575782
string GDS_FILE /home/marwan/clear_signoff_final/openlane/sb_1__0_/runs/sb_1__0_/results/signoff/sb_1__0_.magic.gds
string GDS_START 94420
<< end >>

