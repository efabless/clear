magic
tech sky130A
magscale 1 2
timestamp 1656321138
<< obsli1 >>
rect 16140 21123 492932 574005
<< obsm1 >>
rect 7258 5196 501822 574036
<< metal2 >>
rect 15266 576164 15322 576964
rect 33666 576164 33722 576964
rect 52066 576164 52122 576964
rect 70466 576164 70522 576964
rect 88866 576164 88922 576964
rect 107266 576164 107322 576964
rect 125666 576164 125722 576964
rect 144066 576164 144122 576964
rect 162466 576164 162522 576964
rect 180866 576164 180922 576964
rect 199266 576164 199322 576964
rect 217666 576164 217722 576964
rect 236066 576164 236122 576964
rect 254466 576164 254522 576964
rect 272866 576164 272922 576964
rect 291266 576164 291322 576964
rect 309666 576164 309722 576964
rect 328066 576164 328122 576964
rect 346466 576164 346522 576964
rect 364866 576164 364922 576964
rect 383266 576164 383322 576964
rect 401666 576164 401722 576964
rect 420066 576164 420122 576964
rect 438466 576164 438522 576964
rect 456866 576164 456922 576964
rect 475266 576164 475322 576964
rect 493666 576164 493722 576964
rect 7262 3964 7318 4764
rect 9562 3964 9618 4764
rect 11862 3964 11918 4764
rect 14162 3964 14218 4764
rect 16462 3964 16518 4764
rect 18762 3964 18818 4764
rect 21062 3964 21118 4764
rect 23362 3964 23418 4764
rect 25662 3964 25718 4764
rect 27962 3964 28018 4764
rect 30262 3964 30318 4764
rect 32562 3964 32618 4764
rect 34862 3964 34918 4764
rect 37162 3964 37218 4764
rect 39462 3964 39518 4764
rect 41762 3964 41818 4764
rect 44062 3964 44118 4764
rect 46362 3964 46418 4764
rect 48662 3964 48718 4764
rect 50962 3964 51018 4764
rect 53262 3964 53318 4764
rect 55562 3964 55618 4764
rect 57862 3964 57918 4764
rect 60162 3964 60218 4764
rect 62462 3964 62518 4764
rect 64762 3964 64818 4764
rect 67062 3964 67118 4764
rect 69362 3964 69418 4764
rect 71662 3964 71718 4764
rect 73962 3964 74018 4764
rect 76262 3964 76318 4764
rect 78562 3964 78618 4764
rect 80862 3964 80918 4764
rect 83162 3964 83218 4764
rect 85462 3964 85518 4764
rect 87762 3964 87818 4764
rect 90062 3964 90118 4764
rect 92362 3964 92418 4764
rect 94662 3964 94718 4764
rect 96962 3964 97018 4764
rect 99262 3964 99318 4764
rect 101562 3964 101618 4764
rect 103862 3964 103918 4764
rect 106162 3964 106218 4764
rect 108462 3964 108518 4764
rect 110762 3964 110818 4764
rect 113062 3964 113118 4764
rect 115362 3964 115418 4764
rect 117662 3964 117718 4764
rect 119962 3964 120018 4764
rect 122262 3964 122318 4764
rect 124562 3964 124618 4764
rect 126862 3964 126918 4764
rect 129162 3964 129218 4764
rect 131462 3964 131518 4764
rect 133762 3964 133818 4764
rect 136062 3964 136118 4764
rect 138362 3964 138418 4764
rect 140662 3964 140718 4764
rect 142962 3964 143018 4764
rect 145262 3964 145318 4764
rect 147562 3964 147618 4764
rect 149862 3964 149918 4764
rect 152162 3964 152218 4764
rect 154462 3964 154518 4764
rect 156762 3964 156818 4764
rect 159062 3964 159118 4764
rect 161362 3964 161418 4764
rect 163662 3964 163718 4764
rect 165962 3964 166018 4764
rect 168262 3964 168318 4764
rect 170562 3964 170618 4764
rect 172862 3964 172918 4764
rect 175162 3964 175218 4764
rect 177462 3964 177518 4764
rect 179762 3964 179818 4764
rect 182062 3964 182118 4764
rect 184362 3964 184418 4764
rect 186662 3964 186718 4764
rect 188962 3964 189018 4764
rect 191262 3964 191318 4764
rect 193562 3964 193618 4764
rect 195862 3964 195918 4764
rect 198162 3964 198218 4764
rect 200462 3964 200518 4764
rect 202762 3964 202818 4764
rect 205062 3964 205118 4764
rect 207362 3964 207418 4764
rect 209662 3964 209718 4764
rect 211962 3964 212018 4764
rect 214262 3964 214318 4764
rect 216562 3964 216618 4764
rect 218862 3964 218918 4764
rect 221162 3964 221218 4764
rect 223462 3964 223518 4764
rect 225762 3964 225818 4764
rect 228062 3964 228118 4764
rect 230362 3964 230418 4764
rect 232662 3964 232718 4764
rect 234962 3964 235018 4764
rect 237262 3964 237318 4764
rect 239562 3964 239618 4764
rect 241862 3964 241918 4764
rect 244162 3964 244218 4764
rect 246462 3964 246518 4764
rect 248762 3964 248818 4764
rect 251062 3964 251118 4764
rect 253362 3964 253418 4764
rect 255662 3964 255718 4764
rect 257962 3964 258018 4764
rect 260262 3964 260318 4764
rect 262562 3964 262618 4764
rect 264862 3964 264918 4764
rect 267162 3964 267218 4764
rect 269462 3964 269518 4764
rect 271762 3964 271818 4764
rect 274062 3964 274118 4764
rect 276362 3964 276418 4764
rect 278662 3964 278718 4764
rect 280962 3964 281018 4764
rect 283262 3964 283318 4764
rect 285562 3964 285618 4764
rect 287862 3964 287918 4764
rect 290162 3964 290218 4764
rect 292462 3964 292518 4764
rect 294762 3964 294818 4764
rect 297062 3964 297118 4764
rect 299362 3964 299418 4764
rect 301662 3964 301718 4764
rect 303962 3964 304018 4764
rect 306262 3964 306318 4764
rect 308562 3964 308618 4764
rect 310862 3964 310918 4764
rect 313162 3964 313218 4764
rect 315462 3964 315518 4764
rect 317762 3964 317818 4764
rect 320062 3964 320118 4764
rect 322362 3964 322418 4764
rect 324662 3964 324718 4764
rect 326962 3964 327018 4764
rect 329262 3964 329318 4764
rect 331562 3964 331618 4764
rect 333862 3964 333918 4764
rect 336162 3964 336218 4764
rect 338462 3964 338518 4764
rect 340762 3964 340818 4764
rect 343062 3964 343118 4764
rect 345362 3964 345418 4764
rect 347662 3964 347718 4764
rect 349962 3964 350018 4764
rect 352262 3964 352318 4764
rect 354562 3964 354618 4764
rect 356862 3964 356918 4764
rect 359162 3964 359218 4764
rect 361462 3964 361518 4764
rect 363762 3964 363818 4764
rect 366062 3964 366118 4764
rect 368362 3964 368418 4764
rect 370662 3964 370718 4764
rect 372962 3964 373018 4764
rect 375262 3964 375318 4764
rect 377562 3964 377618 4764
rect 379862 3964 379918 4764
rect 382162 3964 382218 4764
rect 384462 3964 384518 4764
rect 386762 3964 386818 4764
rect 389062 3964 389118 4764
rect 391362 3964 391418 4764
rect 393662 3964 393718 4764
rect 395962 3964 396018 4764
rect 398262 3964 398318 4764
rect 400562 3964 400618 4764
rect 402862 3964 402918 4764
rect 405162 3964 405218 4764
rect 407462 3964 407518 4764
rect 409762 3964 409818 4764
rect 412062 3964 412118 4764
rect 414362 3964 414418 4764
rect 416662 3964 416718 4764
rect 418962 3964 419018 4764
rect 421262 3964 421318 4764
rect 423562 3964 423618 4764
rect 425862 3964 425918 4764
rect 428162 3964 428218 4764
rect 430462 3964 430518 4764
rect 432762 3964 432818 4764
rect 435062 3964 435118 4764
rect 437362 3964 437418 4764
rect 439662 3964 439718 4764
rect 441962 3964 442018 4764
rect 444262 3964 444318 4764
rect 446562 3964 446618 4764
rect 448862 3964 448918 4764
rect 451162 3964 451218 4764
rect 453462 3964 453518 4764
rect 455762 3964 455818 4764
rect 458062 3964 458118 4764
rect 460362 3964 460418 4764
rect 462662 3964 462718 4764
rect 464962 3964 465018 4764
rect 467262 3964 467318 4764
rect 469562 3964 469618 4764
rect 471862 3964 471918 4764
rect 474162 3964 474218 4764
rect 476462 3964 476518 4764
rect 478762 3964 478818 4764
rect 481062 3964 481118 4764
rect 483362 3964 483418 4764
rect 485662 3964 485718 4764
rect 487962 3964 488018 4764
rect 490262 3964 490318 4764
rect 492562 3964 492618 4764
rect 494862 3964 494918 4764
rect 497162 3964 497218 4764
rect 499462 3964 499518 4764
rect 501762 3964 501818 4764
<< obsm2 >>
rect 7264 576108 15210 576198
rect 15378 576108 33610 576198
rect 33778 576108 52010 576198
rect 52178 576108 70410 576198
rect 70578 576108 88810 576198
rect 88978 576108 107210 576198
rect 107378 576108 125610 576198
rect 125778 576108 144010 576198
rect 144178 576108 162410 576198
rect 162578 576108 180810 576198
rect 180978 576108 199210 576198
rect 199378 576108 217610 576198
rect 217778 576108 236010 576198
rect 236178 576108 254410 576198
rect 254578 576108 272810 576198
rect 272978 576108 291210 576198
rect 291378 576108 309610 576198
rect 309778 576108 328010 576198
rect 328178 576108 346410 576198
rect 346578 576108 364810 576198
rect 364978 576108 383210 576198
rect 383378 576108 401610 576198
rect 401778 576108 420010 576198
rect 420178 576108 438410 576198
rect 438578 576108 456810 576198
rect 456978 576108 475210 576198
rect 475378 576108 493610 576198
rect 493778 576108 501816 576198
rect 7264 4820 501816 576108
rect 7374 4698 9506 4820
rect 9674 4698 11806 4820
rect 11974 4698 14106 4820
rect 14274 4698 16406 4820
rect 16574 4698 18706 4820
rect 18874 4698 21006 4820
rect 21174 4698 23306 4820
rect 23474 4698 25606 4820
rect 25774 4698 27906 4820
rect 28074 4698 30206 4820
rect 30374 4698 32506 4820
rect 32674 4698 34806 4820
rect 34974 4698 37106 4820
rect 37274 4698 39406 4820
rect 39574 4698 41706 4820
rect 41874 4698 44006 4820
rect 44174 4698 46306 4820
rect 46474 4698 48606 4820
rect 48774 4698 50906 4820
rect 51074 4698 53206 4820
rect 53374 4698 55506 4820
rect 55674 4698 57806 4820
rect 57974 4698 60106 4820
rect 60274 4698 62406 4820
rect 62574 4698 64706 4820
rect 64874 4698 67006 4820
rect 67174 4698 69306 4820
rect 69474 4698 71606 4820
rect 71774 4698 73906 4820
rect 74074 4698 76206 4820
rect 76374 4698 78506 4820
rect 78674 4698 80806 4820
rect 80974 4698 83106 4820
rect 83274 4698 85406 4820
rect 85574 4698 87706 4820
rect 87874 4698 90006 4820
rect 90174 4698 92306 4820
rect 92474 4698 94606 4820
rect 94774 4698 96906 4820
rect 97074 4698 99206 4820
rect 99374 4698 101506 4820
rect 101674 4698 103806 4820
rect 103974 4698 106106 4820
rect 106274 4698 108406 4820
rect 108574 4698 110706 4820
rect 110874 4698 113006 4820
rect 113174 4698 115306 4820
rect 115474 4698 117606 4820
rect 117774 4698 119906 4820
rect 120074 4698 122206 4820
rect 122374 4698 124506 4820
rect 124674 4698 126806 4820
rect 126974 4698 129106 4820
rect 129274 4698 131406 4820
rect 131574 4698 133706 4820
rect 133874 4698 136006 4820
rect 136174 4698 138306 4820
rect 138474 4698 140606 4820
rect 140774 4698 142906 4820
rect 143074 4698 145206 4820
rect 145374 4698 147506 4820
rect 147674 4698 149806 4820
rect 149974 4698 152106 4820
rect 152274 4698 154406 4820
rect 154574 4698 156706 4820
rect 156874 4698 159006 4820
rect 159174 4698 161306 4820
rect 161474 4698 163606 4820
rect 163774 4698 165906 4820
rect 166074 4698 168206 4820
rect 168374 4698 170506 4820
rect 170674 4698 172806 4820
rect 172974 4698 175106 4820
rect 175274 4698 177406 4820
rect 177574 4698 179706 4820
rect 179874 4698 182006 4820
rect 182174 4698 184306 4820
rect 184474 4698 186606 4820
rect 186774 4698 188906 4820
rect 189074 4698 191206 4820
rect 191374 4698 193506 4820
rect 193674 4698 195806 4820
rect 195974 4698 198106 4820
rect 198274 4698 200406 4820
rect 200574 4698 202706 4820
rect 202874 4698 205006 4820
rect 205174 4698 207306 4820
rect 207474 4698 209606 4820
rect 209774 4698 211906 4820
rect 212074 4698 214206 4820
rect 214374 4698 216506 4820
rect 216674 4698 218806 4820
rect 218974 4698 221106 4820
rect 221274 4698 223406 4820
rect 223574 4698 225706 4820
rect 225874 4698 228006 4820
rect 228174 4698 230306 4820
rect 230474 4698 232606 4820
rect 232774 4698 234906 4820
rect 235074 4698 237206 4820
rect 237374 4698 239506 4820
rect 239674 4698 241806 4820
rect 241974 4698 244106 4820
rect 244274 4698 246406 4820
rect 246574 4698 248706 4820
rect 248874 4698 251006 4820
rect 251174 4698 253306 4820
rect 253474 4698 255606 4820
rect 255774 4698 257906 4820
rect 258074 4698 260206 4820
rect 260374 4698 262506 4820
rect 262674 4698 264806 4820
rect 264974 4698 267106 4820
rect 267274 4698 269406 4820
rect 269574 4698 271706 4820
rect 271874 4698 274006 4820
rect 274174 4698 276306 4820
rect 276474 4698 278606 4820
rect 278774 4698 280906 4820
rect 281074 4698 283206 4820
rect 283374 4698 285506 4820
rect 285674 4698 287806 4820
rect 287974 4698 290106 4820
rect 290274 4698 292406 4820
rect 292574 4698 294706 4820
rect 294874 4698 297006 4820
rect 297174 4698 299306 4820
rect 299474 4698 301606 4820
rect 301774 4698 303906 4820
rect 304074 4698 306206 4820
rect 306374 4698 308506 4820
rect 308674 4698 310806 4820
rect 310974 4698 313106 4820
rect 313274 4698 315406 4820
rect 315574 4698 317706 4820
rect 317874 4698 320006 4820
rect 320174 4698 322306 4820
rect 322474 4698 324606 4820
rect 324774 4698 326906 4820
rect 327074 4698 329206 4820
rect 329374 4698 331506 4820
rect 331674 4698 333806 4820
rect 333974 4698 336106 4820
rect 336274 4698 338406 4820
rect 338574 4698 340706 4820
rect 340874 4698 343006 4820
rect 343174 4698 345306 4820
rect 345474 4698 347606 4820
rect 347774 4698 349906 4820
rect 350074 4698 352206 4820
rect 352374 4698 354506 4820
rect 354674 4698 356806 4820
rect 356974 4698 359106 4820
rect 359274 4698 361406 4820
rect 361574 4698 363706 4820
rect 363874 4698 366006 4820
rect 366174 4698 368306 4820
rect 368474 4698 370606 4820
rect 370774 4698 372906 4820
rect 373074 4698 375206 4820
rect 375374 4698 377506 4820
rect 377674 4698 379806 4820
rect 379974 4698 382106 4820
rect 382274 4698 384406 4820
rect 384574 4698 386706 4820
rect 386874 4698 389006 4820
rect 389174 4698 391306 4820
rect 391474 4698 393606 4820
rect 393774 4698 395906 4820
rect 396074 4698 398206 4820
rect 398374 4698 400506 4820
rect 400674 4698 402806 4820
rect 402974 4698 405106 4820
rect 405274 4698 407406 4820
rect 407574 4698 409706 4820
rect 409874 4698 412006 4820
rect 412174 4698 414306 4820
rect 414474 4698 416606 4820
rect 416774 4698 418906 4820
rect 419074 4698 421206 4820
rect 421374 4698 423506 4820
rect 423674 4698 425806 4820
rect 425974 4698 428106 4820
rect 428274 4698 430406 4820
rect 430574 4698 432706 4820
rect 432874 4698 435006 4820
rect 435174 4698 437306 4820
rect 437474 4698 439606 4820
rect 439774 4698 441906 4820
rect 442074 4698 444206 4820
rect 444374 4698 446506 4820
rect 446674 4698 448806 4820
rect 448974 4698 451106 4820
rect 451274 4698 453406 4820
rect 453574 4698 455706 4820
rect 455874 4698 458006 4820
rect 458174 4698 460306 4820
rect 460474 4698 462606 4820
rect 462774 4698 464906 4820
rect 465074 4698 467206 4820
rect 467374 4698 469506 4820
rect 469674 4698 471806 4820
rect 471974 4698 474106 4820
rect 474274 4698 476406 4820
rect 476574 4698 478706 4820
rect 478874 4698 481006 4820
rect 481174 4698 483306 4820
rect 483474 4698 485606 4820
rect 485774 4698 487906 4820
rect 488074 4698 490206 4820
rect 490374 4698 492506 4820
rect 492674 4698 494806 4820
rect 494974 4698 497106 4820
rect 497274 4698 499406 4820
rect 499574 4698 501706 4820
<< metal3 >>
rect 5036 566468 5836 566588
rect 503236 564020 504036 564140
rect 5036 546748 5836 546868
rect 503236 540220 504036 540340
rect 5036 527028 5836 527148
rect 503236 516420 504036 516540
rect 5036 507308 5836 507428
rect 503236 492620 504036 492740
rect 5036 487588 5836 487708
rect 503236 468820 504036 468940
rect 5036 467868 5836 467988
rect 5036 448148 5836 448268
rect 503236 445020 504036 445140
rect 5036 428428 5836 428548
rect 503236 421220 504036 421340
rect 5036 408708 5836 408828
rect 503236 397420 504036 397540
rect 5036 388988 5836 389108
rect 503236 373620 504036 373740
rect 5036 369268 5836 369388
rect 503236 349820 504036 349940
rect 5036 349548 5836 349668
rect 5036 329828 5836 329948
rect 503236 326020 504036 326140
rect 5036 310108 5836 310228
rect 503236 302220 504036 302340
rect 5036 290388 5836 290508
rect 503236 278420 504036 278540
rect 5036 270668 5836 270788
rect 503236 254620 504036 254740
rect 5036 250948 5836 251068
rect 5036 231228 5836 231348
rect 503236 230820 504036 230940
rect 5036 211508 5836 211628
rect 503236 207020 504036 207140
rect 5036 191788 5836 191908
rect 503236 183220 504036 183340
rect 5036 172068 5836 172188
rect 503236 159420 504036 159540
rect 5036 152348 5836 152468
rect 503236 135620 504036 135740
rect 5036 132628 5836 132748
rect 5036 112908 5836 113028
rect 503236 111820 504036 111940
rect 5036 93188 5836 93308
rect 503236 88020 504036 88140
rect 5036 73468 5836 73588
rect 503236 64220 504036 64340
rect 5036 53748 5836 53868
rect 503236 40420 504036 40540
rect 5036 34028 5836 34148
rect 503236 16620 504036 16740
rect 5036 14308 5836 14428
<< obsm3 >>
rect 5836 566668 503236 574021
rect 5916 566388 503236 566668
rect 5836 564220 503236 566388
rect 5836 563940 503156 564220
rect 5836 546948 503236 563940
rect 5916 546668 503236 546948
rect 5836 540420 503236 546668
rect 5836 540140 503156 540420
rect 5836 527228 503236 540140
rect 5916 526948 503236 527228
rect 5836 516620 503236 526948
rect 5836 516340 503156 516620
rect 5836 507508 503236 516340
rect 5916 507228 503236 507508
rect 5836 492820 503236 507228
rect 5836 492540 503156 492820
rect 5836 487788 503236 492540
rect 5916 487508 503236 487788
rect 5836 469020 503236 487508
rect 5836 468740 503156 469020
rect 5836 468068 503236 468740
rect 5916 467788 503236 468068
rect 5836 448348 503236 467788
rect 5916 448068 503236 448348
rect 5836 445220 503236 448068
rect 5836 444940 503156 445220
rect 5836 428628 503236 444940
rect 5916 428348 503236 428628
rect 5836 421420 503236 428348
rect 5836 421140 503156 421420
rect 5836 408908 503236 421140
rect 5916 408628 503236 408908
rect 5836 397620 503236 408628
rect 5836 397340 503156 397620
rect 5836 389188 503236 397340
rect 5916 388908 503236 389188
rect 5836 373820 503236 388908
rect 5836 373540 503156 373820
rect 5836 369468 503236 373540
rect 5916 369188 503236 369468
rect 5836 350020 503236 369188
rect 5836 349748 503156 350020
rect 5916 349740 503156 349748
rect 5916 349468 503236 349740
rect 5836 330028 503236 349468
rect 5916 329748 503236 330028
rect 5836 326220 503236 329748
rect 5836 325940 503156 326220
rect 5836 310308 503236 325940
rect 5916 310028 503236 310308
rect 5836 302420 503236 310028
rect 5836 302140 503156 302420
rect 5836 290588 503236 302140
rect 5916 290308 503236 290588
rect 5836 278620 503236 290308
rect 5836 278340 503156 278620
rect 5836 270868 503236 278340
rect 5916 270588 503236 270868
rect 5836 254820 503236 270588
rect 5836 254540 503156 254820
rect 5836 251148 503236 254540
rect 5916 250868 503236 251148
rect 5836 231428 503236 250868
rect 5916 231148 503236 231428
rect 5836 231020 503236 231148
rect 5836 230740 503156 231020
rect 5836 211708 503236 230740
rect 5916 211428 503236 211708
rect 5836 207220 503236 211428
rect 5836 206940 503156 207220
rect 5836 191988 503236 206940
rect 5916 191708 503236 191988
rect 5836 183420 503236 191708
rect 5836 183140 503156 183420
rect 5836 172268 503236 183140
rect 5916 171988 503236 172268
rect 5836 159620 503236 171988
rect 5836 159340 503156 159620
rect 5836 152548 503236 159340
rect 5916 152268 503236 152548
rect 5836 135820 503236 152268
rect 5836 135540 503156 135820
rect 5836 132828 503236 135540
rect 5916 132548 503236 132828
rect 5836 113108 503236 132548
rect 5916 112828 503236 113108
rect 5836 112020 503236 112828
rect 5836 111740 503156 112020
rect 5836 93388 503236 111740
rect 5916 93108 503236 93388
rect 5836 88220 503236 93108
rect 5836 87940 503156 88220
rect 5836 73668 503236 87940
rect 5916 73388 503236 73668
rect 5836 64420 503236 73388
rect 5836 64140 503156 64420
rect 5836 53948 503236 64140
rect 5916 53668 503236 53948
rect 5836 40620 503236 53668
rect 5836 40340 503156 40620
rect 5836 34228 503236 40340
rect 5916 33948 503236 34228
rect 5836 16820 503236 33948
rect 5836 16540 503156 16820
rect 5836 14508 503236 16540
rect 5916 14335 503236 14508
<< metal4 >>
rect 0 0 900 580760
rect 1240 1240 2140 579520
rect 506848 1240 507748 579520
rect 508088 0 508988 580760
<< obsm4 >>
rect 18579 21092 493092 574036
<< metal5 >>
rect 0 579860 508988 580760
rect 1240 578620 507748 579520
rect 0 572690 508988 573590
rect 0 568190 508988 569090
rect 0 563690 508988 564590
rect 0 559190 508988 560090
rect 0 554690 508988 555590
rect 0 550190 508988 551090
rect 0 545690 508988 546590
rect 0 541190 508988 542090
rect 0 536690 508988 537590
rect 0 532190 508988 533090
rect 0 527690 508988 528590
rect 0 523190 508988 524090
rect 0 518690 508988 519590
rect 0 514190 508988 515090
rect 0 509690 508988 510590
rect 0 505190 508988 506090
rect 0 500690 508988 501590
rect 0 496190 508988 497090
rect 0 491690 508988 492590
rect 0 487190 508988 488090
rect 0 482690 508988 483590
rect 0 478190 508988 479090
rect 0 473690 508988 474590
rect 0 469190 508988 470090
rect 0 464690 508988 465590
rect 0 460190 508988 461090
rect 0 455690 508988 456590
rect 0 451190 508988 452090
rect 0 446690 508988 447590
rect 0 442190 508988 443090
rect 0 437690 508988 438590
rect 0 433190 508988 434090
rect 0 428690 508988 429590
rect 0 424190 508988 425090
rect 0 419690 508988 420590
rect 0 415190 508988 416090
rect 0 410690 508988 411590
rect 0 406190 508988 407090
rect 0 401690 508988 402590
rect 0 397190 508988 398090
rect 0 392690 508988 393590
rect 0 388190 508988 389090
rect 0 383690 508988 384590
rect 0 379190 508988 380090
rect 0 374690 508988 375590
rect 0 370190 508988 371090
rect 0 365690 508988 366590
rect 0 361190 508988 362090
rect 0 356690 508988 357590
rect 0 352190 508988 353090
rect 0 347690 508988 348590
rect 0 343190 508988 344090
rect 0 338690 508988 339590
rect 0 334190 508988 335090
rect 0 329690 508988 330590
rect 0 325190 508988 326090
rect 0 320690 508988 321590
rect 0 316190 508988 317090
rect 0 311690 508988 312590
rect 0 307190 508988 308090
rect 0 302690 508988 303590
rect 0 298190 508988 299090
rect 0 293690 508988 294590
rect 0 289190 508988 290090
rect 0 284690 508988 285590
rect 0 280190 508988 281090
rect 0 275690 508988 276590
rect 0 271190 508988 272090
rect 0 266690 508988 267590
rect 0 262190 508988 263090
rect 0 257690 508988 258590
rect 0 253190 508988 254090
rect 0 248690 508988 249590
rect 0 244190 508988 245090
rect 0 239690 508988 240590
rect 0 235190 508988 236090
rect 0 230690 508988 231590
rect 0 226190 508988 227090
rect 0 221690 508988 222590
rect 0 217190 508988 218090
rect 0 212690 508988 213590
rect 0 208190 508988 209090
rect 0 203690 508988 204590
rect 0 199190 508988 200090
rect 0 194690 508988 195590
rect 0 190190 508988 191090
rect 0 185690 508988 186590
rect 0 181190 508988 182090
rect 0 176690 508988 177590
rect 0 172190 508988 173090
rect 0 167690 508988 168590
rect 0 163190 508988 164090
rect 0 158690 508988 159590
rect 0 154190 508988 155090
rect 0 149690 508988 150590
rect 0 145190 508988 146090
rect 0 140690 508988 141590
rect 0 136190 508988 137090
rect 0 131690 508988 132590
rect 0 127190 508988 128090
rect 0 122690 508988 123590
rect 0 118190 508988 119090
rect 0 113690 508988 114590
rect 0 109190 508988 110090
rect 0 104690 508988 105590
rect 0 100190 508988 101090
rect 0 95690 508988 96590
rect 0 91190 508988 92090
rect 0 86690 508988 87590
rect 0 82190 508988 83090
rect 0 77690 508988 78590
rect 0 73190 508988 74090
rect 0 68690 508988 69590
rect 0 64190 508988 65090
rect 0 59690 508988 60590
rect 0 55190 508988 56090
rect 0 50690 508988 51590
rect 0 46190 508988 47090
rect 0 41690 508988 42590
rect 0 37190 508988 38090
rect 0 32690 508988 33590
rect 0 28190 508988 29090
rect 0 23690 508988 24590
rect 1240 1240 507748 2140
rect 0 0 508988 900
<< labels >>
rlabel metal3 s 5036 73468 5836 73588 6 IO_ISOL_N
port 1 nsew signal input
rlabel metal3 s 5036 34028 5836 34148 6 Test_en
port 2 nsew signal input
rlabel metal4 s 0 0 900 580760 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 0 508988 900 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 579860 508988 580760 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 508088 0 508988 580760 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 28190 508988 29090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 37190 508988 38090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 46190 508988 47090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 55190 508988 56090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 64190 508988 65090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 73190 508988 74090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 82190 508988 83090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 91190 508988 92090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 100190 508988 101090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 109190 508988 110090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 118190 508988 119090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 127190 508988 128090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 136190 508988 137090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 145190 508988 146090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 154190 508988 155090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 163190 508988 164090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 172190 508988 173090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 181190 508988 182090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 190190 508988 191090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 199190 508988 200090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 208190 508988 209090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 217190 508988 218090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 226190 508988 227090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 235190 508988 236090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 244190 508988 245090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 253190 508988 254090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 262190 508988 263090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 271190 508988 272090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 280190 508988 281090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 289190 508988 290090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 298190 508988 299090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 307190 508988 308090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 316190 508988 317090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 325190 508988 326090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 334190 508988 335090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 343190 508988 344090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 352190 508988 353090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 361190 508988 362090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 370190 508988 371090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 379190 508988 380090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 388190 508988 389090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 397190 508988 398090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 406190 508988 407090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 415190 508988 416090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 424190 508988 425090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 433190 508988 434090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 442190 508988 443090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 451190 508988 452090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 460190 508988 461090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 469190 508988 470090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 478190 508988 479090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 487190 508988 488090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 496190 508988 497090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 505190 508988 506090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 514190 508988 515090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 523190 508988 524090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 532190 508988 533090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 541190 508988 542090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 550190 508988 551090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 559190 508988 560090 6 VGND
port 3 nsew ground bidirectional
rlabel metal5 s 0 568190 508988 569090 6 VGND
port 3 nsew ground bidirectional
rlabel metal4 s 1240 1240 2140 579520 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 1240 1240 507748 2140 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 1240 578620 507748 579520 6 VPWR
port 4 nsew power bidirectional
rlabel metal4 s 506848 1240 507748 579520 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 23690 508988 24590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 32690 508988 33590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 41690 508988 42590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 50690 508988 51590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 59690 508988 60590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 68690 508988 69590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 77690 508988 78590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 86690 508988 87590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 95690 508988 96590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 104690 508988 105590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 113690 508988 114590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 122690 508988 123590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 131690 508988 132590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 140690 508988 141590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 149690 508988 150590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 158690 508988 159590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 167690 508988 168590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 176690 508988 177590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 185690 508988 186590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 194690 508988 195590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 203690 508988 204590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 212690 508988 213590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 221690 508988 222590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 230690 508988 231590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 239690 508988 240590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 248690 508988 249590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 257690 508988 258590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 266690 508988 267590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 275690 508988 276590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 284690 508988 285590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 293690 508988 294590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 302690 508988 303590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 311690 508988 312590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 320690 508988 321590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 329690 508988 330590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 338690 508988 339590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 347690 508988 348590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 356690 508988 357590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 365690 508988 366590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 374690 508988 375590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 383690 508988 384590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 392690 508988 393590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 401690 508988 402590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 410690 508988 411590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 419690 508988 420590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 428690 508988 429590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 437690 508988 438590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 446690 508988 447590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 455690 508988 456590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 464690 508988 465590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 473690 508988 474590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 482690 508988 483590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 491690 508988 492590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 500690 508988 501590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 509690 508988 510590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 518690 508988 519590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 527690 508988 528590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 536690 508988 537590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 545690 508988 546590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 554690 508988 555590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 563690 508988 564590 6 VPWR
port 4 nsew power bidirectional
rlabel metal5 s 0 572690 508988 573590 6 VPWR
port 4 nsew power bidirectional
rlabel metal3 s 503236 540220 504036 540340 6 ccff_head
port 5 nsew signal input
rlabel metal3 s 5036 14308 5836 14428 6 ccff_tail
port 6 nsew signal output
rlabel metal3 s 5036 53748 5836 53868 6 clk
port 7 nsew signal input
rlabel metal2 s 15266 576164 15322 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
port 8 nsew signal output
rlabel metal3 s 503236 111820 504036 111940 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[10]
port 9 nsew signal output
rlabel metal3 s 503236 183220 504036 183340 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[11]
port 10 nsew signal output
rlabel metal3 s 503236 254620 504036 254740 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[12]
port 11 nsew signal output
rlabel metal3 s 503236 326020 504036 326140 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[13]
port 12 nsew signal output
rlabel metal3 s 503236 397420 504036 397540 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[14]
port 13 nsew signal output
rlabel metal3 s 503236 468820 504036 468940 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[15]
port 14 nsew signal output
rlabel metal2 s 441962 3964 442018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[16]
port 15 nsew signal output
rlabel metal2 s 444262 3964 444318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[17]
port 16 nsew signal output
rlabel metal2 s 446562 3964 446618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[18]
port 17 nsew signal output
rlabel metal2 s 448862 3964 448918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[19]
port 18 nsew signal output
rlabel metal2 s 33666 576164 33722 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
port 19 nsew signal output
rlabel metal2 s 451162 3964 451218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[20]
port 20 nsew signal output
rlabel metal2 s 453462 3964 453518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[21]
port 21 nsew signal output
rlabel metal2 s 455762 3964 455818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[22]
port 22 nsew signal output
rlabel metal2 s 458062 3964 458118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[23]
port 23 nsew signal output
rlabel metal2 s 460362 3964 460418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[24]
port 24 nsew signal output
rlabel metal2 s 379862 3964 379918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[25]
port 25 nsew signal output
rlabel metal2 s 382162 3964 382218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[26]
port 26 nsew signal output
rlabel metal2 s 384462 3964 384518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[27]
port 27 nsew signal output
rlabel metal2 s 386762 3964 386818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[28]
port 28 nsew signal output
rlabel metal2 s 389062 3964 389118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[29]
port 29 nsew signal output
rlabel metal2 s 52066 576164 52122 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
port 30 nsew signal output
rlabel metal2 s 391362 3964 391418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[30]
port 31 nsew signal output
rlabel metal2 s 393662 3964 393718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[31]
port 32 nsew signal output
rlabel metal2 s 395962 3964 396018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[32]
port 33 nsew signal output
rlabel metal2 s 398262 3964 398318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[33]
port 34 nsew signal output
rlabel metal2 s 317762 3964 317818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[34]
port 35 nsew signal output
rlabel metal2 s 320062 3964 320118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[35]
port 36 nsew signal output
rlabel metal2 s 322362 3964 322418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[36]
port 37 nsew signal output
rlabel metal2 s 324662 3964 324718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[37]
port 38 nsew signal output
rlabel metal2 s 326962 3964 327018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[38]
port 39 nsew signal output
rlabel metal2 s 329262 3964 329318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[39]
port 40 nsew signal output
rlabel metal2 s 70466 576164 70522 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
port 41 nsew signal output
rlabel metal2 s 331562 3964 331618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[40]
port 42 nsew signal output
rlabel metal2 s 333862 3964 333918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[41]
port 43 nsew signal output
rlabel metal2 s 336162 3964 336218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[42]
port 44 nsew signal output
rlabel metal2 s 255662 3964 255718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[43]
port 45 nsew signal output
rlabel metal2 s 257962 3964 258018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[44]
port 46 nsew signal output
rlabel metal2 s 260262 3964 260318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[45]
port 47 nsew signal output
rlabel metal2 s 262562 3964 262618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[46]
port 48 nsew signal output
rlabel metal2 s 264862 3964 264918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[47]
port 49 nsew signal output
rlabel metal2 s 267162 3964 267218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[48]
port 50 nsew signal output
rlabel metal2 s 269462 3964 269518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[49]
port 51 nsew signal output
rlabel metal2 s 88866 576164 88922 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
port 52 nsew signal output
rlabel metal2 s 271762 3964 271818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[50]
port 53 nsew signal output
rlabel metal2 s 274062 3964 274118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[51]
port 54 nsew signal output
rlabel metal2 s 193562 3964 193618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[52]
port 55 nsew signal output
rlabel metal2 s 195862 3964 195918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[53]
port 56 nsew signal output
rlabel metal2 s 198162 3964 198218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[54]
port 57 nsew signal output
rlabel metal2 s 200462 3964 200518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[55]
port 58 nsew signal output
rlabel metal2 s 202762 3964 202818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[56]
port 59 nsew signal output
rlabel metal2 s 205062 3964 205118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[57]
port 60 nsew signal output
rlabel metal2 s 207362 3964 207418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[58]
port 61 nsew signal output
rlabel metal2 s 209662 3964 209718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[59]
port 62 nsew signal output
rlabel metal2 s 107266 576164 107322 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
port 63 nsew signal output
rlabel metal2 s 211962 3964 212018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[60]
port 64 nsew signal output
rlabel metal2 s 131462 3964 131518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[61]
port 65 nsew signal output
rlabel metal2 s 133762 3964 133818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[62]
port 66 nsew signal output
rlabel metal2 s 136062 3964 136118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[63]
port 67 nsew signal output
rlabel metal2 s 138362 3964 138418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[64]
port 68 nsew signal output
rlabel metal2 s 140662 3964 140718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[65]
port 69 nsew signal output
rlabel metal2 s 142962 3964 143018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[66]
port 70 nsew signal output
rlabel metal2 s 145262 3964 145318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[67]
port 71 nsew signal output
rlabel metal2 s 147562 3964 147618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[68]
port 72 nsew signal output
rlabel metal2 s 149862 3964 149918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[69]
port 73 nsew signal output
rlabel metal2 s 125666 576164 125722 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
port 74 nsew signal output
rlabel metal2 s 69362 3964 69418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[70]
port 75 nsew signal output
rlabel metal2 s 71662 3964 71718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[71]
port 76 nsew signal output
rlabel metal2 s 73962 3964 74018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[72]
port 77 nsew signal output
rlabel metal2 s 76262 3964 76318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[73]
port 78 nsew signal output
rlabel metal2 s 78562 3964 78618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[74]
port 79 nsew signal output
rlabel metal2 s 80862 3964 80918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[75]
port 80 nsew signal output
rlabel metal2 s 83162 3964 83218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[76]
port 81 nsew signal output
rlabel metal2 s 85462 3964 85518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[77]
port 82 nsew signal output
rlabel metal2 s 87762 3964 87818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[78]
port 83 nsew signal output
rlabel metal2 s 7262 3964 7318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[79]
port 84 nsew signal output
rlabel metal2 s 144066 576164 144122 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
port 85 nsew signal output
rlabel metal2 s 9562 3964 9618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[80]
port 86 nsew signal output
rlabel metal2 s 11862 3964 11918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[81]
port 87 nsew signal output
rlabel metal2 s 14162 3964 14218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[82]
port 88 nsew signal output
rlabel metal2 s 16462 3964 16518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[83]
port 89 nsew signal output
rlabel metal2 s 18762 3964 18818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[84]
port 90 nsew signal output
rlabel metal2 s 21062 3964 21118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[85]
port 91 nsew signal output
rlabel metal2 s 23362 3964 23418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[86]
port 92 nsew signal output
rlabel metal2 s 25662 3964 25718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[87]
port 93 nsew signal output
rlabel metal3 s 5036 93188 5836 93308 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[88]
port 94 nsew signal output
rlabel metal3 s 5036 152348 5836 152468 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[89]
port 95 nsew signal output
rlabel metal2 s 162466 576164 162522 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
port 96 nsew signal output
rlabel metal3 s 5036 211508 5836 211628 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[90]
port 97 nsew signal output
rlabel metal3 s 5036 270668 5836 270788 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[91]
port 98 nsew signal output
rlabel metal3 s 5036 329828 5836 329948 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[92]
port 99 nsew signal output
rlabel metal3 s 5036 388988 5836 389108 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[93]
port 100 nsew signal output
rlabel metal3 s 5036 448148 5836 448268 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[94]
port 101 nsew signal output
rlabel metal3 s 5036 507308 5836 507428 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[95]
port 102 nsew signal output
rlabel metal3 s 503236 40420 504036 40540 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[9]
port 103 nsew signal output
rlabel metal2 s 180866 576164 180922 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
port 104 nsew signal input
rlabel metal3 s 503236 135620 504036 135740 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[10]
port 105 nsew signal input
rlabel metal3 s 503236 207020 504036 207140 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[11]
port 106 nsew signal input
rlabel metal3 s 503236 278420 504036 278540 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[12]
port 107 nsew signal input
rlabel metal3 s 503236 349820 504036 349940 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[13]
port 108 nsew signal input
rlabel metal3 s 503236 421220 504036 421340 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[14]
port 109 nsew signal input
rlabel metal3 s 503236 492620 504036 492740 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[15]
port 110 nsew signal input
rlabel metal2 s 462662 3964 462718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[16]
port 111 nsew signal input
rlabel metal2 s 464962 3964 465018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[17]
port 112 nsew signal input
rlabel metal2 s 467262 3964 467318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[18]
port 113 nsew signal input
rlabel metal2 s 469562 3964 469618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[19]
port 114 nsew signal input
rlabel metal2 s 199266 576164 199322 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
port 115 nsew signal input
rlabel metal2 s 471862 3964 471918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[20]
port 116 nsew signal input
rlabel metal2 s 474162 3964 474218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[21]
port 117 nsew signal input
rlabel metal2 s 476462 3964 476518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[22]
port 118 nsew signal input
rlabel metal2 s 478762 3964 478818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[23]
port 119 nsew signal input
rlabel metal2 s 481062 3964 481118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[24]
port 120 nsew signal input
rlabel metal2 s 400562 3964 400618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[25]
port 121 nsew signal input
rlabel metal2 s 402862 3964 402918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[26]
port 122 nsew signal input
rlabel metal2 s 405162 3964 405218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[27]
port 123 nsew signal input
rlabel metal2 s 407462 3964 407518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[28]
port 124 nsew signal input
rlabel metal2 s 409762 3964 409818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[29]
port 125 nsew signal input
rlabel metal2 s 217666 576164 217722 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
port 126 nsew signal input
rlabel metal2 s 412062 3964 412118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[30]
port 127 nsew signal input
rlabel metal2 s 414362 3964 414418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[31]
port 128 nsew signal input
rlabel metal2 s 416662 3964 416718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[32]
port 129 nsew signal input
rlabel metal2 s 418962 3964 419018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[33]
port 130 nsew signal input
rlabel metal2 s 338462 3964 338518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[34]
port 131 nsew signal input
rlabel metal2 s 340762 3964 340818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[35]
port 132 nsew signal input
rlabel metal2 s 343062 3964 343118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[36]
port 133 nsew signal input
rlabel metal2 s 345362 3964 345418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[37]
port 134 nsew signal input
rlabel metal2 s 347662 3964 347718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[38]
port 135 nsew signal input
rlabel metal2 s 349962 3964 350018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[39]
port 136 nsew signal input
rlabel metal2 s 236066 576164 236122 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
port 137 nsew signal input
rlabel metal2 s 352262 3964 352318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[40]
port 138 nsew signal input
rlabel metal2 s 354562 3964 354618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[41]
port 139 nsew signal input
rlabel metal2 s 356862 3964 356918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[42]
port 140 nsew signal input
rlabel metal2 s 276362 3964 276418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[43]
port 141 nsew signal input
rlabel metal2 s 278662 3964 278718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[44]
port 142 nsew signal input
rlabel metal2 s 280962 3964 281018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[45]
port 143 nsew signal input
rlabel metal2 s 283262 3964 283318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[46]
port 144 nsew signal input
rlabel metal2 s 285562 3964 285618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[47]
port 145 nsew signal input
rlabel metal2 s 287862 3964 287918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[48]
port 146 nsew signal input
rlabel metal2 s 290162 3964 290218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[49]
port 147 nsew signal input
rlabel metal2 s 254466 576164 254522 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
port 148 nsew signal input
rlabel metal2 s 292462 3964 292518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[50]
port 149 nsew signal input
rlabel metal2 s 294762 3964 294818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[51]
port 150 nsew signal input
rlabel metal2 s 214262 3964 214318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[52]
port 151 nsew signal input
rlabel metal2 s 216562 3964 216618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[53]
port 152 nsew signal input
rlabel metal2 s 218862 3964 218918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[54]
port 153 nsew signal input
rlabel metal2 s 221162 3964 221218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[55]
port 154 nsew signal input
rlabel metal2 s 223462 3964 223518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[56]
port 155 nsew signal input
rlabel metal2 s 225762 3964 225818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[57]
port 156 nsew signal input
rlabel metal2 s 228062 3964 228118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[58]
port 157 nsew signal input
rlabel metal2 s 230362 3964 230418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[59]
port 158 nsew signal input
rlabel metal2 s 272866 576164 272922 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
port 159 nsew signal input
rlabel metal2 s 232662 3964 232718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[60]
port 160 nsew signal input
rlabel metal2 s 152162 3964 152218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[61]
port 161 nsew signal input
rlabel metal2 s 154462 3964 154518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[62]
port 162 nsew signal input
rlabel metal2 s 156762 3964 156818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[63]
port 163 nsew signal input
rlabel metal2 s 159062 3964 159118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[64]
port 164 nsew signal input
rlabel metal2 s 161362 3964 161418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[65]
port 165 nsew signal input
rlabel metal2 s 163662 3964 163718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[66]
port 166 nsew signal input
rlabel metal2 s 165962 3964 166018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[67]
port 167 nsew signal input
rlabel metal2 s 168262 3964 168318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[68]
port 168 nsew signal input
rlabel metal2 s 170562 3964 170618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[69]
port 169 nsew signal input
rlabel metal2 s 291266 576164 291322 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
port 170 nsew signal input
rlabel metal2 s 90062 3964 90118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[70]
port 171 nsew signal input
rlabel metal2 s 92362 3964 92418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[71]
port 172 nsew signal input
rlabel metal2 s 94662 3964 94718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[72]
port 173 nsew signal input
rlabel metal2 s 96962 3964 97018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[73]
port 174 nsew signal input
rlabel metal2 s 99262 3964 99318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[74]
port 175 nsew signal input
rlabel metal2 s 101562 3964 101618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[75]
port 176 nsew signal input
rlabel metal2 s 103862 3964 103918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[76]
port 177 nsew signal input
rlabel metal2 s 106162 3964 106218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[77]
port 178 nsew signal input
rlabel metal2 s 108462 3964 108518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[78]
port 179 nsew signal input
rlabel metal2 s 27962 3964 28018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[79]
port 180 nsew signal input
rlabel metal2 s 309666 576164 309722 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
port 181 nsew signal input
rlabel metal2 s 30262 3964 30318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[80]
port 182 nsew signal input
rlabel metal2 s 32562 3964 32618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[81]
port 183 nsew signal input
rlabel metal2 s 34862 3964 34918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[82]
port 184 nsew signal input
rlabel metal2 s 37162 3964 37218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[83]
port 185 nsew signal input
rlabel metal2 s 39462 3964 39518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[84]
port 186 nsew signal input
rlabel metal2 s 41762 3964 41818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[85]
port 187 nsew signal input
rlabel metal2 s 44062 3964 44118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[86]
port 188 nsew signal input
rlabel metal2 s 46362 3964 46418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[87]
port 189 nsew signal input
rlabel metal3 s 5036 112908 5836 113028 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[88]
port 190 nsew signal input
rlabel metal3 s 5036 172068 5836 172188 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[89]
port 191 nsew signal input
rlabel metal2 s 328066 576164 328122 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
port 192 nsew signal input
rlabel metal3 s 5036 231228 5836 231348 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[90]
port 193 nsew signal input
rlabel metal3 s 5036 290388 5836 290508 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[91]
port 194 nsew signal input
rlabel metal3 s 5036 349548 5836 349668 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[92]
port 195 nsew signal input
rlabel metal3 s 5036 408708 5836 408828 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[93]
port 196 nsew signal input
rlabel metal3 s 5036 467868 5836 467988 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[94]
port 197 nsew signal input
rlabel metal3 s 5036 527028 5836 527148 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[95]
port 198 nsew signal input
rlabel metal3 s 503236 64220 504036 64340 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[9]
port 199 nsew signal input
rlabel metal2 s 346466 576164 346522 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
port 200 nsew signal output
rlabel metal3 s 503236 159420 504036 159540 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[10]
port 201 nsew signal output
rlabel metal3 s 503236 230820 504036 230940 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[11]
port 202 nsew signal output
rlabel metal3 s 503236 302220 504036 302340 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[12]
port 203 nsew signal output
rlabel metal3 s 503236 373620 504036 373740 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[13]
port 204 nsew signal output
rlabel metal3 s 503236 445020 504036 445140 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[14]
port 205 nsew signal output
rlabel metal3 s 503236 516420 504036 516540 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[15]
port 206 nsew signal output
rlabel metal2 s 483362 3964 483418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[16]
port 207 nsew signal output
rlabel metal2 s 485662 3964 485718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[17]
port 208 nsew signal output
rlabel metal2 s 487962 3964 488018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[18]
port 209 nsew signal output
rlabel metal2 s 490262 3964 490318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[19]
port 210 nsew signal output
rlabel metal2 s 364866 576164 364922 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
port 211 nsew signal output
rlabel metal2 s 492562 3964 492618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[20]
port 212 nsew signal output
rlabel metal2 s 494862 3964 494918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[21]
port 213 nsew signal output
rlabel metal2 s 497162 3964 497218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[22]
port 214 nsew signal output
rlabel metal2 s 499462 3964 499518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[23]
port 215 nsew signal output
rlabel metal2 s 501762 3964 501818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[24]
port 216 nsew signal output
rlabel metal2 s 421262 3964 421318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[25]
port 217 nsew signal output
rlabel metal2 s 423562 3964 423618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[26]
port 218 nsew signal output
rlabel metal2 s 425862 3964 425918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[27]
port 219 nsew signal output
rlabel metal2 s 428162 3964 428218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[28]
port 220 nsew signal output
rlabel metal2 s 430462 3964 430518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[29]
port 221 nsew signal output
rlabel metal2 s 383266 576164 383322 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
port 222 nsew signal output
rlabel metal2 s 432762 3964 432818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[30]
port 223 nsew signal output
rlabel metal2 s 435062 3964 435118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[31]
port 224 nsew signal output
rlabel metal2 s 437362 3964 437418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[32]
port 225 nsew signal output
rlabel metal2 s 439662 3964 439718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[33]
port 226 nsew signal output
rlabel metal2 s 359162 3964 359218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[34]
port 227 nsew signal output
rlabel metal2 s 361462 3964 361518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[35]
port 228 nsew signal output
rlabel metal2 s 363762 3964 363818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[36]
port 229 nsew signal output
rlabel metal2 s 366062 3964 366118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[37]
port 230 nsew signal output
rlabel metal2 s 368362 3964 368418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[38]
port 231 nsew signal output
rlabel metal2 s 370662 3964 370718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[39]
port 232 nsew signal output
rlabel metal2 s 401666 576164 401722 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
port 233 nsew signal output
rlabel metal2 s 372962 3964 373018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[40]
port 234 nsew signal output
rlabel metal2 s 375262 3964 375318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[41]
port 235 nsew signal output
rlabel metal2 s 377562 3964 377618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[42]
port 236 nsew signal output
rlabel metal2 s 297062 3964 297118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[43]
port 237 nsew signal output
rlabel metal2 s 299362 3964 299418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[44]
port 238 nsew signal output
rlabel metal2 s 301662 3964 301718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[45]
port 239 nsew signal output
rlabel metal2 s 303962 3964 304018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[46]
port 240 nsew signal output
rlabel metal2 s 306262 3964 306318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[47]
port 241 nsew signal output
rlabel metal2 s 308562 3964 308618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[48]
port 242 nsew signal output
rlabel metal2 s 310862 3964 310918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[49]
port 243 nsew signal output
rlabel metal2 s 420066 576164 420122 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
port 244 nsew signal output
rlabel metal2 s 313162 3964 313218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[50]
port 245 nsew signal output
rlabel metal2 s 315462 3964 315518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[51]
port 246 nsew signal output
rlabel metal2 s 234962 3964 235018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[52]
port 247 nsew signal output
rlabel metal2 s 237262 3964 237318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[53]
port 248 nsew signal output
rlabel metal2 s 239562 3964 239618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[54]
port 249 nsew signal output
rlabel metal2 s 241862 3964 241918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[55]
port 250 nsew signal output
rlabel metal2 s 244162 3964 244218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[56]
port 251 nsew signal output
rlabel metal2 s 246462 3964 246518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[57]
port 252 nsew signal output
rlabel metal2 s 248762 3964 248818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[58]
port 253 nsew signal output
rlabel metal2 s 251062 3964 251118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[59]
port 254 nsew signal output
rlabel metal2 s 438466 576164 438522 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
port 255 nsew signal output
rlabel metal2 s 253362 3964 253418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[60]
port 256 nsew signal output
rlabel metal2 s 172862 3964 172918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[61]
port 257 nsew signal output
rlabel metal2 s 175162 3964 175218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[62]
port 258 nsew signal output
rlabel metal2 s 177462 3964 177518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[63]
port 259 nsew signal output
rlabel metal2 s 179762 3964 179818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[64]
port 260 nsew signal output
rlabel metal2 s 182062 3964 182118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[65]
port 261 nsew signal output
rlabel metal2 s 184362 3964 184418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[66]
port 262 nsew signal output
rlabel metal2 s 186662 3964 186718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[67]
port 263 nsew signal output
rlabel metal2 s 188962 3964 189018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[68]
port 264 nsew signal output
rlabel metal2 s 191262 3964 191318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[69]
port 265 nsew signal output
rlabel metal2 s 456866 576164 456922 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
port 266 nsew signal output
rlabel metal2 s 110762 3964 110818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[70]
port 267 nsew signal output
rlabel metal2 s 113062 3964 113118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[71]
port 268 nsew signal output
rlabel metal2 s 115362 3964 115418 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[72]
port 269 nsew signal output
rlabel metal2 s 117662 3964 117718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[73]
port 270 nsew signal output
rlabel metal2 s 119962 3964 120018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[74]
port 271 nsew signal output
rlabel metal2 s 122262 3964 122318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[75]
port 272 nsew signal output
rlabel metal2 s 124562 3964 124618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[76]
port 273 nsew signal output
rlabel metal2 s 126862 3964 126918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[77]
port 274 nsew signal output
rlabel metal2 s 129162 3964 129218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[78]
port 275 nsew signal output
rlabel metal2 s 48662 3964 48718 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[79]
port 276 nsew signal output
rlabel metal2 s 475266 576164 475322 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
port 277 nsew signal output
rlabel metal2 s 50962 3964 51018 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[80]
port 278 nsew signal output
rlabel metal2 s 53262 3964 53318 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[81]
port 279 nsew signal output
rlabel metal2 s 55562 3964 55618 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[82]
port 280 nsew signal output
rlabel metal2 s 57862 3964 57918 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[83]
port 281 nsew signal output
rlabel metal2 s 60162 3964 60218 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[84]
port 282 nsew signal output
rlabel metal2 s 62462 3964 62518 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[85]
port 283 nsew signal output
rlabel metal2 s 64762 3964 64818 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[86]
port 284 nsew signal output
rlabel metal2 s 67062 3964 67118 4764 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[87]
port 285 nsew signal output
rlabel metal3 s 5036 132628 5836 132748 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[88]
port 286 nsew signal output
rlabel metal3 s 5036 191788 5836 191908 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[89]
port 287 nsew signal output
rlabel metal2 s 493666 576164 493722 576964 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
port 288 nsew signal output
rlabel metal3 s 5036 250948 5836 251068 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[90]
port 289 nsew signal output
rlabel metal3 s 5036 310108 5836 310228 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[91]
port 290 nsew signal output
rlabel metal3 s 5036 369268 5836 369388 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[92]
port 291 nsew signal output
rlabel metal3 s 5036 428428 5836 428548 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[93]
port 292 nsew signal output
rlabel metal3 s 5036 487588 5836 487708 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[94]
port 293 nsew signal output
rlabel metal3 s 5036 546748 5836 546868 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[95]
port 294 nsew signal output
rlabel metal3 s 503236 88020 504036 88140 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[9]
port 295 nsew signal output
rlabel metal3 s 503236 16620 504036 16740 6 prog_clk
port 296 nsew signal input
rlabel metal3 s 5036 566468 5836 566588 6 sc_head
port 297 nsew signal input
rlabel metal3 s 503236 564020 504036 564140 6 sc_tail
port 298 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 508988 580760
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 39104070
string GDS_FILE /home/marwan/clear_signoff_final/openlane/fpga_core/runs/fpga_core/results/signoff/fpga_core.magic.gds
string GDS_START 21725804
<< end >>

