magic
tech sky130A
magscale 1 2
timestamp 1681685900
<< obsli1 >>
rect 368 2159 494592 540753
<< obsm1 >>
rect 368 1368 494592 540784
<< metal2 >>
rect 6734 542200 6790 543000
rect 11150 542200 11206 543000
rect 15566 542200 15622 543000
rect 19982 542200 20038 543000
rect 24398 542200 24454 543000
rect 28814 542200 28870 543000
rect 33230 542200 33286 543000
rect 37646 542200 37702 543000
rect 42062 542200 42118 543000
rect 46478 542200 46534 543000
rect 50894 542200 50950 543000
rect 55310 542200 55366 543000
rect 59726 542200 59782 543000
rect 64142 542200 64198 543000
rect 68558 542200 68614 543000
rect 72974 542200 73030 543000
rect 77390 542200 77446 543000
rect 81806 542200 81862 543000
rect 86222 542200 86278 543000
rect 90638 542200 90694 543000
rect 95054 542200 95110 543000
rect 99470 542200 99526 543000
rect 103886 542200 103942 543000
rect 108302 542200 108358 543000
rect 112718 542200 112774 543000
rect 117134 542200 117190 543000
rect 121550 542200 121606 543000
rect 125966 542200 126022 543000
rect 130382 542200 130438 543000
rect 134798 542200 134854 543000
rect 139214 542200 139270 543000
rect 143630 542200 143686 543000
rect 148046 542200 148102 543000
rect 152462 542200 152518 543000
rect 156878 542200 156934 543000
rect 161294 542200 161350 543000
rect 165710 542200 165766 543000
rect 170126 542200 170182 543000
rect 174542 542200 174598 543000
rect 178958 542200 179014 543000
rect 183374 542200 183430 543000
rect 187790 542200 187846 543000
rect 192206 542200 192262 543000
rect 196622 542200 196678 543000
rect 201038 542200 201094 543000
rect 205454 542200 205510 543000
rect 209870 542200 209926 543000
rect 214286 542200 214342 543000
rect 218702 542200 218758 543000
rect 223118 542200 223174 543000
rect 227534 542200 227590 543000
rect 231950 542200 232006 543000
rect 236366 542200 236422 543000
rect 240782 542200 240838 543000
rect 245198 542200 245254 543000
rect 249614 542200 249670 543000
rect 254030 542200 254086 543000
rect 258446 542200 258502 543000
rect 262862 542200 262918 543000
rect 267278 542200 267334 543000
rect 271694 542200 271750 543000
rect 276110 542200 276166 543000
rect 280526 542200 280582 543000
rect 284942 542200 284998 543000
rect 289358 542200 289414 543000
rect 293774 542200 293830 543000
rect 298190 542200 298246 543000
rect 302606 542200 302662 543000
rect 307022 542200 307078 543000
rect 311438 542200 311494 543000
rect 315854 542200 315910 543000
rect 320270 542200 320326 543000
rect 324686 542200 324742 543000
rect 329102 542200 329158 543000
rect 333518 542200 333574 543000
rect 337934 542200 337990 543000
rect 342350 542200 342406 543000
rect 346766 542200 346822 543000
rect 351182 542200 351238 543000
rect 355598 542200 355654 543000
rect 360014 542200 360070 543000
rect 364430 542200 364486 543000
rect 368846 542200 368902 543000
rect 373262 542200 373318 543000
rect 377678 542200 377734 543000
rect 382094 542200 382150 543000
rect 386510 542200 386566 543000
rect 390926 542200 390982 543000
rect 395342 542200 395398 543000
rect 399758 542200 399814 543000
rect 404174 542200 404230 543000
rect 408590 542200 408646 543000
rect 413006 542200 413062 543000
rect 417422 542200 417478 543000
rect 421838 542200 421894 543000
rect 426254 542200 426310 543000
rect 430670 542200 430726 543000
rect 435086 542200 435142 543000
rect 439502 542200 439558 543000
rect 443918 542200 443974 543000
rect 448334 542200 448390 543000
rect 452750 542200 452806 543000
rect 457166 542200 457222 543000
rect 461582 542200 461638 543000
rect 465998 542200 466054 543000
rect 470414 542200 470470 543000
rect 474830 542200 474886 543000
rect 479246 542200 479302 543000
rect 483662 542200 483718 543000
rect 488078 542200 488134 543000
rect 3974 0 4030 800
rect 9770 0 9826 800
rect 15566 0 15622 800
rect 21362 0 21418 800
rect 27158 0 27214 800
rect 32954 0 33010 800
rect 38750 0 38806 800
rect 44546 0 44602 800
rect 50342 0 50398 800
rect 56138 0 56194 800
rect 61934 0 61990 800
rect 67730 0 67786 800
rect 73526 0 73582 800
rect 79322 0 79378 800
rect 85118 0 85174 800
rect 90914 0 90970 800
rect 96710 0 96766 800
rect 102506 0 102562 800
rect 108302 0 108358 800
rect 114098 0 114154 800
rect 119894 0 119950 800
rect 125690 0 125746 800
rect 131486 0 131542 800
rect 137282 0 137338 800
rect 143078 0 143134 800
rect 148874 0 148930 800
rect 154670 0 154726 800
rect 160466 0 160522 800
rect 166262 0 166318 800
rect 172058 0 172114 800
rect 177854 0 177910 800
rect 183650 0 183706 800
rect 189446 0 189502 800
rect 195242 0 195298 800
rect 201038 0 201094 800
rect 206834 0 206890 800
rect 212630 0 212686 800
rect 218426 0 218482 800
rect 224222 0 224278 800
rect 230018 0 230074 800
rect 235814 0 235870 800
rect 241610 0 241666 800
rect 247406 0 247462 800
rect 253202 0 253258 800
rect 258998 0 259054 800
rect 264794 0 264850 800
rect 270590 0 270646 800
rect 276386 0 276442 800
rect 282182 0 282238 800
rect 287978 0 288034 800
rect 293774 0 293830 800
rect 299570 0 299626 800
rect 305366 0 305422 800
rect 311162 0 311218 800
rect 316958 0 317014 800
rect 322754 0 322810 800
rect 328550 0 328606 800
rect 334346 0 334402 800
rect 340142 0 340198 800
rect 345938 0 345994 800
rect 351734 0 351790 800
rect 357530 0 357586 800
rect 363326 0 363382 800
rect 369122 0 369178 800
rect 374918 0 374974 800
rect 380714 0 380770 800
rect 386510 0 386566 800
rect 392306 0 392362 800
rect 398102 0 398158 800
rect 403898 0 403954 800
rect 409694 0 409750 800
rect 415490 0 415546 800
rect 421286 0 421342 800
rect 427082 0 427138 800
rect 432878 0 432934 800
rect 438674 0 438730 800
rect 444470 0 444526 800
rect 450266 0 450322 800
rect 456062 0 456118 800
rect 461858 0 461914 800
rect 467654 0 467710 800
rect 473450 0 473506 800
rect 479246 0 479302 800
rect 485042 0 485098 800
rect 490838 0 490894 800
<< obsm2 >>
rect 572 542144 6678 542314
rect 6846 542144 11094 542314
rect 11262 542144 15510 542314
rect 15678 542144 19926 542314
rect 20094 542144 24342 542314
rect 24510 542144 28758 542314
rect 28926 542144 33174 542314
rect 33342 542144 37590 542314
rect 37758 542144 42006 542314
rect 42174 542144 46422 542314
rect 46590 542144 50838 542314
rect 51006 542144 55254 542314
rect 55422 542144 59670 542314
rect 59838 542144 64086 542314
rect 64254 542144 68502 542314
rect 68670 542144 72918 542314
rect 73086 542144 77334 542314
rect 77502 542144 81750 542314
rect 81918 542144 86166 542314
rect 86334 542144 90582 542314
rect 90750 542144 94998 542314
rect 95166 542144 99414 542314
rect 99582 542144 103830 542314
rect 103998 542144 108246 542314
rect 108414 542144 112662 542314
rect 112830 542144 117078 542314
rect 117246 542144 121494 542314
rect 121662 542144 125910 542314
rect 126078 542144 130326 542314
rect 130494 542144 134742 542314
rect 134910 542144 139158 542314
rect 139326 542144 143574 542314
rect 143742 542144 147990 542314
rect 148158 542144 152406 542314
rect 152574 542144 156822 542314
rect 156990 542144 161238 542314
rect 161406 542144 165654 542314
rect 165822 542144 170070 542314
rect 170238 542144 174486 542314
rect 174654 542144 178902 542314
rect 179070 542144 183318 542314
rect 183486 542144 187734 542314
rect 187902 542144 192150 542314
rect 192318 542144 196566 542314
rect 196734 542144 200982 542314
rect 201150 542144 205398 542314
rect 205566 542144 209814 542314
rect 209982 542144 214230 542314
rect 214398 542144 218646 542314
rect 218814 542144 223062 542314
rect 223230 542144 227478 542314
rect 227646 542144 231894 542314
rect 232062 542144 236310 542314
rect 236478 542144 240726 542314
rect 240894 542144 245142 542314
rect 245310 542144 249558 542314
rect 249726 542144 253974 542314
rect 254142 542144 258390 542314
rect 258558 542144 262806 542314
rect 262974 542144 267222 542314
rect 267390 542144 271638 542314
rect 271806 542144 276054 542314
rect 276222 542144 280470 542314
rect 280638 542144 284886 542314
rect 285054 542144 289302 542314
rect 289470 542144 293718 542314
rect 293886 542144 298134 542314
rect 298302 542144 302550 542314
rect 302718 542144 306966 542314
rect 307134 542144 311382 542314
rect 311550 542144 315798 542314
rect 315966 542144 320214 542314
rect 320382 542144 324630 542314
rect 324798 542144 329046 542314
rect 329214 542144 333462 542314
rect 333630 542144 337878 542314
rect 338046 542144 342294 542314
rect 342462 542144 346710 542314
rect 346878 542144 351126 542314
rect 351294 542144 355542 542314
rect 355710 542144 359958 542314
rect 360126 542144 364374 542314
rect 364542 542144 368790 542314
rect 368958 542144 373206 542314
rect 373374 542144 377622 542314
rect 377790 542144 382038 542314
rect 382206 542144 386454 542314
rect 386622 542144 390870 542314
rect 391038 542144 395286 542314
rect 395454 542144 399702 542314
rect 399870 542144 404118 542314
rect 404286 542144 408534 542314
rect 408702 542144 412950 542314
rect 413118 542144 417366 542314
rect 417534 542144 421782 542314
rect 421950 542144 426198 542314
rect 426366 542144 430614 542314
rect 430782 542144 435030 542314
rect 435198 542144 439446 542314
rect 439614 542144 443862 542314
rect 444030 542144 448278 542314
rect 448446 542144 452694 542314
rect 452862 542144 457110 542314
rect 457278 542144 461526 542314
rect 461694 542144 465942 542314
rect 466110 542144 470358 542314
rect 470526 542144 474774 542314
rect 474942 542144 479190 542314
rect 479358 542144 483606 542314
rect 483774 542144 488022 542314
rect 488190 542144 494572 542314
rect 572 856 494572 542144
rect 572 734 3918 856
rect 4086 734 9714 856
rect 9882 734 15510 856
rect 15678 734 21306 856
rect 21474 734 27102 856
rect 27270 734 32898 856
rect 33066 734 38694 856
rect 38862 734 44490 856
rect 44658 734 50286 856
rect 50454 734 56082 856
rect 56250 734 61878 856
rect 62046 734 67674 856
rect 67842 734 73470 856
rect 73638 734 79266 856
rect 79434 734 85062 856
rect 85230 734 90858 856
rect 91026 734 96654 856
rect 96822 734 102450 856
rect 102618 734 108246 856
rect 108414 734 114042 856
rect 114210 734 119838 856
rect 120006 734 125634 856
rect 125802 734 131430 856
rect 131598 734 137226 856
rect 137394 734 143022 856
rect 143190 734 148818 856
rect 148986 734 154614 856
rect 154782 734 160410 856
rect 160578 734 166206 856
rect 166374 734 172002 856
rect 172170 734 177798 856
rect 177966 734 183594 856
rect 183762 734 189390 856
rect 189558 734 195186 856
rect 195354 734 200982 856
rect 201150 734 206778 856
rect 206946 734 212574 856
rect 212742 734 218370 856
rect 218538 734 224166 856
rect 224334 734 229962 856
rect 230130 734 235758 856
rect 235926 734 241554 856
rect 241722 734 247350 856
rect 247518 734 253146 856
rect 253314 734 258942 856
rect 259110 734 264738 856
rect 264906 734 270534 856
rect 270702 734 276330 856
rect 276498 734 282126 856
rect 282294 734 287922 856
rect 288090 734 293718 856
rect 293886 734 299514 856
rect 299682 734 305310 856
rect 305478 734 311106 856
rect 311274 734 316902 856
rect 317070 734 322698 856
rect 322866 734 328494 856
rect 328662 734 334290 856
rect 334458 734 340086 856
rect 340254 734 345882 856
rect 346050 734 351678 856
rect 351846 734 357474 856
rect 357642 734 363270 856
rect 363438 734 369066 856
rect 369234 734 374862 856
rect 375030 734 380658 856
rect 380826 734 386454 856
rect 386622 734 392250 856
rect 392418 734 398046 856
rect 398214 734 403842 856
rect 404010 734 409638 856
rect 409806 734 415434 856
rect 415602 734 421230 856
rect 421398 734 427026 856
rect 427194 734 432822 856
rect 432990 734 438618 856
rect 438786 734 444414 856
rect 444582 734 450210 856
rect 450378 734 456006 856
rect 456174 734 461802 856
rect 461970 734 467598 856
rect 467766 734 473394 856
rect 473562 734 479190 856
rect 479358 734 484986 856
rect 485154 734 490782 856
rect 490950 734 494572 856
<< metal3 >>
rect 0 537888 800 538008
rect 494200 533944 495000 534064
rect 0 532448 800 532568
rect 494200 528640 495000 528760
rect 0 527008 800 527128
rect 494200 523336 495000 523456
rect 0 521568 800 521688
rect 494200 518032 495000 518152
rect 0 516128 800 516248
rect 494200 512728 495000 512848
rect 0 510688 800 510808
rect 494200 507424 495000 507544
rect 0 505248 800 505368
rect 494200 502120 495000 502240
rect 0 499808 800 499928
rect 494200 496816 495000 496936
rect 0 494368 800 494488
rect 494200 491512 495000 491632
rect 0 488928 800 489048
rect 494200 486208 495000 486328
rect 0 483488 800 483608
rect 494200 480904 495000 481024
rect 0 478048 800 478168
rect 494200 475600 495000 475720
rect 0 472608 800 472728
rect 494200 470296 495000 470416
rect 0 467168 800 467288
rect 494200 464992 495000 465112
rect 0 461728 800 461848
rect 494200 459688 495000 459808
rect 0 456288 800 456408
rect 494200 454384 495000 454504
rect 0 450848 800 450968
rect 494200 449080 495000 449200
rect 0 445408 800 445528
rect 494200 443776 495000 443896
rect 0 439968 800 440088
rect 494200 438472 495000 438592
rect 0 434528 800 434648
rect 494200 433168 495000 433288
rect 0 429088 800 429208
rect 494200 427864 495000 427984
rect 0 423648 800 423768
rect 494200 422560 495000 422680
rect 0 418208 800 418328
rect 494200 417256 495000 417376
rect 0 412768 800 412888
rect 494200 411952 495000 412072
rect 0 407328 800 407448
rect 494200 406648 495000 406768
rect 0 401888 800 402008
rect 494200 401344 495000 401464
rect 0 396448 800 396568
rect 494200 396040 495000 396160
rect 0 391008 800 391128
rect 494200 390736 495000 390856
rect 0 385568 800 385688
rect 494200 385432 495000 385552
rect 0 380128 800 380248
rect 494200 380128 495000 380248
rect 0 374688 800 374808
rect 494200 374824 495000 374944
rect 494200 369520 495000 369640
rect 0 369248 800 369368
rect 494200 364216 495000 364336
rect 0 363808 800 363928
rect 494200 358912 495000 359032
rect 0 358368 800 358488
rect 494200 353608 495000 353728
rect 0 352928 800 353048
rect 494200 348304 495000 348424
rect 0 347488 800 347608
rect 494200 343000 495000 343120
rect 0 342048 800 342168
rect 494200 337696 495000 337816
rect 0 336608 800 336728
rect 494200 332392 495000 332512
rect 0 331168 800 331288
rect 494200 327088 495000 327208
rect 0 325728 800 325848
rect 494200 321784 495000 321904
rect 0 320288 800 320408
rect 494200 316480 495000 316600
rect 0 314848 800 314968
rect 494200 311176 495000 311296
rect 0 309408 800 309528
rect 494200 305872 495000 305992
rect 0 303968 800 304088
rect 494200 300568 495000 300688
rect 0 298528 800 298648
rect 494200 295264 495000 295384
rect 0 293088 800 293208
rect 494200 289960 495000 290080
rect 0 287648 800 287768
rect 494200 284656 495000 284776
rect 0 282208 800 282328
rect 494200 279352 495000 279472
rect 0 276768 800 276888
rect 494200 274048 495000 274168
rect 0 271328 800 271448
rect 494200 268744 495000 268864
rect 0 265888 800 266008
rect 494200 263440 495000 263560
rect 0 260448 800 260568
rect 494200 258136 495000 258256
rect 0 255008 800 255128
rect 494200 252832 495000 252952
rect 0 249568 800 249688
rect 494200 247528 495000 247648
rect 0 244128 800 244248
rect 494200 242224 495000 242344
rect 0 238688 800 238808
rect 494200 236920 495000 237040
rect 0 233248 800 233368
rect 494200 231616 495000 231736
rect 0 227808 800 227928
rect 494200 226312 495000 226432
rect 0 222368 800 222488
rect 494200 221008 495000 221128
rect 0 216928 800 217048
rect 494200 215704 495000 215824
rect 0 211488 800 211608
rect 494200 210400 495000 210520
rect 0 206048 800 206168
rect 494200 205096 495000 205216
rect 0 200608 800 200728
rect 494200 199792 495000 199912
rect 0 195168 800 195288
rect 494200 194488 495000 194608
rect 0 189728 800 189848
rect 494200 189184 495000 189304
rect 0 184288 800 184408
rect 494200 183880 495000 184000
rect 0 178848 800 178968
rect 494200 178576 495000 178696
rect 0 173408 800 173528
rect 494200 173272 495000 173392
rect 0 167968 800 168088
rect 494200 167968 495000 168088
rect 0 162528 800 162648
rect 494200 162664 495000 162784
rect 494200 157360 495000 157480
rect 0 157088 800 157208
rect 494200 152056 495000 152176
rect 0 151648 800 151768
rect 494200 146752 495000 146872
rect 0 146208 800 146328
rect 494200 141448 495000 141568
rect 0 140768 800 140888
rect 494200 136144 495000 136264
rect 0 135328 800 135448
rect 494200 130840 495000 130960
rect 0 129888 800 130008
rect 494200 125536 495000 125656
rect 0 124448 800 124568
rect 494200 120232 495000 120352
rect 0 119008 800 119128
rect 494200 114928 495000 115048
rect 0 113568 800 113688
rect 494200 109624 495000 109744
rect 0 108128 800 108248
rect 494200 104320 495000 104440
rect 0 102688 800 102808
rect 494200 99016 495000 99136
rect 0 97248 800 97368
rect 494200 93712 495000 93832
rect 0 91808 800 91928
rect 494200 88408 495000 88528
rect 0 86368 800 86488
rect 494200 83104 495000 83224
rect 0 80928 800 81048
rect 494200 77800 495000 77920
rect 0 75488 800 75608
rect 494200 72496 495000 72616
rect 0 70048 800 70168
rect 494200 67192 495000 67312
rect 0 64608 800 64728
rect 494200 61888 495000 62008
rect 0 59168 800 59288
rect 494200 56584 495000 56704
rect 0 53728 800 53848
rect 494200 51280 495000 51400
rect 0 48288 800 48408
rect 494200 45976 495000 46096
rect 0 42848 800 42968
rect 494200 40672 495000 40792
rect 0 37408 800 37528
rect 494200 35368 495000 35488
rect 0 31968 800 32088
rect 494200 30064 495000 30184
rect 0 26528 800 26648
rect 494200 24760 495000 24880
rect 0 21088 800 21208
rect 494200 19456 495000 19576
rect 0 15648 800 15768
rect 494200 14152 495000 14272
rect 0 10208 800 10328
rect 494200 8848 495000 8968
rect 0 4768 800 4888
<< obsm3 >>
rect 657 538088 494200 540769
rect 880 537808 494200 538088
rect 657 534144 494200 537808
rect 657 533864 494120 534144
rect 657 532648 494200 533864
rect 880 532368 494200 532648
rect 657 528840 494200 532368
rect 657 528560 494120 528840
rect 657 527208 494200 528560
rect 880 526928 494200 527208
rect 657 523536 494200 526928
rect 657 523256 494120 523536
rect 657 521768 494200 523256
rect 880 521488 494200 521768
rect 657 518232 494200 521488
rect 657 517952 494120 518232
rect 657 516328 494200 517952
rect 880 516048 494200 516328
rect 657 512928 494200 516048
rect 657 512648 494120 512928
rect 657 510888 494200 512648
rect 880 510608 494200 510888
rect 657 507624 494200 510608
rect 657 507344 494120 507624
rect 657 505448 494200 507344
rect 880 505168 494200 505448
rect 657 502320 494200 505168
rect 657 502040 494120 502320
rect 657 500008 494200 502040
rect 880 499728 494200 500008
rect 657 497016 494200 499728
rect 657 496736 494120 497016
rect 657 494568 494200 496736
rect 880 494288 494200 494568
rect 657 491712 494200 494288
rect 657 491432 494120 491712
rect 657 489128 494200 491432
rect 880 488848 494200 489128
rect 657 486408 494200 488848
rect 657 486128 494120 486408
rect 657 483688 494200 486128
rect 880 483408 494200 483688
rect 657 481104 494200 483408
rect 657 480824 494120 481104
rect 657 478248 494200 480824
rect 880 477968 494200 478248
rect 657 475800 494200 477968
rect 657 475520 494120 475800
rect 657 472808 494200 475520
rect 880 472528 494200 472808
rect 657 470496 494200 472528
rect 657 470216 494120 470496
rect 657 467368 494200 470216
rect 880 467088 494200 467368
rect 657 465192 494200 467088
rect 657 464912 494120 465192
rect 657 461928 494200 464912
rect 880 461648 494200 461928
rect 657 459888 494200 461648
rect 657 459608 494120 459888
rect 657 456488 494200 459608
rect 880 456208 494200 456488
rect 657 454584 494200 456208
rect 657 454304 494120 454584
rect 657 451048 494200 454304
rect 880 450768 494200 451048
rect 657 449280 494200 450768
rect 657 449000 494120 449280
rect 657 445608 494200 449000
rect 880 445328 494200 445608
rect 657 443976 494200 445328
rect 657 443696 494120 443976
rect 657 440168 494200 443696
rect 880 439888 494200 440168
rect 657 438672 494200 439888
rect 657 438392 494120 438672
rect 657 434728 494200 438392
rect 880 434448 494200 434728
rect 657 433368 494200 434448
rect 657 433088 494120 433368
rect 657 429288 494200 433088
rect 880 429008 494200 429288
rect 657 428064 494200 429008
rect 657 427784 494120 428064
rect 657 423848 494200 427784
rect 880 423568 494200 423848
rect 657 422760 494200 423568
rect 657 422480 494120 422760
rect 657 418408 494200 422480
rect 880 418128 494200 418408
rect 657 417456 494200 418128
rect 657 417176 494120 417456
rect 657 412968 494200 417176
rect 880 412688 494200 412968
rect 657 412152 494200 412688
rect 657 411872 494120 412152
rect 657 407528 494200 411872
rect 880 407248 494200 407528
rect 657 406848 494200 407248
rect 657 406568 494120 406848
rect 657 402088 494200 406568
rect 880 401808 494200 402088
rect 657 401544 494200 401808
rect 657 401264 494120 401544
rect 657 396648 494200 401264
rect 880 396368 494200 396648
rect 657 396240 494200 396368
rect 657 395960 494120 396240
rect 657 391208 494200 395960
rect 880 390936 494200 391208
rect 880 390928 494120 390936
rect 657 390656 494120 390928
rect 657 385768 494200 390656
rect 880 385632 494200 385768
rect 880 385488 494120 385632
rect 657 385352 494120 385488
rect 657 380328 494200 385352
rect 880 380048 494120 380328
rect 657 375024 494200 380048
rect 657 374888 494120 375024
rect 880 374744 494120 374888
rect 880 374608 494200 374744
rect 657 369720 494200 374608
rect 657 369448 494120 369720
rect 880 369440 494120 369448
rect 880 369168 494200 369440
rect 657 364416 494200 369168
rect 657 364136 494120 364416
rect 657 364008 494200 364136
rect 880 363728 494200 364008
rect 657 359112 494200 363728
rect 657 358832 494120 359112
rect 657 358568 494200 358832
rect 880 358288 494200 358568
rect 657 353808 494200 358288
rect 657 353528 494120 353808
rect 657 353128 494200 353528
rect 880 352848 494200 353128
rect 657 348504 494200 352848
rect 657 348224 494120 348504
rect 657 347688 494200 348224
rect 880 347408 494200 347688
rect 657 343200 494200 347408
rect 657 342920 494120 343200
rect 657 342248 494200 342920
rect 880 341968 494200 342248
rect 657 337896 494200 341968
rect 657 337616 494120 337896
rect 657 336808 494200 337616
rect 880 336528 494200 336808
rect 657 332592 494200 336528
rect 657 332312 494120 332592
rect 657 331368 494200 332312
rect 880 331088 494200 331368
rect 657 327288 494200 331088
rect 657 327008 494120 327288
rect 657 325928 494200 327008
rect 880 325648 494200 325928
rect 657 321984 494200 325648
rect 657 321704 494120 321984
rect 657 320488 494200 321704
rect 880 320208 494200 320488
rect 657 316680 494200 320208
rect 657 316400 494120 316680
rect 657 315048 494200 316400
rect 880 314768 494200 315048
rect 657 311376 494200 314768
rect 657 311096 494120 311376
rect 657 309608 494200 311096
rect 880 309328 494200 309608
rect 657 306072 494200 309328
rect 657 305792 494120 306072
rect 657 304168 494200 305792
rect 880 303888 494200 304168
rect 657 300768 494200 303888
rect 657 300488 494120 300768
rect 657 298728 494200 300488
rect 880 298448 494200 298728
rect 657 295464 494200 298448
rect 657 295184 494120 295464
rect 657 293288 494200 295184
rect 880 293008 494200 293288
rect 657 290160 494200 293008
rect 657 289880 494120 290160
rect 657 287848 494200 289880
rect 880 287568 494200 287848
rect 657 284856 494200 287568
rect 657 284576 494120 284856
rect 657 282408 494200 284576
rect 880 282128 494200 282408
rect 657 279552 494200 282128
rect 657 279272 494120 279552
rect 657 276968 494200 279272
rect 880 276688 494200 276968
rect 657 274248 494200 276688
rect 657 273968 494120 274248
rect 657 271528 494200 273968
rect 880 271248 494200 271528
rect 657 268944 494200 271248
rect 657 268664 494120 268944
rect 657 266088 494200 268664
rect 880 265808 494200 266088
rect 657 263640 494200 265808
rect 657 263360 494120 263640
rect 657 260648 494200 263360
rect 880 260368 494200 260648
rect 657 258336 494200 260368
rect 657 258056 494120 258336
rect 657 255208 494200 258056
rect 880 254928 494200 255208
rect 657 253032 494200 254928
rect 657 252752 494120 253032
rect 657 249768 494200 252752
rect 880 249488 494200 249768
rect 657 247728 494200 249488
rect 657 247448 494120 247728
rect 657 244328 494200 247448
rect 880 244048 494200 244328
rect 657 242424 494200 244048
rect 657 242144 494120 242424
rect 657 238888 494200 242144
rect 880 238608 494200 238888
rect 657 237120 494200 238608
rect 657 236840 494120 237120
rect 657 233448 494200 236840
rect 880 233168 494200 233448
rect 657 231816 494200 233168
rect 657 231536 494120 231816
rect 657 228008 494200 231536
rect 880 227728 494200 228008
rect 657 226512 494200 227728
rect 657 226232 494120 226512
rect 657 222568 494200 226232
rect 880 222288 494200 222568
rect 657 221208 494200 222288
rect 657 220928 494120 221208
rect 657 217128 494200 220928
rect 880 216848 494200 217128
rect 657 215904 494200 216848
rect 657 215624 494120 215904
rect 657 211688 494200 215624
rect 880 211408 494200 211688
rect 657 210600 494200 211408
rect 657 210320 494120 210600
rect 657 206248 494200 210320
rect 880 205968 494200 206248
rect 657 205296 494200 205968
rect 657 205016 494120 205296
rect 657 200808 494200 205016
rect 880 200528 494200 200808
rect 657 199992 494200 200528
rect 657 199712 494120 199992
rect 657 195368 494200 199712
rect 880 195088 494200 195368
rect 657 194688 494200 195088
rect 657 194408 494120 194688
rect 657 189928 494200 194408
rect 880 189648 494200 189928
rect 657 189384 494200 189648
rect 657 189104 494120 189384
rect 657 184488 494200 189104
rect 880 184208 494200 184488
rect 657 184080 494200 184208
rect 657 183800 494120 184080
rect 657 179048 494200 183800
rect 880 178776 494200 179048
rect 880 178768 494120 178776
rect 657 178496 494120 178768
rect 657 173608 494200 178496
rect 880 173472 494200 173608
rect 880 173328 494120 173472
rect 657 173192 494120 173328
rect 657 168168 494200 173192
rect 880 167888 494120 168168
rect 657 162864 494200 167888
rect 657 162728 494120 162864
rect 880 162584 494120 162728
rect 880 162448 494200 162584
rect 657 157560 494200 162448
rect 657 157288 494120 157560
rect 880 157280 494120 157288
rect 880 157008 494200 157280
rect 657 152256 494200 157008
rect 657 151976 494120 152256
rect 657 151848 494200 151976
rect 880 151568 494200 151848
rect 657 146952 494200 151568
rect 657 146672 494120 146952
rect 657 146408 494200 146672
rect 880 146128 494200 146408
rect 657 141648 494200 146128
rect 657 141368 494120 141648
rect 657 140968 494200 141368
rect 880 140688 494200 140968
rect 657 136344 494200 140688
rect 657 136064 494120 136344
rect 657 135528 494200 136064
rect 880 135248 494200 135528
rect 657 131040 494200 135248
rect 657 130760 494120 131040
rect 657 130088 494200 130760
rect 880 129808 494200 130088
rect 657 125736 494200 129808
rect 657 125456 494120 125736
rect 657 124648 494200 125456
rect 880 124368 494200 124648
rect 657 120432 494200 124368
rect 657 120152 494120 120432
rect 657 119208 494200 120152
rect 880 118928 494200 119208
rect 657 115128 494200 118928
rect 657 114848 494120 115128
rect 657 113768 494200 114848
rect 880 113488 494200 113768
rect 657 109824 494200 113488
rect 657 109544 494120 109824
rect 657 108328 494200 109544
rect 880 108048 494200 108328
rect 657 104520 494200 108048
rect 657 104240 494120 104520
rect 657 102888 494200 104240
rect 880 102608 494200 102888
rect 657 99216 494200 102608
rect 657 98936 494120 99216
rect 657 97448 494200 98936
rect 880 97168 494200 97448
rect 657 93912 494200 97168
rect 657 93632 494120 93912
rect 657 92008 494200 93632
rect 880 91728 494200 92008
rect 657 88608 494200 91728
rect 657 88328 494120 88608
rect 657 86568 494200 88328
rect 880 86288 494200 86568
rect 657 83304 494200 86288
rect 657 83024 494120 83304
rect 657 81128 494200 83024
rect 880 80848 494200 81128
rect 657 78000 494200 80848
rect 657 77720 494120 78000
rect 657 75688 494200 77720
rect 880 75408 494200 75688
rect 657 72696 494200 75408
rect 657 72416 494120 72696
rect 657 70248 494200 72416
rect 880 69968 494200 70248
rect 657 67392 494200 69968
rect 657 67112 494120 67392
rect 657 64808 494200 67112
rect 880 64528 494200 64808
rect 657 62088 494200 64528
rect 657 61808 494120 62088
rect 657 59368 494200 61808
rect 880 59088 494200 59368
rect 657 56784 494200 59088
rect 657 56504 494120 56784
rect 657 53928 494200 56504
rect 880 53648 494200 53928
rect 657 51480 494200 53648
rect 657 51200 494120 51480
rect 657 48488 494200 51200
rect 880 48208 494200 48488
rect 657 46176 494200 48208
rect 657 45896 494120 46176
rect 657 43048 494200 45896
rect 880 42768 494200 43048
rect 657 40872 494200 42768
rect 657 40592 494120 40872
rect 657 37608 494200 40592
rect 880 37328 494200 37608
rect 657 35568 494200 37328
rect 657 35288 494120 35568
rect 657 32168 494200 35288
rect 880 31888 494200 32168
rect 657 30264 494200 31888
rect 657 29984 494120 30264
rect 657 26728 494200 29984
rect 880 26448 494200 26728
rect 657 24960 494200 26448
rect 657 24680 494120 24960
rect 657 21288 494200 24680
rect 880 21008 494200 21288
rect 657 19656 494200 21008
rect 657 19376 494120 19656
rect 657 15848 494200 19376
rect 880 15568 494200 15848
rect 657 14352 494200 15568
rect 657 14072 494120 14352
rect 657 10408 494200 14072
rect 880 10128 494200 10408
rect 657 9048 494200 10128
rect 657 8768 494120 9048
rect 657 4968 494200 8768
rect 880 4688 494200 4968
rect 657 2143 494200 4688
<< metal4 >>
rect -2552 -744 -1592 543656
rect -1192 616 -232 542296
rect 1024 -744 1664 543656
rect 1984 -744 2624 543656
rect 12424 471657 13064 543656
rect 13384 536508 14024 543656
rect 23824 536508 24464 543656
rect 24784 520921 25424 543656
rect 13384 473508 14024 480068
rect 23824 473508 24464 480068
rect 24784 471657 25424 481375
rect 12424 408657 13064 418919
rect 13384 410508 14024 417068
rect 23824 410508 24464 417068
rect 24784 408657 25424 418919
rect 12424 345657 13064 355919
rect 13384 347508 14024 354068
rect 23824 347508 24464 354068
rect 24784 345657 25424 355919
rect 12424 282657 13064 292919
rect 13384 284508 14024 291068
rect 23824 284508 24464 291068
rect 24784 282657 25424 292919
rect 12424 219657 13064 229919
rect 13384 221508 14024 228068
rect 23824 221508 24464 228068
rect 24784 219657 25424 229919
rect 12424 156657 13064 166919
rect 13384 158508 14024 165068
rect 23824 158508 24464 165068
rect 24784 156657 25424 166919
rect 12424 93657 13064 103919
rect 13384 95508 14024 102068
rect 23824 95508 24464 102068
rect 24784 93657 25424 103919
rect 12424 34409 13064 40919
rect 13384 34409 14024 39068
rect 23824 34409 24464 39068
rect 24784 34409 25424 40919
rect 12424 -744 13064 12271
rect 13384 -744 14024 6068
rect 23824 -744 24464 6068
rect 24784 -744 25424 12271
rect 35224 -744 35864 543656
rect 36184 -744 36824 543656
rect 46624 536508 47264 543656
rect 47584 535609 48224 543656
rect 58024 535609 58664 543656
rect 58984 535609 59624 543656
rect 69424 535609 70064 543656
rect 70384 535609 71024 543656
rect 80824 535609 81464 543656
rect 81784 536508 82424 543656
rect 46624 473508 47264 480068
rect 47584 473153 48224 480423
rect 58024 473153 58664 480423
rect 58984 473153 59624 480423
rect 69424 473153 70064 480423
rect 70384 473153 71024 480423
rect 80824 473153 81464 480423
rect 81784 473508 82424 480068
rect 46624 410508 47264 417068
rect 47584 410153 48224 417423
rect 58024 410153 58664 417423
rect 58984 410153 59624 417423
rect 69424 410153 70064 417423
rect 70384 410153 71024 417423
rect 80824 410153 81464 417423
rect 81784 410508 82424 417068
rect 46624 347508 47264 354068
rect 47584 347153 48224 354423
rect 58024 347153 58664 354423
rect 58984 347153 59624 354423
rect 69424 347153 70064 354423
rect 70384 347153 71024 354423
rect 80824 347153 81464 354423
rect 81784 347508 82424 354068
rect 46624 284508 47264 291068
rect 47584 284153 48224 291423
rect 58024 284153 58664 291423
rect 58984 284153 59624 291423
rect 69424 284153 70064 291423
rect 70384 284153 71024 291423
rect 80824 284153 81464 291423
rect 81784 284508 82424 291068
rect 46624 221508 47264 228068
rect 47584 221153 48224 228423
rect 58024 221153 58664 228423
rect 58984 221153 59624 228423
rect 69424 221153 70064 228423
rect 70384 221153 71024 228423
rect 80824 221153 81464 228423
rect 81784 221508 82424 228068
rect 46624 158508 47264 165068
rect 47584 158153 48224 165423
rect 58024 158153 58664 165423
rect 58984 158153 59624 165423
rect 69424 158153 70064 165423
rect 70384 158153 71024 165423
rect 80824 158153 81464 165423
rect 81784 158508 82424 165068
rect 46624 95508 47264 102068
rect 47584 95153 48224 102423
rect 58024 95153 58664 102423
rect 58984 95153 59624 102423
rect 69424 95153 70064 102423
rect 70384 95153 71024 102423
rect 80824 95153 81464 102423
rect 81784 95508 82424 102068
rect 46624 32588 47264 39068
rect 46624 -744 47264 6068
rect 47584 -744 48224 39423
rect 58024 32233 58664 39423
rect 58984 32233 59624 39423
rect 69424 32233 70064 39423
rect 70384 32233 71024 39423
rect 58024 -744 58664 10639
rect 58984 -744 59624 10639
rect 69424 -744 70064 10639
rect 70384 -744 71024 10639
rect 80824 -744 81464 39423
rect 81784 32588 82424 39068
rect 81784 -744 82424 6068
rect 92224 -744 92864 543656
rect 93184 -744 93824 543656
rect 103624 536508 104264 543656
rect 104584 535609 105224 543656
rect 115024 535609 115664 543656
rect 115984 535609 116624 543656
rect 126424 535609 127064 543656
rect 127384 535609 128024 543656
rect 137824 535609 138464 543656
rect 138784 536508 139424 543656
rect 103624 473508 104264 480068
rect 104584 473153 105224 480423
rect 115024 473153 115664 480423
rect 115984 473153 116624 480423
rect 126424 473153 127064 480423
rect 127384 473153 128024 480423
rect 137824 473153 138464 480423
rect 138784 473508 139424 480068
rect 103624 410508 104264 417068
rect 104584 410153 105224 417423
rect 115024 410153 115664 417423
rect 115984 410153 116624 417423
rect 126424 410153 127064 417423
rect 127384 410153 128024 417423
rect 137824 410153 138464 417423
rect 138784 410508 139424 417068
rect 103624 347508 104264 354068
rect 104584 347153 105224 354423
rect 115024 347153 115664 354423
rect 115984 347153 116624 354423
rect 126424 347153 127064 354423
rect 127384 347153 128024 354423
rect 137824 347153 138464 354423
rect 138784 347508 139424 354068
rect 103624 284508 104264 291068
rect 104584 284153 105224 291423
rect 115024 284153 115664 291423
rect 115984 284153 116624 291423
rect 126424 284153 127064 291423
rect 127384 284153 128024 291423
rect 137824 284153 138464 291423
rect 138784 284508 139424 291068
rect 103624 221508 104264 228068
rect 104584 221153 105224 228423
rect 115024 221153 115664 228423
rect 115984 221153 116624 228423
rect 126424 221153 127064 228423
rect 127384 221153 128024 228423
rect 137824 221153 138464 228423
rect 138784 221508 139424 228068
rect 103624 158508 104264 165068
rect 104584 158153 105224 165423
rect 115024 158153 115664 165423
rect 115984 158153 116624 165423
rect 126424 158153 127064 165423
rect 127384 158153 128024 165423
rect 137824 158153 138464 165423
rect 138784 158508 139424 165068
rect 103624 95508 104264 102068
rect 104584 95153 105224 102423
rect 115024 95153 115664 102423
rect 115984 95153 116624 102423
rect 126424 95153 127064 102423
rect 127384 95153 128024 102423
rect 137824 95153 138464 102423
rect 138784 95508 139424 102068
rect 103624 32588 104264 39068
rect 103624 -744 104264 6068
rect 104584 -744 105224 39423
rect 115024 32233 115664 39423
rect 115984 32233 116624 39423
rect 126424 32233 127064 39423
rect 127384 32233 128024 39423
rect 115024 -744 115664 10639
rect 115984 -744 116624 10639
rect 126424 -744 127064 10639
rect 127384 -744 128024 10639
rect 137824 -744 138464 39423
rect 138784 32588 139424 39068
rect 138784 -744 139424 6068
rect 149224 -744 149864 543656
rect 150184 -744 150824 543656
rect 160624 536508 161264 543656
rect 161584 535609 162224 543656
rect 172024 535609 172664 543656
rect 172984 535609 173624 543656
rect 183424 535609 184064 543656
rect 184384 535609 185024 543656
rect 194824 535609 195464 543656
rect 195784 536508 196424 543656
rect 160624 473508 161264 480068
rect 161584 473153 162224 480423
rect 172024 473153 172664 480423
rect 172984 473153 173624 480423
rect 183424 473153 184064 480423
rect 184384 473153 185024 480423
rect 194824 473153 195464 480423
rect 195784 473508 196424 480068
rect 160624 410508 161264 417068
rect 161584 410153 162224 417423
rect 172024 410153 172664 417423
rect 172984 410153 173624 417423
rect 183424 410153 184064 417423
rect 184384 410153 185024 417423
rect 194824 410153 195464 417423
rect 195784 410508 196424 417068
rect 160624 347508 161264 354068
rect 161584 347153 162224 354423
rect 172024 347153 172664 354423
rect 172984 347153 173624 354423
rect 183424 347153 184064 354423
rect 184384 347153 185024 354423
rect 194824 347153 195464 354423
rect 195784 347508 196424 354068
rect 160624 284508 161264 291068
rect 161584 284153 162224 291423
rect 172024 284153 172664 291423
rect 172984 284153 173624 291423
rect 183424 284153 184064 291423
rect 184384 284153 185024 291423
rect 194824 284153 195464 291423
rect 195784 284508 196424 291068
rect 160624 221508 161264 228068
rect 161584 221153 162224 228423
rect 172024 221153 172664 228423
rect 172984 221153 173624 228423
rect 183424 221153 184064 228423
rect 184384 221153 185024 228423
rect 194824 221153 195464 228423
rect 195784 221508 196424 228068
rect 160624 158508 161264 165068
rect 161584 158153 162224 165423
rect 172024 158153 172664 165423
rect 172984 158153 173624 165423
rect 183424 158153 184064 165423
rect 184384 158153 185024 165423
rect 194824 158153 195464 165423
rect 195784 158508 196424 165068
rect 160624 95508 161264 102068
rect 161584 95153 162224 102423
rect 172024 95153 172664 102423
rect 172984 95153 173624 102423
rect 183424 95153 184064 102423
rect 184384 95153 185024 102423
rect 194824 95153 195464 102423
rect 195784 95508 196424 102068
rect 160624 32588 161264 39068
rect 160624 -744 161264 6068
rect 161584 -744 162224 39423
rect 172024 32233 172664 39423
rect 172984 32233 173624 39423
rect 183424 32233 184064 39423
rect 184384 32233 185024 39423
rect 172024 -744 172664 10639
rect 172984 -744 173624 10639
rect 183424 -744 184064 10639
rect 184384 -744 185024 10639
rect 194824 -744 195464 39423
rect 195784 32588 196424 39068
rect 195784 -744 196424 6068
rect 206224 -744 206864 543656
rect 207184 -744 207824 543656
rect 217624 536508 218264 543656
rect 218584 535609 219224 543656
rect 229024 535609 229664 543656
rect 229984 535609 230624 543656
rect 240424 535609 241064 543656
rect 241384 535609 242024 543656
rect 251824 535609 252464 543656
rect 252784 536508 253424 543656
rect 217624 473508 218264 480068
rect 218584 473153 219224 480423
rect 229024 473153 229664 480423
rect 229984 473153 230624 480423
rect 240424 473153 241064 480423
rect 241384 473153 242024 480423
rect 251824 473153 252464 480423
rect 252784 473508 253424 480068
rect 217624 410508 218264 417068
rect 218584 410153 219224 417423
rect 229024 410153 229664 417423
rect 229984 410153 230624 417423
rect 240424 410153 241064 417423
rect 241384 410153 242024 417423
rect 251824 410153 252464 417423
rect 252784 410508 253424 417068
rect 217624 347508 218264 354068
rect 218584 347153 219224 354423
rect 229024 347153 229664 354423
rect 229984 347153 230624 354423
rect 240424 347153 241064 354423
rect 241384 347153 242024 354423
rect 251824 347153 252464 354423
rect 252784 347508 253424 354068
rect 217624 284508 218264 291068
rect 218584 284153 219224 291423
rect 229024 284153 229664 291423
rect 229984 284153 230624 291423
rect 240424 284153 241064 291423
rect 241384 284153 242024 291423
rect 251824 284153 252464 291423
rect 252784 284508 253424 291068
rect 217624 221508 218264 228068
rect 218584 221153 219224 228423
rect 229024 221153 229664 228423
rect 229984 221153 230624 228423
rect 240424 221153 241064 228423
rect 241384 221153 242024 228423
rect 251824 221153 252464 228423
rect 252784 221508 253424 228068
rect 217624 158508 218264 165068
rect 218584 158153 219224 165423
rect 229024 158153 229664 165423
rect 229984 158153 230624 165423
rect 240424 158153 241064 165423
rect 241384 158153 242024 165423
rect 251824 158153 252464 165423
rect 252784 158508 253424 165068
rect 217624 95508 218264 102068
rect 218584 95153 219224 102423
rect 229024 95153 229664 102423
rect 229984 95153 230624 102423
rect 240424 95153 241064 102423
rect 241384 95153 242024 102423
rect 251824 95153 252464 102423
rect 252784 95508 253424 102068
rect 217624 32588 218264 39068
rect 217624 -744 218264 6068
rect 218584 -744 219224 39423
rect 229024 32233 229664 39423
rect 229984 32233 230624 39423
rect 240424 32233 241064 39423
rect 241384 32233 242024 39423
rect 229024 -744 229664 10639
rect 229984 -744 230624 10639
rect 240424 -744 241064 10639
rect 241384 -744 242024 10639
rect 251824 -744 252464 39423
rect 252784 32588 253424 39068
rect 252784 -744 253424 6068
rect 263224 -744 263864 543656
rect 264184 -744 264824 543656
rect 274624 536508 275264 543656
rect 275584 535609 276224 543656
rect 286024 535609 286664 543656
rect 286984 535609 287624 543656
rect 297424 535609 298064 543656
rect 298384 535609 299024 543656
rect 308824 535609 309464 543656
rect 309784 536508 310424 543656
rect 274624 473508 275264 480068
rect 275584 473153 276224 480423
rect 286024 473153 286664 480423
rect 286984 473153 287624 480423
rect 297424 473153 298064 480423
rect 298384 473153 299024 480423
rect 308824 473153 309464 480423
rect 309784 473508 310424 480068
rect 274624 410508 275264 417068
rect 275584 410153 276224 417423
rect 286024 410153 286664 417423
rect 286984 410153 287624 417423
rect 297424 410153 298064 417423
rect 298384 410153 299024 417423
rect 308824 410153 309464 417423
rect 309784 410508 310424 417068
rect 274624 347508 275264 354068
rect 275584 347153 276224 354423
rect 286024 347153 286664 354423
rect 286984 347153 287624 354423
rect 297424 347153 298064 354423
rect 298384 347153 299024 354423
rect 308824 347153 309464 354423
rect 309784 347508 310424 354068
rect 274624 284508 275264 291068
rect 275584 284153 276224 291423
rect 286024 284153 286664 291423
rect 286984 284153 287624 291423
rect 297424 284153 298064 291423
rect 298384 284153 299024 291423
rect 308824 284153 309464 291423
rect 309784 284508 310424 291068
rect 274624 221508 275264 228068
rect 275584 221153 276224 228423
rect 286024 221153 286664 228423
rect 286984 221153 287624 228423
rect 297424 221153 298064 228423
rect 298384 221153 299024 228423
rect 308824 221153 309464 228423
rect 309784 221508 310424 228068
rect 274624 158508 275264 165068
rect 275584 158153 276224 165423
rect 286024 158153 286664 165423
rect 286984 158153 287624 165423
rect 297424 158153 298064 165423
rect 298384 158153 299024 165423
rect 308824 158153 309464 165423
rect 309784 158508 310424 165068
rect 274624 95508 275264 102068
rect 275584 95153 276224 102423
rect 286024 95153 286664 102423
rect 286984 95153 287624 102423
rect 297424 95153 298064 102423
rect 298384 95153 299024 102423
rect 308824 95153 309464 102423
rect 309784 95508 310424 102068
rect 274624 32588 275264 39068
rect 274624 -744 275264 6068
rect 275584 -744 276224 39423
rect 286024 32233 286664 39423
rect 286984 32233 287624 39423
rect 297424 32233 298064 39423
rect 298384 32233 299024 39423
rect 286024 -744 286664 10639
rect 286984 -744 287624 10639
rect 297424 -744 298064 10639
rect 298384 -744 299024 10639
rect 308824 -744 309464 39423
rect 309784 32588 310424 39068
rect 309784 -744 310424 6068
rect 320224 -744 320864 543656
rect 321184 -744 321824 543656
rect 331624 536508 332264 543656
rect 332584 535609 333224 543656
rect 343024 535609 343664 543656
rect 343984 535609 344624 543656
rect 354424 535609 355064 543656
rect 355384 535609 356024 543656
rect 365824 535609 366464 543656
rect 366784 536508 367424 543656
rect 331624 473508 332264 480068
rect 332584 473153 333224 480423
rect 343024 473153 343664 480423
rect 343984 473153 344624 480423
rect 354424 473153 355064 480423
rect 355384 473153 356024 480423
rect 365824 473153 366464 480423
rect 366784 473508 367424 480068
rect 331624 410508 332264 417068
rect 332584 410153 333224 417423
rect 343024 410153 343664 417423
rect 343984 410153 344624 417423
rect 354424 410153 355064 417423
rect 355384 410153 356024 417423
rect 365824 410153 366464 417423
rect 366784 410508 367424 417068
rect 331624 347508 332264 354068
rect 332584 347153 333224 354423
rect 343024 347153 343664 354423
rect 343984 347153 344624 354423
rect 354424 347153 355064 354423
rect 355384 347153 356024 354423
rect 365824 347153 366464 354423
rect 366784 347508 367424 354068
rect 331624 284508 332264 291068
rect 332584 284153 333224 291423
rect 343024 284153 343664 291423
rect 343984 284153 344624 291423
rect 354424 284153 355064 291423
rect 355384 284153 356024 291423
rect 365824 284153 366464 291423
rect 366784 284508 367424 291068
rect 331624 221508 332264 228068
rect 332584 221153 333224 228423
rect 343024 221153 343664 228423
rect 343984 221153 344624 228423
rect 354424 221153 355064 228423
rect 355384 221153 356024 228423
rect 365824 221153 366464 228423
rect 366784 221508 367424 228068
rect 331624 158508 332264 165068
rect 332584 158153 333224 165423
rect 343024 158153 343664 165423
rect 343984 158153 344624 165423
rect 354424 158153 355064 165423
rect 355384 158153 356024 165423
rect 365824 158153 366464 165423
rect 366784 158508 367424 165068
rect 331624 95508 332264 102068
rect 332584 95153 333224 102423
rect 343024 95153 343664 102423
rect 343984 95153 344624 102423
rect 354424 95153 355064 102423
rect 355384 95153 356024 102423
rect 365824 95153 366464 102423
rect 366784 95508 367424 102068
rect 331624 32588 332264 39068
rect 331624 -744 332264 6068
rect 332584 -744 333224 39423
rect 343024 32233 343664 39423
rect 343984 32233 344624 39423
rect 354424 32233 355064 39423
rect 355384 32233 356024 39423
rect 343024 -744 343664 10639
rect 343984 -744 344624 10639
rect 354424 -744 355064 10639
rect 355384 -744 356024 10639
rect 365824 -744 366464 39423
rect 366784 32588 367424 39068
rect 366784 -744 367424 6068
rect 377224 -744 377864 543656
rect 378184 -744 378824 543656
rect 388624 536508 389264 543656
rect 389584 535609 390224 543656
rect 400024 535609 400664 543656
rect 400984 535609 401624 543656
rect 411424 535609 412064 543656
rect 412384 535609 413024 543656
rect 422824 535609 423464 543656
rect 423784 536508 424424 543656
rect 388624 473508 389264 480068
rect 389584 473153 390224 480423
rect 400024 473153 400664 480423
rect 400984 473153 401624 480423
rect 411424 473153 412064 480423
rect 412384 473153 413024 480423
rect 422824 473153 423464 480423
rect 423784 473508 424424 480068
rect 388624 410508 389264 417068
rect 389584 410153 390224 417423
rect 400024 410153 400664 417423
rect 400984 410153 401624 417423
rect 411424 410153 412064 417423
rect 412384 410153 413024 417423
rect 422824 410153 423464 417423
rect 423784 410508 424424 417068
rect 388624 347508 389264 354068
rect 389584 347153 390224 354423
rect 400024 347153 400664 354423
rect 400984 347153 401624 354423
rect 411424 347153 412064 354423
rect 412384 347153 413024 354423
rect 422824 347153 423464 354423
rect 423784 347508 424424 354068
rect 388624 284508 389264 291068
rect 389584 284153 390224 291423
rect 400024 284153 400664 291423
rect 400984 284153 401624 291423
rect 411424 284153 412064 291423
rect 412384 284153 413024 291423
rect 422824 284153 423464 291423
rect 423784 284508 424424 291068
rect 388624 221508 389264 228068
rect 389584 221153 390224 228423
rect 400024 221153 400664 228423
rect 400984 221153 401624 228423
rect 411424 221153 412064 228423
rect 412384 221153 413024 228423
rect 422824 221153 423464 228423
rect 423784 221508 424424 228068
rect 388624 158508 389264 165068
rect 389584 158153 390224 165423
rect 400024 158153 400664 165423
rect 400984 158153 401624 165423
rect 411424 158153 412064 165423
rect 412384 158153 413024 165423
rect 422824 158153 423464 165423
rect 423784 158508 424424 165068
rect 388624 95508 389264 102068
rect 389584 95153 390224 102423
rect 400024 95153 400664 102423
rect 400984 95153 401624 102423
rect 411424 95153 412064 102423
rect 412384 95153 413024 102423
rect 422824 95153 423464 102423
rect 423784 95508 424424 102068
rect 388624 32588 389264 39068
rect 388624 -744 389264 6068
rect 389584 -744 390224 39423
rect 400024 32233 400664 39423
rect 400984 32233 401624 39423
rect 411424 32233 412064 39423
rect 412384 32233 413024 39423
rect 400024 -744 400664 10639
rect 400984 -744 401624 10639
rect 411424 -744 412064 10639
rect 412384 -744 413024 10639
rect 422824 -744 423464 39423
rect 423784 32588 424424 39068
rect 423784 -744 424424 6068
rect 434224 -744 434864 543656
rect 435184 -744 435824 543656
rect 445624 536508 446264 543656
rect 446584 535473 447224 543656
rect 457024 535473 457664 543656
rect 457984 535473 458624 543656
rect 468424 535473 469064 543656
rect 469384 535473 470024 543656
rect 479824 535473 480464 543656
rect 480784 536508 481424 543656
rect 445624 473508 446264 480068
rect 446584 471657 447224 481375
rect 457024 471657 457664 481375
rect 457984 471657 458624 481375
rect 468424 471657 469064 481375
rect 469384 471657 470024 481375
rect 479824 471657 480464 481375
rect 480784 473508 481424 480068
rect 445624 410508 446264 417068
rect 446584 408657 447224 418919
rect 457024 408657 457664 418919
rect 457984 408657 458624 418919
rect 468424 408657 469064 418919
rect 469384 408657 470024 418919
rect 479824 408657 480464 418919
rect 480784 410508 481424 417068
rect 445624 347508 446264 354068
rect 446584 345657 447224 355919
rect 457024 345657 457664 355919
rect 457984 345657 458624 355919
rect 468424 345657 469064 355919
rect 469384 345657 470024 355919
rect 479824 345657 480464 355919
rect 480784 347508 481424 354068
rect 445624 284508 446264 291068
rect 446584 282657 447224 292919
rect 457024 282657 457664 292919
rect 457984 282657 458624 292919
rect 468424 282657 469064 292919
rect 469384 282657 470024 292919
rect 479824 282657 480464 292919
rect 480784 284508 481424 291068
rect 445624 221508 446264 228068
rect 446584 219657 447224 229919
rect 457024 219657 457664 229919
rect 457984 219657 458624 229919
rect 468424 219657 469064 229919
rect 469384 219657 470024 229919
rect 479824 219657 480464 229919
rect 480784 221508 481424 228068
rect 445624 158508 446264 165068
rect 446584 156657 447224 166919
rect 457024 156657 457664 166919
rect 457984 156657 458624 166919
rect 468424 156657 469064 166919
rect 469384 156657 470024 166919
rect 479824 156657 480464 166919
rect 480784 158508 481424 165068
rect 445624 95508 446264 102068
rect 446584 93657 447224 103919
rect 457024 93657 457664 103919
rect 457984 93657 458624 103919
rect 468424 93657 469064 103919
rect 469384 93657 470024 103919
rect 479824 93657 480464 103919
rect 480784 95508 481424 102068
rect 445624 33049 446264 39068
rect 446584 33049 447224 40919
rect 457024 33049 457664 40919
rect 457984 33049 458624 40919
rect 468424 33049 469064 40919
rect 469384 33049 470024 40919
rect 445624 -744 446264 6068
rect 446584 -744 447224 11183
rect 457024 -744 457664 11183
rect 457984 -744 458624 11183
rect 468424 -744 469064 11183
rect 469384 -744 470024 11183
rect 479824 -744 480464 40919
rect 480784 32588 481424 39068
rect 480784 -744 481424 6068
rect 491224 -744 491864 543656
rect 492184 -744 492824 543656
rect 495192 616 496152 542296
rect 496552 -744 497512 543656
<< obsm4 >>
rect 8267 471577 12344 534448
rect 13144 520841 24704 534448
rect 25504 520841 35144 534448
rect 13144 481455 35144 520841
rect 13144 480148 24704 481455
rect 13144 473428 13304 480148
rect 14104 473428 23744 480148
rect 24544 473428 24704 480148
rect 13144 471577 24704 473428
rect 25504 471577 35144 481455
rect 8267 418999 35144 471577
rect 8267 408577 12344 418999
rect 13144 417148 24704 418999
rect 13144 410428 13304 417148
rect 14104 410428 23744 417148
rect 24544 410428 24704 417148
rect 13144 408577 24704 410428
rect 25504 408577 35144 418999
rect 8267 355999 35144 408577
rect 8267 345577 12344 355999
rect 13144 354148 24704 355999
rect 13144 347428 13304 354148
rect 14104 347428 23744 354148
rect 24544 347428 24704 354148
rect 13144 345577 24704 347428
rect 25504 345577 35144 355999
rect 8267 292999 35144 345577
rect 8267 282577 12344 292999
rect 13144 291148 24704 292999
rect 13144 284428 13304 291148
rect 14104 284428 23744 291148
rect 24544 284428 24704 291148
rect 13144 282577 24704 284428
rect 25504 282577 35144 292999
rect 8267 229999 35144 282577
rect 8267 219577 12344 229999
rect 13144 228148 24704 229999
rect 13144 221428 13304 228148
rect 14104 221428 23744 228148
rect 24544 221428 24704 228148
rect 13144 219577 24704 221428
rect 25504 219577 35144 229999
rect 8267 166999 35144 219577
rect 8267 156577 12344 166999
rect 13144 165148 24704 166999
rect 13144 158428 13304 165148
rect 14104 158428 23744 165148
rect 24544 158428 24704 165148
rect 13144 156577 24704 158428
rect 25504 156577 35144 166999
rect 8267 103999 35144 156577
rect 8267 93577 12344 103999
rect 13144 102148 24704 103999
rect 13144 95428 13304 102148
rect 14104 95428 23744 102148
rect 24544 95428 24704 102148
rect 13144 93577 24704 95428
rect 25504 93577 35144 103999
rect 8267 40999 35144 93577
rect 8267 34329 12344 40999
rect 13144 39148 24704 40999
rect 13144 34329 13304 39148
rect 14104 34329 23744 39148
rect 24544 34329 24704 39148
rect 25504 34329 35144 40999
rect 8267 12351 35144 34329
rect 8267 8128 12344 12351
rect 13144 8128 24704 12351
rect 25504 8128 35144 12351
rect 35944 8128 36104 534448
rect 36904 480503 92144 534448
rect 36904 480148 47504 480503
rect 36904 473428 46544 480148
rect 47344 473428 47504 480148
rect 36904 473073 47504 473428
rect 48304 473073 57944 480503
rect 58744 473073 58904 480503
rect 59704 473073 69344 480503
rect 70144 473073 70304 480503
rect 71104 473073 80744 480503
rect 81544 480148 92144 480503
rect 81544 473428 81704 480148
rect 82504 473428 92144 480148
rect 81544 473073 92144 473428
rect 36904 417503 92144 473073
rect 36904 417148 47504 417503
rect 36904 410428 46544 417148
rect 47344 410428 47504 417148
rect 36904 410073 47504 410428
rect 48304 410073 57944 417503
rect 58744 410073 58904 417503
rect 59704 410073 69344 417503
rect 70144 410073 70304 417503
rect 71104 410073 80744 417503
rect 81544 417148 92144 417503
rect 81544 410428 81704 417148
rect 82504 410428 92144 417148
rect 81544 410073 92144 410428
rect 36904 354503 92144 410073
rect 36904 354148 47504 354503
rect 36904 347428 46544 354148
rect 47344 347428 47504 354148
rect 36904 347073 47504 347428
rect 48304 347073 57944 354503
rect 58744 347073 58904 354503
rect 59704 347073 69344 354503
rect 70144 347073 70304 354503
rect 71104 347073 80744 354503
rect 81544 354148 92144 354503
rect 81544 347428 81704 354148
rect 82504 347428 92144 354148
rect 81544 347073 92144 347428
rect 36904 291503 92144 347073
rect 36904 291148 47504 291503
rect 36904 284428 46544 291148
rect 47344 284428 47504 291148
rect 36904 284073 47504 284428
rect 48304 284073 57944 291503
rect 58744 284073 58904 291503
rect 59704 284073 69344 291503
rect 70144 284073 70304 291503
rect 71104 284073 80744 291503
rect 81544 291148 92144 291503
rect 81544 284428 81704 291148
rect 82504 284428 92144 291148
rect 81544 284073 92144 284428
rect 36904 228503 92144 284073
rect 36904 228148 47504 228503
rect 36904 221428 46544 228148
rect 47344 221428 47504 228148
rect 36904 221073 47504 221428
rect 48304 221073 57944 228503
rect 58744 221073 58904 228503
rect 59704 221073 69344 228503
rect 70144 221073 70304 228503
rect 71104 221073 80744 228503
rect 81544 228148 92144 228503
rect 81544 221428 81704 228148
rect 82504 221428 92144 228148
rect 81544 221073 92144 221428
rect 36904 165503 92144 221073
rect 36904 165148 47504 165503
rect 36904 158428 46544 165148
rect 47344 158428 47504 165148
rect 36904 158073 47504 158428
rect 48304 158073 57944 165503
rect 58744 158073 58904 165503
rect 59704 158073 69344 165503
rect 70144 158073 70304 165503
rect 71104 158073 80744 165503
rect 81544 165148 92144 165503
rect 81544 158428 81704 165148
rect 82504 158428 92144 165148
rect 81544 158073 92144 158428
rect 36904 102503 92144 158073
rect 36904 102148 47504 102503
rect 36904 95428 46544 102148
rect 47344 95428 47504 102148
rect 36904 95073 47504 95428
rect 48304 95073 57944 102503
rect 58744 95073 58904 102503
rect 59704 95073 69344 102503
rect 70144 95073 70304 102503
rect 71104 95073 80744 102503
rect 81544 102148 92144 102503
rect 81544 95428 81704 102148
rect 82504 95428 92144 102148
rect 81544 95073 92144 95428
rect 36904 39503 92144 95073
rect 36904 39148 47504 39503
rect 36904 32508 46544 39148
rect 47344 32508 47504 39148
rect 36904 8128 47504 32508
rect 48304 32153 57944 39503
rect 58744 32153 58904 39503
rect 59704 32153 69344 39503
rect 70144 32153 70304 39503
rect 71104 32153 80744 39503
rect 48304 10719 80744 32153
rect 48304 8128 57944 10719
rect 58744 8128 58904 10719
rect 59704 8128 69344 10719
rect 70144 8128 70304 10719
rect 71104 8128 80744 10719
rect 81544 39148 92144 39503
rect 81544 32508 81704 39148
rect 82504 32508 92144 39148
rect 81544 8128 92144 32508
rect 92944 8128 93104 534448
rect 93904 480503 149144 534448
rect 93904 480148 104504 480503
rect 93904 473428 103544 480148
rect 104344 473428 104504 480148
rect 93904 473073 104504 473428
rect 105304 473073 114944 480503
rect 115744 473073 115904 480503
rect 116704 473073 126344 480503
rect 127144 473073 127304 480503
rect 128104 473073 137744 480503
rect 138544 480148 149144 480503
rect 138544 473428 138704 480148
rect 139504 473428 149144 480148
rect 138544 473073 149144 473428
rect 93904 417503 149144 473073
rect 93904 417148 104504 417503
rect 93904 410428 103544 417148
rect 104344 410428 104504 417148
rect 93904 410073 104504 410428
rect 105304 410073 114944 417503
rect 115744 410073 115904 417503
rect 116704 410073 126344 417503
rect 127144 410073 127304 417503
rect 128104 410073 137744 417503
rect 138544 417148 149144 417503
rect 138544 410428 138704 417148
rect 139504 410428 149144 417148
rect 138544 410073 149144 410428
rect 93904 354503 149144 410073
rect 93904 354148 104504 354503
rect 93904 347428 103544 354148
rect 104344 347428 104504 354148
rect 93904 347073 104504 347428
rect 105304 347073 114944 354503
rect 115744 347073 115904 354503
rect 116704 347073 126344 354503
rect 127144 347073 127304 354503
rect 128104 347073 137744 354503
rect 138544 354148 149144 354503
rect 138544 347428 138704 354148
rect 139504 347428 149144 354148
rect 138544 347073 149144 347428
rect 93904 291503 149144 347073
rect 93904 291148 104504 291503
rect 93904 284428 103544 291148
rect 104344 284428 104504 291148
rect 93904 284073 104504 284428
rect 105304 284073 114944 291503
rect 115744 284073 115904 291503
rect 116704 284073 126344 291503
rect 127144 284073 127304 291503
rect 128104 284073 137744 291503
rect 138544 291148 149144 291503
rect 138544 284428 138704 291148
rect 139504 284428 149144 291148
rect 138544 284073 149144 284428
rect 93904 228503 149144 284073
rect 93904 228148 104504 228503
rect 93904 221428 103544 228148
rect 104344 221428 104504 228148
rect 93904 221073 104504 221428
rect 105304 221073 114944 228503
rect 115744 221073 115904 228503
rect 116704 221073 126344 228503
rect 127144 221073 127304 228503
rect 128104 221073 137744 228503
rect 138544 228148 149144 228503
rect 138544 221428 138704 228148
rect 139504 221428 149144 228148
rect 138544 221073 149144 221428
rect 93904 165503 149144 221073
rect 93904 165148 104504 165503
rect 93904 158428 103544 165148
rect 104344 158428 104504 165148
rect 93904 158073 104504 158428
rect 105304 158073 114944 165503
rect 115744 158073 115904 165503
rect 116704 158073 126344 165503
rect 127144 158073 127304 165503
rect 128104 158073 137744 165503
rect 138544 165148 149144 165503
rect 138544 158428 138704 165148
rect 139504 158428 149144 165148
rect 138544 158073 149144 158428
rect 93904 102503 149144 158073
rect 93904 102148 104504 102503
rect 93904 95428 103544 102148
rect 104344 95428 104504 102148
rect 93904 95073 104504 95428
rect 105304 95073 114944 102503
rect 115744 95073 115904 102503
rect 116704 95073 126344 102503
rect 127144 95073 127304 102503
rect 128104 95073 137744 102503
rect 138544 102148 149144 102503
rect 138544 95428 138704 102148
rect 139504 95428 149144 102148
rect 138544 95073 149144 95428
rect 93904 39503 149144 95073
rect 93904 39148 104504 39503
rect 93904 32508 103544 39148
rect 104344 32508 104504 39148
rect 93904 8128 104504 32508
rect 105304 32153 114944 39503
rect 115744 32153 115904 39503
rect 116704 32153 126344 39503
rect 127144 32153 127304 39503
rect 128104 32153 137744 39503
rect 105304 10719 137744 32153
rect 105304 8128 114944 10719
rect 115744 8128 115904 10719
rect 116704 8128 126344 10719
rect 127144 8128 127304 10719
rect 128104 8128 137744 10719
rect 138544 39148 149144 39503
rect 138544 32508 138704 39148
rect 139504 32508 149144 39148
rect 138544 8128 149144 32508
rect 149944 8128 150104 534448
rect 150904 480503 206144 534448
rect 150904 480148 161504 480503
rect 150904 473428 160544 480148
rect 161344 473428 161504 480148
rect 150904 473073 161504 473428
rect 162304 473073 171944 480503
rect 172744 473073 172904 480503
rect 173704 473073 183344 480503
rect 184144 473073 184304 480503
rect 185104 473073 194744 480503
rect 195544 480148 206144 480503
rect 195544 473428 195704 480148
rect 196504 473428 206144 480148
rect 195544 473073 206144 473428
rect 150904 417503 206144 473073
rect 150904 417148 161504 417503
rect 150904 410428 160544 417148
rect 161344 410428 161504 417148
rect 150904 410073 161504 410428
rect 162304 410073 171944 417503
rect 172744 410073 172904 417503
rect 173704 410073 183344 417503
rect 184144 410073 184304 417503
rect 185104 410073 194744 417503
rect 195544 417148 206144 417503
rect 195544 410428 195704 417148
rect 196504 410428 206144 417148
rect 195544 410073 206144 410428
rect 150904 354503 206144 410073
rect 150904 354148 161504 354503
rect 150904 347428 160544 354148
rect 161344 347428 161504 354148
rect 150904 347073 161504 347428
rect 162304 347073 171944 354503
rect 172744 347073 172904 354503
rect 173704 347073 183344 354503
rect 184144 347073 184304 354503
rect 185104 347073 194744 354503
rect 195544 354148 206144 354503
rect 195544 347428 195704 354148
rect 196504 347428 206144 354148
rect 195544 347073 206144 347428
rect 150904 291503 206144 347073
rect 150904 291148 161504 291503
rect 150904 284428 160544 291148
rect 161344 284428 161504 291148
rect 150904 284073 161504 284428
rect 162304 284073 171944 291503
rect 172744 284073 172904 291503
rect 173704 284073 183344 291503
rect 184144 284073 184304 291503
rect 185104 284073 194744 291503
rect 195544 291148 206144 291503
rect 195544 284428 195704 291148
rect 196504 284428 206144 291148
rect 195544 284073 206144 284428
rect 150904 228503 206144 284073
rect 150904 228148 161504 228503
rect 150904 221428 160544 228148
rect 161344 221428 161504 228148
rect 150904 221073 161504 221428
rect 162304 221073 171944 228503
rect 172744 221073 172904 228503
rect 173704 221073 183344 228503
rect 184144 221073 184304 228503
rect 185104 221073 194744 228503
rect 195544 228148 206144 228503
rect 195544 221428 195704 228148
rect 196504 221428 206144 228148
rect 195544 221073 206144 221428
rect 150904 165503 206144 221073
rect 150904 165148 161504 165503
rect 150904 158428 160544 165148
rect 161344 158428 161504 165148
rect 150904 158073 161504 158428
rect 162304 158073 171944 165503
rect 172744 158073 172904 165503
rect 173704 158073 183344 165503
rect 184144 158073 184304 165503
rect 185104 158073 194744 165503
rect 195544 165148 206144 165503
rect 195544 158428 195704 165148
rect 196504 158428 206144 165148
rect 195544 158073 206144 158428
rect 150904 102503 206144 158073
rect 150904 102148 161504 102503
rect 150904 95428 160544 102148
rect 161344 95428 161504 102148
rect 150904 95073 161504 95428
rect 162304 95073 171944 102503
rect 172744 95073 172904 102503
rect 173704 95073 183344 102503
rect 184144 95073 184304 102503
rect 185104 95073 194744 102503
rect 195544 102148 206144 102503
rect 195544 95428 195704 102148
rect 196504 95428 206144 102148
rect 195544 95073 206144 95428
rect 150904 39503 206144 95073
rect 150904 39148 161504 39503
rect 150904 32508 160544 39148
rect 161344 32508 161504 39148
rect 150904 8128 161504 32508
rect 162304 32153 171944 39503
rect 172744 32153 172904 39503
rect 173704 32153 183344 39503
rect 184144 32153 184304 39503
rect 185104 32153 194744 39503
rect 162304 10719 194744 32153
rect 162304 8128 171944 10719
rect 172744 8128 172904 10719
rect 173704 8128 183344 10719
rect 184144 8128 184304 10719
rect 185104 8128 194744 10719
rect 195544 39148 206144 39503
rect 195544 32508 195704 39148
rect 196504 32508 206144 39148
rect 195544 8128 206144 32508
rect 206944 8128 207104 534448
rect 207904 480503 263144 534448
rect 207904 480148 218504 480503
rect 207904 473428 217544 480148
rect 218344 473428 218504 480148
rect 207904 473073 218504 473428
rect 219304 473073 228944 480503
rect 229744 473073 229904 480503
rect 230704 473073 240344 480503
rect 241144 473073 241304 480503
rect 242104 473073 251744 480503
rect 252544 480148 263144 480503
rect 252544 473428 252704 480148
rect 253504 473428 263144 480148
rect 252544 473073 263144 473428
rect 207904 417503 263144 473073
rect 207904 417148 218504 417503
rect 207904 410428 217544 417148
rect 218344 410428 218504 417148
rect 207904 410073 218504 410428
rect 219304 410073 228944 417503
rect 229744 410073 229904 417503
rect 230704 410073 240344 417503
rect 241144 410073 241304 417503
rect 242104 410073 251744 417503
rect 252544 417148 263144 417503
rect 252544 410428 252704 417148
rect 253504 410428 263144 417148
rect 252544 410073 263144 410428
rect 207904 354503 263144 410073
rect 207904 354148 218504 354503
rect 207904 347428 217544 354148
rect 218344 347428 218504 354148
rect 207904 347073 218504 347428
rect 219304 347073 228944 354503
rect 229744 347073 229904 354503
rect 230704 347073 240344 354503
rect 241144 347073 241304 354503
rect 242104 347073 251744 354503
rect 252544 354148 263144 354503
rect 252544 347428 252704 354148
rect 253504 347428 263144 354148
rect 252544 347073 263144 347428
rect 207904 291503 263144 347073
rect 207904 291148 218504 291503
rect 207904 284428 217544 291148
rect 218344 284428 218504 291148
rect 207904 284073 218504 284428
rect 219304 284073 228944 291503
rect 229744 284073 229904 291503
rect 230704 284073 240344 291503
rect 241144 284073 241304 291503
rect 242104 284073 251744 291503
rect 252544 291148 263144 291503
rect 252544 284428 252704 291148
rect 253504 284428 263144 291148
rect 252544 284073 263144 284428
rect 207904 228503 263144 284073
rect 207904 228148 218504 228503
rect 207904 221428 217544 228148
rect 218344 221428 218504 228148
rect 207904 221073 218504 221428
rect 219304 221073 228944 228503
rect 229744 221073 229904 228503
rect 230704 221073 240344 228503
rect 241144 221073 241304 228503
rect 242104 221073 251744 228503
rect 252544 228148 263144 228503
rect 252544 221428 252704 228148
rect 253504 221428 263144 228148
rect 252544 221073 263144 221428
rect 207904 165503 263144 221073
rect 207904 165148 218504 165503
rect 207904 158428 217544 165148
rect 218344 158428 218504 165148
rect 207904 158073 218504 158428
rect 219304 158073 228944 165503
rect 229744 158073 229904 165503
rect 230704 158073 240344 165503
rect 241144 158073 241304 165503
rect 242104 158073 251744 165503
rect 252544 165148 263144 165503
rect 252544 158428 252704 165148
rect 253504 158428 263144 165148
rect 252544 158073 263144 158428
rect 207904 102503 263144 158073
rect 207904 102148 218504 102503
rect 207904 95428 217544 102148
rect 218344 95428 218504 102148
rect 207904 95073 218504 95428
rect 219304 95073 228944 102503
rect 229744 95073 229904 102503
rect 230704 95073 240344 102503
rect 241144 95073 241304 102503
rect 242104 95073 251744 102503
rect 252544 102148 263144 102503
rect 252544 95428 252704 102148
rect 253504 95428 263144 102148
rect 252544 95073 263144 95428
rect 207904 39503 263144 95073
rect 207904 39148 218504 39503
rect 207904 32508 217544 39148
rect 218344 32508 218504 39148
rect 207904 8128 218504 32508
rect 219304 32153 228944 39503
rect 229744 32153 229904 39503
rect 230704 32153 240344 39503
rect 241144 32153 241304 39503
rect 242104 32153 251744 39503
rect 219304 10719 251744 32153
rect 219304 8128 228944 10719
rect 229744 8128 229904 10719
rect 230704 8128 240344 10719
rect 241144 8128 241304 10719
rect 242104 8128 251744 10719
rect 252544 39148 263144 39503
rect 252544 32508 252704 39148
rect 253504 32508 263144 39148
rect 252544 8128 263144 32508
rect 263944 8128 264104 534448
rect 264904 480503 320144 534448
rect 264904 480148 275504 480503
rect 264904 473428 274544 480148
rect 275344 473428 275504 480148
rect 264904 473073 275504 473428
rect 276304 473073 285944 480503
rect 286744 473073 286904 480503
rect 287704 473073 297344 480503
rect 298144 473073 298304 480503
rect 299104 473073 308744 480503
rect 309544 480148 320144 480503
rect 309544 473428 309704 480148
rect 310504 473428 320144 480148
rect 309544 473073 320144 473428
rect 264904 417503 320144 473073
rect 264904 417148 275504 417503
rect 264904 410428 274544 417148
rect 275344 410428 275504 417148
rect 264904 410073 275504 410428
rect 276304 410073 285944 417503
rect 286744 410073 286904 417503
rect 287704 410073 297344 417503
rect 298144 410073 298304 417503
rect 299104 410073 308744 417503
rect 309544 417148 320144 417503
rect 309544 410428 309704 417148
rect 310504 410428 320144 417148
rect 309544 410073 320144 410428
rect 264904 354503 320144 410073
rect 264904 354148 275504 354503
rect 264904 347428 274544 354148
rect 275344 347428 275504 354148
rect 264904 347073 275504 347428
rect 276304 347073 285944 354503
rect 286744 347073 286904 354503
rect 287704 347073 297344 354503
rect 298144 347073 298304 354503
rect 299104 347073 308744 354503
rect 309544 354148 320144 354503
rect 309544 347428 309704 354148
rect 310504 347428 320144 354148
rect 309544 347073 320144 347428
rect 264904 291503 320144 347073
rect 264904 291148 275504 291503
rect 264904 284428 274544 291148
rect 275344 284428 275504 291148
rect 264904 284073 275504 284428
rect 276304 284073 285944 291503
rect 286744 284073 286904 291503
rect 287704 284073 297344 291503
rect 298144 284073 298304 291503
rect 299104 284073 308744 291503
rect 309544 291148 320144 291503
rect 309544 284428 309704 291148
rect 310504 284428 320144 291148
rect 309544 284073 320144 284428
rect 264904 228503 320144 284073
rect 264904 228148 275504 228503
rect 264904 221428 274544 228148
rect 275344 221428 275504 228148
rect 264904 221073 275504 221428
rect 276304 221073 285944 228503
rect 286744 221073 286904 228503
rect 287704 221073 297344 228503
rect 298144 221073 298304 228503
rect 299104 221073 308744 228503
rect 309544 228148 320144 228503
rect 309544 221428 309704 228148
rect 310504 221428 320144 228148
rect 309544 221073 320144 221428
rect 264904 165503 320144 221073
rect 264904 165148 275504 165503
rect 264904 158428 274544 165148
rect 275344 158428 275504 165148
rect 264904 158073 275504 158428
rect 276304 158073 285944 165503
rect 286744 158073 286904 165503
rect 287704 158073 297344 165503
rect 298144 158073 298304 165503
rect 299104 158073 308744 165503
rect 309544 165148 320144 165503
rect 309544 158428 309704 165148
rect 310504 158428 320144 165148
rect 309544 158073 320144 158428
rect 264904 102503 320144 158073
rect 264904 102148 275504 102503
rect 264904 95428 274544 102148
rect 275344 95428 275504 102148
rect 264904 95073 275504 95428
rect 276304 95073 285944 102503
rect 286744 95073 286904 102503
rect 287704 95073 297344 102503
rect 298144 95073 298304 102503
rect 299104 95073 308744 102503
rect 309544 102148 320144 102503
rect 309544 95428 309704 102148
rect 310504 95428 320144 102148
rect 309544 95073 320144 95428
rect 264904 39503 320144 95073
rect 264904 39148 275504 39503
rect 264904 32508 274544 39148
rect 275344 32508 275504 39148
rect 264904 8128 275504 32508
rect 276304 32153 285944 39503
rect 286744 32153 286904 39503
rect 287704 32153 297344 39503
rect 298144 32153 298304 39503
rect 299104 32153 308744 39503
rect 276304 10719 308744 32153
rect 276304 8128 285944 10719
rect 286744 8128 286904 10719
rect 287704 8128 297344 10719
rect 298144 8128 298304 10719
rect 299104 8128 308744 10719
rect 309544 39148 320144 39503
rect 309544 32508 309704 39148
rect 310504 32508 320144 39148
rect 309544 8128 320144 32508
rect 320944 8128 321104 534448
rect 321904 480503 377144 534448
rect 321904 480148 332504 480503
rect 321904 473428 331544 480148
rect 332344 473428 332504 480148
rect 321904 473073 332504 473428
rect 333304 473073 342944 480503
rect 343744 473073 343904 480503
rect 344704 473073 354344 480503
rect 355144 473073 355304 480503
rect 356104 473073 365744 480503
rect 366544 480148 377144 480503
rect 366544 473428 366704 480148
rect 367504 473428 377144 480148
rect 366544 473073 377144 473428
rect 321904 417503 377144 473073
rect 321904 417148 332504 417503
rect 321904 410428 331544 417148
rect 332344 410428 332504 417148
rect 321904 410073 332504 410428
rect 333304 410073 342944 417503
rect 343744 410073 343904 417503
rect 344704 410073 354344 417503
rect 355144 410073 355304 417503
rect 356104 410073 365744 417503
rect 366544 417148 377144 417503
rect 366544 410428 366704 417148
rect 367504 410428 377144 417148
rect 366544 410073 377144 410428
rect 321904 354503 377144 410073
rect 321904 354148 332504 354503
rect 321904 347428 331544 354148
rect 332344 347428 332504 354148
rect 321904 347073 332504 347428
rect 333304 347073 342944 354503
rect 343744 347073 343904 354503
rect 344704 347073 354344 354503
rect 355144 347073 355304 354503
rect 356104 347073 365744 354503
rect 366544 354148 377144 354503
rect 366544 347428 366704 354148
rect 367504 347428 377144 354148
rect 366544 347073 377144 347428
rect 321904 291503 377144 347073
rect 321904 291148 332504 291503
rect 321904 284428 331544 291148
rect 332344 284428 332504 291148
rect 321904 284073 332504 284428
rect 333304 284073 342944 291503
rect 343744 284073 343904 291503
rect 344704 284073 354344 291503
rect 355144 284073 355304 291503
rect 356104 284073 365744 291503
rect 366544 291148 377144 291503
rect 366544 284428 366704 291148
rect 367504 284428 377144 291148
rect 366544 284073 377144 284428
rect 321904 228503 377144 284073
rect 321904 228148 332504 228503
rect 321904 221428 331544 228148
rect 332344 221428 332504 228148
rect 321904 221073 332504 221428
rect 333304 221073 342944 228503
rect 343744 221073 343904 228503
rect 344704 221073 354344 228503
rect 355144 221073 355304 228503
rect 356104 221073 365744 228503
rect 366544 228148 377144 228503
rect 366544 221428 366704 228148
rect 367504 221428 377144 228148
rect 366544 221073 377144 221428
rect 321904 165503 377144 221073
rect 321904 165148 332504 165503
rect 321904 158428 331544 165148
rect 332344 158428 332504 165148
rect 321904 158073 332504 158428
rect 333304 158073 342944 165503
rect 343744 158073 343904 165503
rect 344704 158073 354344 165503
rect 355144 158073 355304 165503
rect 356104 158073 365744 165503
rect 366544 165148 377144 165503
rect 366544 158428 366704 165148
rect 367504 158428 377144 165148
rect 366544 158073 377144 158428
rect 321904 102503 377144 158073
rect 321904 102148 332504 102503
rect 321904 95428 331544 102148
rect 332344 95428 332504 102148
rect 321904 95073 332504 95428
rect 333304 95073 342944 102503
rect 343744 95073 343904 102503
rect 344704 95073 354344 102503
rect 355144 95073 355304 102503
rect 356104 95073 365744 102503
rect 366544 102148 377144 102503
rect 366544 95428 366704 102148
rect 367504 95428 377144 102148
rect 366544 95073 377144 95428
rect 321904 39503 377144 95073
rect 321904 39148 332504 39503
rect 321904 32508 331544 39148
rect 332344 32508 332504 39148
rect 321904 8128 332504 32508
rect 333304 32153 342944 39503
rect 343744 32153 343904 39503
rect 344704 32153 354344 39503
rect 355144 32153 355304 39503
rect 356104 32153 365744 39503
rect 333304 10719 365744 32153
rect 333304 8128 342944 10719
rect 343744 8128 343904 10719
rect 344704 8128 354344 10719
rect 355144 8128 355304 10719
rect 356104 8128 365744 10719
rect 366544 39148 377144 39503
rect 366544 32508 366704 39148
rect 367504 32508 377144 39148
rect 366544 8128 377144 32508
rect 377944 8128 378104 534448
rect 378904 480503 434144 534448
rect 378904 480148 389504 480503
rect 378904 473428 388544 480148
rect 389344 473428 389504 480148
rect 378904 473073 389504 473428
rect 390304 473073 399944 480503
rect 400744 473073 400904 480503
rect 401704 473073 411344 480503
rect 412144 473073 412304 480503
rect 413104 473073 422744 480503
rect 423544 480148 434144 480503
rect 423544 473428 423704 480148
rect 424504 473428 434144 480148
rect 423544 473073 434144 473428
rect 378904 417503 434144 473073
rect 378904 417148 389504 417503
rect 378904 410428 388544 417148
rect 389344 410428 389504 417148
rect 378904 410073 389504 410428
rect 390304 410073 399944 417503
rect 400744 410073 400904 417503
rect 401704 410073 411344 417503
rect 412144 410073 412304 417503
rect 413104 410073 422744 417503
rect 423544 417148 434144 417503
rect 423544 410428 423704 417148
rect 424504 410428 434144 417148
rect 423544 410073 434144 410428
rect 378904 354503 434144 410073
rect 378904 354148 389504 354503
rect 378904 347428 388544 354148
rect 389344 347428 389504 354148
rect 378904 347073 389504 347428
rect 390304 347073 399944 354503
rect 400744 347073 400904 354503
rect 401704 347073 411344 354503
rect 412144 347073 412304 354503
rect 413104 347073 422744 354503
rect 423544 354148 434144 354503
rect 423544 347428 423704 354148
rect 424504 347428 434144 354148
rect 423544 347073 434144 347428
rect 378904 291503 434144 347073
rect 378904 291148 389504 291503
rect 378904 284428 388544 291148
rect 389344 284428 389504 291148
rect 378904 284073 389504 284428
rect 390304 284073 399944 291503
rect 400744 284073 400904 291503
rect 401704 284073 411344 291503
rect 412144 284073 412304 291503
rect 413104 284073 422744 291503
rect 423544 291148 434144 291503
rect 423544 284428 423704 291148
rect 424504 284428 434144 291148
rect 423544 284073 434144 284428
rect 378904 228503 434144 284073
rect 378904 228148 389504 228503
rect 378904 221428 388544 228148
rect 389344 221428 389504 228148
rect 378904 221073 389504 221428
rect 390304 221073 399944 228503
rect 400744 221073 400904 228503
rect 401704 221073 411344 228503
rect 412144 221073 412304 228503
rect 413104 221073 422744 228503
rect 423544 228148 434144 228503
rect 423544 221428 423704 228148
rect 424504 221428 434144 228148
rect 423544 221073 434144 221428
rect 378904 165503 434144 221073
rect 378904 165148 389504 165503
rect 378904 158428 388544 165148
rect 389344 158428 389504 165148
rect 378904 158073 389504 158428
rect 390304 158073 399944 165503
rect 400744 158073 400904 165503
rect 401704 158073 411344 165503
rect 412144 158073 412304 165503
rect 413104 158073 422744 165503
rect 423544 165148 434144 165503
rect 423544 158428 423704 165148
rect 424504 158428 434144 165148
rect 423544 158073 434144 158428
rect 378904 102503 434144 158073
rect 378904 102148 389504 102503
rect 378904 95428 388544 102148
rect 389344 95428 389504 102148
rect 378904 95073 389504 95428
rect 390304 95073 399944 102503
rect 400744 95073 400904 102503
rect 401704 95073 411344 102503
rect 412144 95073 412304 102503
rect 413104 95073 422744 102503
rect 423544 102148 434144 102503
rect 423544 95428 423704 102148
rect 424504 95428 434144 102148
rect 423544 95073 434144 95428
rect 378904 39503 434144 95073
rect 378904 39148 389504 39503
rect 378904 32508 388544 39148
rect 389344 32508 389504 39148
rect 378904 8128 389504 32508
rect 390304 32153 399944 39503
rect 400744 32153 400904 39503
rect 401704 32153 411344 39503
rect 412144 32153 412304 39503
rect 413104 32153 422744 39503
rect 390304 10719 422744 32153
rect 390304 8128 399944 10719
rect 400744 8128 400904 10719
rect 401704 8128 411344 10719
rect 412144 8128 412304 10719
rect 413104 8128 422744 10719
rect 423544 39148 434144 39503
rect 423544 32508 423704 39148
rect 424504 32508 434144 39148
rect 423544 8128 434144 32508
rect 434944 8128 435104 534448
rect 435904 481455 486264 534448
rect 435904 480148 446504 481455
rect 435904 473428 445544 480148
rect 446344 473428 446504 480148
rect 435904 471577 446504 473428
rect 447304 471577 456944 481455
rect 457744 471577 457904 481455
rect 458704 471577 468344 481455
rect 469144 471577 469304 481455
rect 470104 471577 479744 481455
rect 480544 480148 486264 481455
rect 480544 473428 480704 480148
rect 481504 473428 486264 480148
rect 480544 471577 486264 473428
rect 435904 418999 486264 471577
rect 435904 417148 446504 418999
rect 435904 410428 445544 417148
rect 446344 410428 446504 417148
rect 435904 408577 446504 410428
rect 447304 408577 456944 418999
rect 457744 408577 457904 418999
rect 458704 408577 468344 418999
rect 469144 408577 469304 418999
rect 470104 408577 479744 418999
rect 480544 417148 486264 418999
rect 480544 410428 480704 417148
rect 481504 410428 486264 417148
rect 480544 408577 486264 410428
rect 435904 355999 486264 408577
rect 435904 354148 446504 355999
rect 435904 347428 445544 354148
rect 446344 347428 446504 354148
rect 435904 345577 446504 347428
rect 447304 345577 456944 355999
rect 457744 345577 457904 355999
rect 458704 345577 468344 355999
rect 469144 345577 469304 355999
rect 470104 345577 479744 355999
rect 480544 354148 486264 355999
rect 480544 347428 480704 354148
rect 481504 347428 486264 354148
rect 480544 345577 486264 347428
rect 435904 292999 486264 345577
rect 435904 291148 446504 292999
rect 435904 284428 445544 291148
rect 446344 284428 446504 291148
rect 435904 282577 446504 284428
rect 447304 282577 456944 292999
rect 457744 282577 457904 292999
rect 458704 282577 468344 292999
rect 469144 282577 469304 292999
rect 470104 282577 479744 292999
rect 480544 291148 486264 292999
rect 480544 284428 480704 291148
rect 481504 284428 486264 291148
rect 480544 282577 486264 284428
rect 435904 229999 486264 282577
rect 435904 228148 446504 229999
rect 435904 221428 445544 228148
rect 446344 221428 446504 228148
rect 435904 219577 446504 221428
rect 447304 219577 456944 229999
rect 457744 219577 457904 229999
rect 458704 219577 468344 229999
rect 469144 219577 469304 229999
rect 470104 219577 479744 229999
rect 480544 228148 486264 229999
rect 480544 221428 480704 228148
rect 481504 221428 486264 228148
rect 480544 219577 486264 221428
rect 435904 166999 486264 219577
rect 435904 165148 446504 166999
rect 435904 158428 445544 165148
rect 446344 158428 446504 165148
rect 435904 156577 446504 158428
rect 447304 156577 456944 166999
rect 457744 156577 457904 166999
rect 458704 156577 468344 166999
rect 469144 156577 469304 166999
rect 470104 156577 479744 166999
rect 480544 165148 486264 166999
rect 480544 158428 480704 165148
rect 481504 158428 486264 165148
rect 480544 156577 486264 158428
rect 435904 103999 486264 156577
rect 435904 102148 446504 103999
rect 435904 95428 445544 102148
rect 446344 95428 446504 102148
rect 435904 93577 446504 95428
rect 447304 93577 456944 103999
rect 457744 93577 457904 103999
rect 458704 93577 468344 103999
rect 469144 93577 469304 103999
rect 470104 93577 479744 103999
rect 480544 102148 486264 103999
rect 480544 95428 480704 102148
rect 481504 95428 486264 102148
rect 480544 93577 486264 95428
rect 435904 40999 486264 93577
rect 435904 39148 446504 40999
rect 435904 32969 445544 39148
rect 446344 32969 446504 39148
rect 447304 32969 456944 40999
rect 457744 32969 457904 40999
rect 458704 32969 468344 40999
rect 469144 32969 469304 40999
rect 470104 32969 479744 40999
rect 435904 11263 479744 32969
rect 435904 8128 446504 11263
rect 447304 8128 456944 11263
rect 457744 8128 457904 11263
rect 458704 8128 468344 11263
rect 469144 8128 469304 11263
rect 470104 8128 479744 11263
rect 480544 39148 486264 40999
rect 480544 32508 480704 39148
rect 481504 32508 486264 39148
rect 480544 8128 486264 32508
<< metal5 >>
rect -2552 542696 497512 543656
rect -1192 541336 496152 542296
rect -2552 539356 497512 539996
rect -2552 530136 497512 530776
rect -2552 528856 497512 529496
rect -2552 519636 497512 520276
rect -2552 518356 497512 518996
rect -2552 509136 497512 509776
rect -2552 507856 497512 508496
rect -2552 498636 497512 499276
rect -2552 497356 497512 497996
rect -2552 488136 497512 488776
rect -2552 486856 497512 487496
rect -2552 477636 497512 478276
rect -2552 476356 497512 476996
rect -2552 467136 497512 467776
rect -2552 465856 497512 466496
rect -2552 456636 497512 457276
rect -2552 455356 497512 455996
rect -2552 446136 497512 446776
rect -2552 444856 497512 445496
rect -2552 435636 497512 436276
rect -2552 434356 497512 434996
rect -2552 425136 497512 425776
rect -2552 423856 497512 424496
rect -2552 414636 497512 415276
rect -2552 413356 497512 413996
rect -2552 404136 497512 404776
rect -2552 402856 497512 403496
rect -2552 393636 497512 394276
rect -2552 392356 497512 392996
rect -2552 383136 497512 383776
rect -2552 381856 497512 382496
rect -2552 372636 497512 373276
rect -2552 371356 497512 371996
rect -2552 362136 497512 362776
rect -2552 360856 497512 361496
rect -2552 351636 497512 352276
rect -2552 350356 497512 350996
rect -2552 341136 497512 341776
rect -2552 339856 497512 340496
rect -2552 330636 497512 331276
rect -2552 329356 497512 329996
rect -2552 320136 497512 320776
rect -2552 318856 497512 319496
rect -2552 309636 497512 310276
rect -2552 308356 497512 308996
rect -2552 299136 497512 299776
rect -2552 297856 497512 298496
rect -2552 288636 497512 289276
rect -2552 287356 497512 287996
rect -2552 278136 497512 278776
rect -2552 276856 497512 277496
rect -2552 267636 497512 268276
rect -2552 266356 497512 266996
rect -2552 257136 497512 257776
rect -2552 255856 497512 256496
rect -2552 246636 497512 247276
rect -2552 245356 497512 245996
rect -2552 236136 497512 236776
rect -2552 234856 497512 235496
rect -2552 225636 497512 226276
rect -2552 224356 497512 224996
rect -2552 215136 497512 215776
rect -2552 213856 497512 214496
rect -2552 204636 497512 205276
rect -2552 203356 497512 203996
rect -2552 194136 497512 194776
rect -2552 192856 497512 193496
rect -2552 183636 497512 184276
rect -2552 182356 497512 182996
rect -2552 173136 497512 173776
rect -2552 171856 497512 172496
rect -2552 162636 497512 163276
rect -2552 161356 497512 161996
rect -2552 152136 497512 152776
rect -2552 150856 497512 151496
rect -2552 141636 497512 142276
rect -2552 140356 497512 140996
rect -2552 131136 497512 131776
rect -2552 129856 497512 130496
rect -2552 120636 497512 121276
rect -2552 119356 497512 119996
rect -2552 110136 497512 110776
rect -2552 108856 497512 109496
rect -2552 99636 497512 100276
rect -2552 98356 497512 98996
rect -2552 89136 497512 89776
rect -2552 87856 497512 88496
rect -2552 78636 497512 79276
rect -2552 77356 497512 77996
rect -2552 68136 497512 68776
rect -2552 66856 497512 67496
rect -2552 57636 497512 58276
rect -2552 56356 497512 56996
rect -2552 47136 497512 47776
rect -2552 45856 497512 46496
rect -2552 36636 497512 37276
rect -2552 35356 497512 35996
rect -2552 26136 497512 26776
rect -2552 24856 497512 25496
rect -2552 15636 497512 16276
rect -2552 14356 497512 14996
rect -2552 5136 497512 5776
rect -2552 3856 497512 4496
rect -1192 616 496152 1576
rect -2552 -744 497512 216
<< labels >>
rlabel metal4 s -2552 -744 -1592 543656 4 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 -744 497512 216 8 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 542696 497512 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 496552 -744 497512 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1984 -744 2624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 -744 14024 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 34409 14024 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 95508 14024 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 158508 14024 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 221508 14024 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 284508 14024 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 347508 14024 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 410508 14024 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 473508 14024 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13384 536508 14024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 -744 25424 12271 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 34409 25424 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 93657 25424 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 156657 25424 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 219657 25424 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 282657 25424 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 345657 25424 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 408657 25424 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 471657 25424 481375 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 24784 520921 25424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 36184 -744 36824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 -744 48224 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 95153 48224 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 158153 48224 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 221153 48224 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 284153 48224 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 347153 48224 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 410153 48224 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 473153 48224 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47584 535609 48224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 -744 59624 10639 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 32233 59624 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 95153 59624 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 158153 59624 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 221153 59624 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 284153 59624 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 347153 59624 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 410153 59624 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 473153 59624 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 58984 535609 59624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 -744 71024 10639 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 32233 71024 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 95153 71024 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 158153 71024 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 221153 71024 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 284153 71024 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 347153 71024 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 410153 71024 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 473153 71024 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 70384 535609 71024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 -744 82424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 32588 82424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 95508 82424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 158508 82424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 221508 82424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 284508 82424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 347508 82424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 410508 82424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 473508 82424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81784 536508 82424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 93184 -744 93824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 -744 105224 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 95153 105224 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 158153 105224 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 221153 105224 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 284153 105224 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 347153 105224 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 410153 105224 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 473153 105224 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 104584 535609 105224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 -744 116624 10639 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 32233 116624 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 95153 116624 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 158153 116624 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 221153 116624 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 284153 116624 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 347153 116624 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 410153 116624 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 473153 116624 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 115984 535609 116624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 -744 128024 10639 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 32233 128024 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 95153 128024 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 158153 128024 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 221153 128024 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 284153 128024 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 347153 128024 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 410153 128024 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 473153 128024 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 127384 535609 128024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 -744 139424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 32588 139424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 95508 139424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 158508 139424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 221508 139424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 284508 139424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 347508 139424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 410508 139424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 473508 139424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 138784 536508 139424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 150184 -744 150824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 -744 162224 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 95153 162224 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 158153 162224 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 221153 162224 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 284153 162224 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 347153 162224 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 410153 162224 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 473153 162224 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 161584 535609 162224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 -744 173624 10639 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 32233 173624 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 95153 173624 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 158153 173624 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 221153 173624 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 284153 173624 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 347153 173624 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 410153 173624 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 473153 173624 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 172984 535609 173624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 -744 185024 10639 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 32233 185024 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 95153 185024 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 158153 185024 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 221153 185024 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 284153 185024 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 347153 185024 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 410153 185024 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 473153 185024 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 184384 535609 185024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 -744 196424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 32588 196424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 95508 196424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 158508 196424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 221508 196424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 284508 196424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 347508 196424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 410508 196424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 473508 196424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 195784 536508 196424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 207184 -744 207824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 -744 219224 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 95153 219224 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 158153 219224 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 221153 219224 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 284153 219224 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 347153 219224 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 410153 219224 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 473153 219224 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 218584 535609 219224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 -744 230624 10639 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 32233 230624 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 95153 230624 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 158153 230624 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 221153 230624 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 284153 230624 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 347153 230624 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 410153 230624 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 473153 230624 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 229984 535609 230624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 -744 242024 10639 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 32233 242024 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 95153 242024 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 158153 242024 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 221153 242024 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 284153 242024 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 347153 242024 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 410153 242024 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 473153 242024 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 241384 535609 242024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 -744 253424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 32588 253424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 95508 253424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 158508 253424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 221508 253424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 284508 253424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 347508 253424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 410508 253424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 473508 253424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 252784 536508 253424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 264184 -744 264824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 -744 276224 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 95153 276224 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 158153 276224 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 221153 276224 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 284153 276224 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 347153 276224 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 410153 276224 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 473153 276224 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 275584 535609 276224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 -744 287624 10639 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 32233 287624 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 95153 287624 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 158153 287624 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 221153 287624 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 284153 287624 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 347153 287624 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 410153 287624 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 473153 287624 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 286984 535609 287624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 -744 299024 10639 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 32233 299024 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 95153 299024 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 158153 299024 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 221153 299024 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 284153 299024 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 347153 299024 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 410153 299024 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 473153 299024 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 298384 535609 299024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 -744 310424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 32588 310424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 95508 310424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 158508 310424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 221508 310424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 284508 310424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 347508 310424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 410508 310424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 473508 310424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 309784 536508 310424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 321184 -744 321824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 -744 333224 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 95153 333224 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 158153 333224 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 221153 333224 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 284153 333224 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 347153 333224 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 410153 333224 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 473153 333224 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 332584 535609 333224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 -744 344624 10639 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 32233 344624 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 95153 344624 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 158153 344624 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 221153 344624 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 284153 344624 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 347153 344624 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 410153 344624 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 473153 344624 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 343984 535609 344624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 -744 356024 10639 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 32233 356024 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 95153 356024 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 158153 356024 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 221153 356024 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 284153 356024 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 347153 356024 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 410153 356024 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 473153 356024 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 355384 535609 356024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 -744 367424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 32588 367424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 95508 367424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 158508 367424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 221508 367424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 284508 367424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 347508 367424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 410508 367424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 473508 367424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 366784 536508 367424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 378184 -744 378824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 -744 390224 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 95153 390224 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 158153 390224 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 221153 390224 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 284153 390224 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 347153 390224 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 410153 390224 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 473153 390224 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 389584 535609 390224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 -744 401624 10639 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 32233 401624 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 95153 401624 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 158153 401624 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 221153 401624 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 284153 401624 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 347153 401624 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 410153 401624 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 473153 401624 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 400984 535609 401624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 -744 413024 10639 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 32233 413024 39423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 95153 413024 102423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 158153 413024 165423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 221153 413024 228423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 284153 413024 291423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 347153 413024 354423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 410153 413024 417423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 473153 413024 480423 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 412384 535609 413024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 -744 424424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 32588 424424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 95508 424424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 158508 424424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 221508 424424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 284508 424424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 347508 424424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 410508 424424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 473508 424424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 423784 536508 424424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 435184 -744 435824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 -744 447224 11183 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 33049 447224 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 93657 447224 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 156657 447224 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 219657 447224 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 282657 447224 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 345657 447224 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 408657 447224 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 471657 447224 481375 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 446584 535473 447224 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 -744 458624 11183 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 33049 458624 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 93657 458624 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 156657 458624 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 219657 458624 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 282657 458624 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 345657 458624 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 408657 458624 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 471657 458624 481375 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 457984 535473 458624 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 -744 470024 11183 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 33049 470024 40919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 93657 470024 103919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 156657 470024 166919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 219657 470024 229919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 282657 470024 292919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 345657 470024 355919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 408657 470024 418919 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 471657 470024 481375 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 469384 535473 470024 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 -744 481424 6068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 32588 481424 39068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 95508 481424 102068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 158508 481424 165068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 221508 481424 228068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 284508 481424 291068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 347508 481424 354068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 410508 481424 417068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 473508 481424 480068 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 480784 536508 481424 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 492184 -744 492824 543656 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 5136 497512 5776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 15636 497512 16276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 26136 497512 26776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 36636 497512 37276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 47136 497512 47776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 57636 497512 58276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 68136 497512 68776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 78636 497512 79276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 89136 497512 89776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 99636 497512 100276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 110136 497512 110776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 120636 497512 121276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 131136 497512 131776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 141636 497512 142276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 152136 497512 152776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 162636 497512 163276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 173136 497512 173776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 183636 497512 184276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 194136 497512 194776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 204636 497512 205276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 215136 497512 215776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 225636 497512 226276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 236136 497512 236776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 246636 497512 247276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 257136 497512 257776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 267636 497512 268276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 278136 497512 278776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 288636 497512 289276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 299136 497512 299776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 309636 497512 310276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 320136 497512 320776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 330636 497512 331276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 341136 497512 341776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 351636 497512 352276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 362136 497512 362776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 372636 497512 373276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 383136 497512 383776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 393636 497512 394276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 404136 497512 404776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 414636 497512 415276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 425136 497512 425776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 435636 497512 436276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 446136 497512 446776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 456636 497512 457276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 467136 497512 467776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 477636 497512 478276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 488136 497512 488776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 498636 497512 499276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 509136 497512 509776 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 519636 497512 520276 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s -2552 530136 497512 530776 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s -1192 616 -232 542296 4 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -1192 616 496152 1576 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -1192 541336 496152 542296 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 495192 616 496152 542296 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 1024 -744 1664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12424 -744 13064 12271 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12424 34409 13064 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12424 93657 13064 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12424 156657 13064 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12424 219657 13064 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12424 282657 13064 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12424 345657 13064 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12424 408657 13064 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12424 471657 13064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 -744 24464 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 34409 24464 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 95508 24464 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 158508 24464 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 221508 24464 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 284508 24464 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 347508 24464 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 410508 24464 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 473508 24464 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 23824 536508 24464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 35224 -744 35864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 -744 47264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 32588 47264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 95508 47264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 158508 47264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 221508 47264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 284508 47264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 347508 47264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 410508 47264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 473508 47264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 46624 536508 47264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 -744 58664 10639 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 32233 58664 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 95153 58664 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 158153 58664 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 221153 58664 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 284153 58664 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 347153 58664 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 410153 58664 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 473153 58664 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 58024 535609 58664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 -744 70064 10639 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 32233 70064 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 95153 70064 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 158153 70064 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 221153 70064 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 284153 70064 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 347153 70064 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 410153 70064 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 473153 70064 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 69424 535609 70064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 -744 81464 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 95153 81464 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 158153 81464 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 221153 81464 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 284153 81464 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 347153 81464 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 410153 81464 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 473153 81464 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 80824 535609 81464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 92224 -744 92864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 -744 104264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 32588 104264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 95508 104264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 158508 104264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 221508 104264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 284508 104264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 347508 104264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 410508 104264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 473508 104264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 103624 536508 104264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 -744 115664 10639 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 32233 115664 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 95153 115664 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 158153 115664 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 221153 115664 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 284153 115664 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 347153 115664 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 410153 115664 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 473153 115664 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 115024 535609 115664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 -744 127064 10639 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 32233 127064 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 95153 127064 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 158153 127064 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 221153 127064 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 284153 127064 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 347153 127064 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 410153 127064 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 473153 127064 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 126424 535609 127064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 -744 138464 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 95153 138464 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 158153 138464 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 221153 138464 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 284153 138464 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 347153 138464 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 410153 138464 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 473153 138464 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 137824 535609 138464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 149224 -744 149864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 -744 161264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 32588 161264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 95508 161264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 158508 161264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 221508 161264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 284508 161264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 347508 161264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 410508 161264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 473508 161264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 160624 536508 161264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 -744 172664 10639 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 32233 172664 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 95153 172664 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 158153 172664 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 221153 172664 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 284153 172664 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 347153 172664 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 410153 172664 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 473153 172664 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 172024 535609 172664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 -744 184064 10639 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 32233 184064 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 95153 184064 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 158153 184064 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 221153 184064 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 284153 184064 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 347153 184064 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 410153 184064 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 473153 184064 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 183424 535609 184064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 -744 195464 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 95153 195464 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 158153 195464 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 221153 195464 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 284153 195464 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 347153 195464 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 410153 195464 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 473153 195464 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 194824 535609 195464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 206224 -744 206864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 -744 218264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 32588 218264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 95508 218264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 158508 218264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 221508 218264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 284508 218264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 347508 218264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 410508 218264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 473508 218264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 217624 536508 218264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 -744 229664 10639 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 32233 229664 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 95153 229664 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 158153 229664 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 221153 229664 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 284153 229664 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 347153 229664 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 410153 229664 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 473153 229664 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 229024 535609 229664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 -744 241064 10639 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 32233 241064 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 95153 241064 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 158153 241064 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 221153 241064 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 284153 241064 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 347153 241064 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 410153 241064 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 473153 241064 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 240424 535609 241064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 -744 252464 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 95153 252464 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 158153 252464 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 221153 252464 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 284153 252464 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 347153 252464 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 410153 252464 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 473153 252464 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 251824 535609 252464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 263224 -744 263864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 -744 275264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 32588 275264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 95508 275264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 158508 275264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 221508 275264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 284508 275264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 347508 275264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 410508 275264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 473508 275264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 274624 536508 275264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 -744 286664 10639 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 32233 286664 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 95153 286664 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 158153 286664 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 221153 286664 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 284153 286664 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 347153 286664 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 410153 286664 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 473153 286664 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 286024 535609 286664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 -744 298064 10639 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 32233 298064 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 95153 298064 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 158153 298064 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 221153 298064 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 284153 298064 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 347153 298064 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 410153 298064 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 473153 298064 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 297424 535609 298064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 -744 309464 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 95153 309464 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 158153 309464 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 221153 309464 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 284153 309464 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 347153 309464 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 410153 309464 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 473153 309464 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 308824 535609 309464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 320224 -744 320864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 -744 332264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 32588 332264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 95508 332264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 158508 332264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 221508 332264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 284508 332264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 347508 332264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 410508 332264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 473508 332264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 331624 536508 332264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 -744 343664 10639 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 32233 343664 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 95153 343664 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 158153 343664 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 221153 343664 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 284153 343664 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 347153 343664 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 410153 343664 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 473153 343664 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 343024 535609 343664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 -744 355064 10639 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 32233 355064 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 95153 355064 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 158153 355064 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 221153 355064 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 284153 355064 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 347153 355064 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 410153 355064 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 473153 355064 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 354424 535609 355064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 -744 366464 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 95153 366464 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 158153 366464 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 221153 366464 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 284153 366464 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 347153 366464 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 410153 366464 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 473153 366464 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 365824 535609 366464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 377224 -744 377864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 -744 389264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 32588 389264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 95508 389264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 158508 389264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 221508 389264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 284508 389264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 347508 389264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 410508 389264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 473508 389264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 388624 536508 389264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 -744 400664 10639 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 32233 400664 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 95153 400664 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 158153 400664 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 221153 400664 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 284153 400664 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 347153 400664 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 410153 400664 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 473153 400664 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 400024 535609 400664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 -744 412064 10639 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 32233 412064 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 95153 412064 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 158153 412064 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 221153 412064 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 284153 412064 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 347153 412064 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 410153 412064 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 473153 412064 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 411424 535609 412064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 -744 423464 39423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 95153 423464 102423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 158153 423464 165423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 221153 423464 228423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 284153 423464 291423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 347153 423464 354423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 410153 423464 417423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 473153 423464 480423 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 422824 535609 423464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 434224 -744 434864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 -744 446264 6068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 33049 446264 39068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 95508 446264 102068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 158508 446264 165068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 221508 446264 228068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 284508 446264 291068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 347508 446264 354068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 410508 446264 417068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 473508 446264 480068 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 445624 536508 446264 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 -744 457664 11183 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 33049 457664 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 93657 457664 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 156657 457664 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 219657 457664 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 282657 457664 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 345657 457664 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 408657 457664 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 471657 457664 481375 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 457024 535473 457664 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 -744 469064 11183 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 33049 469064 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 93657 469064 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 156657 469064 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 219657 469064 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 282657 469064 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 345657 469064 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 408657 469064 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 471657 469064 481375 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 468424 535473 469064 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 -744 480464 40919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 93657 480464 103919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 156657 480464 166919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 219657 480464 229919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 282657 480464 292919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 345657 480464 355919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 408657 480464 418919 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 471657 480464 481375 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 479824 535473 480464 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 491224 -744 491864 543656 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 3856 497512 4496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 14356 497512 14996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 24856 497512 25496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 35356 497512 35996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 45856 497512 46496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 56356 497512 56996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 66856 497512 67496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 77356 497512 77996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 87856 497512 88496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 98356 497512 98996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 108856 497512 109496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 119356 497512 119996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 129856 497512 130496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 140356 497512 140996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 150856 497512 151496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 161356 497512 161996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 171856 497512 172496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 182356 497512 182996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 192856 497512 193496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 203356 497512 203996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 213856 497512 214496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 224356 497512 224996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 234856 497512 235496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 245356 497512 245996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 255856 497512 256496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 266356 497512 266996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 276856 497512 277496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 287356 497512 287996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 297856 497512 298496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 308356 497512 308996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 318856 497512 319496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 329356 497512 329996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 339856 497512 340496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 350356 497512 350996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 360856 497512 361496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 371356 497512 371996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 381856 497512 382496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 392356 497512 392996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 402856 497512 403496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 413356 497512 413996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 423856 497512 424496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 434356 497512 434996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 444856 497512 445496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 455356 497512 455996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 465856 497512 466496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 476356 497512 476996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 486856 497512 487496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 497356 497512 497996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 507856 497512 508496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 518356 497512 518996 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 528856 497512 529496 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s -2552 539356 497512 539996 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 73526 0 73582 800 6 ccff_head
port 3 nsew signal input
rlabel metal2 s 59726 542200 59782 543000 6 ccff_tail
port 4 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 clk
port 5 nsew signal input
rlabel metal2 s 15566 542200 15622 543000 6 gfpga_pad_io_soc_dir[0]
port 6 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 gfpga_pad_io_soc_dir[100]
port 7 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 gfpga_pad_io_soc_dir[101]
port 8 nsew signal output
rlabel metal3 s 0 124448 800 124568 6 gfpga_pad_io_soc_dir[102]
port 9 nsew signal output
rlabel metal3 s 0 140768 800 140888 6 gfpga_pad_io_soc_dir[103]
port 10 nsew signal output
rlabel metal3 s 0 157088 800 157208 6 gfpga_pad_io_soc_dir[104]
port 11 nsew signal output
rlabel metal3 s 0 173408 800 173528 6 gfpga_pad_io_soc_dir[105]
port 12 nsew signal output
rlabel metal3 s 0 189728 800 189848 6 gfpga_pad_io_soc_dir[106]
port 13 nsew signal output
rlabel metal3 s 0 206048 800 206168 6 gfpga_pad_io_soc_dir[107]
port 14 nsew signal output
rlabel metal3 s 0 222368 800 222488 6 gfpga_pad_io_soc_dir[108]
port 15 nsew signal output
rlabel metal3 s 0 238688 800 238808 6 gfpga_pad_io_soc_dir[109]
port 16 nsew signal output
rlabel metal2 s 156878 542200 156934 543000 6 gfpga_pad_io_soc_dir[10]
port 17 nsew signal output
rlabel metal3 s 0 255008 800 255128 6 gfpga_pad_io_soc_dir[110]
port 18 nsew signal output
rlabel metal3 s 0 276768 800 276888 6 gfpga_pad_io_soc_dir[111]
port 19 nsew signal output
rlabel metal3 s 0 293088 800 293208 6 gfpga_pad_io_soc_dir[112]
port 20 nsew signal output
rlabel metal3 s 0 309408 800 309528 6 gfpga_pad_io_soc_dir[113]
port 21 nsew signal output
rlabel metal3 s 0 325728 800 325848 6 gfpga_pad_io_soc_dir[114]
port 22 nsew signal output
rlabel metal3 s 0 342048 800 342168 6 gfpga_pad_io_soc_dir[115]
port 23 nsew signal output
rlabel metal3 s 0 358368 800 358488 6 gfpga_pad_io_soc_dir[116]
port 24 nsew signal output
rlabel metal3 s 0 374688 800 374808 6 gfpga_pad_io_soc_dir[117]
port 25 nsew signal output
rlabel metal3 s 0 391008 800 391128 6 gfpga_pad_io_soc_dir[118]
port 26 nsew signal output
rlabel metal3 s 0 407328 800 407448 6 gfpga_pad_io_soc_dir[119]
port 27 nsew signal output
rlabel metal2 s 170126 542200 170182 543000 6 gfpga_pad_io_soc_dir[11]
port 28 nsew signal output
rlabel metal3 s 0 423648 800 423768 6 gfpga_pad_io_soc_dir[120]
port 29 nsew signal output
rlabel metal3 s 0 439968 800 440088 6 gfpga_pad_io_soc_dir[121]
port 30 nsew signal output
rlabel metal3 s 0 456288 800 456408 6 gfpga_pad_io_soc_dir[122]
port 31 nsew signal output
rlabel metal3 s 0 472608 800 472728 6 gfpga_pad_io_soc_dir[123]
port 32 nsew signal output
rlabel metal3 s 0 488928 800 489048 6 gfpga_pad_io_soc_dir[124]
port 33 nsew signal output
rlabel metal3 s 0 505248 800 505368 6 gfpga_pad_io_soc_dir[125]
port 34 nsew signal output
rlabel metal3 s 0 521568 800 521688 6 gfpga_pad_io_soc_dir[126]
port 35 nsew signal output
rlabel metal3 s 0 537888 800 538008 6 gfpga_pad_io_soc_dir[127]
port 36 nsew signal output
rlabel metal2 s 183374 542200 183430 543000 6 gfpga_pad_io_soc_dir[12]
port 37 nsew signal output
rlabel metal2 s 196622 542200 196678 543000 6 gfpga_pad_io_soc_dir[13]
port 38 nsew signal output
rlabel metal2 s 209870 542200 209926 543000 6 gfpga_pad_io_soc_dir[14]
port 39 nsew signal output
rlabel metal2 s 223118 542200 223174 543000 6 gfpga_pad_io_soc_dir[15]
port 40 nsew signal output
rlabel metal2 s 236366 542200 236422 543000 6 gfpga_pad_io_soc_dir[16]
port 41 nsew signal output
rlabel metal2 s 249614 542200 249670 543000 6 gfpga_pad_io_soc_dir[17]
port 42 nsew signal output
rlabel metal2 s 262862 542200 262918 543000 6 gfpga_pad_io_soc_dir[18]
port 43 nsew signal output
rlabel metal2 s 276110 542200 276166 543000 6 gfpga_pad_io_soc_dir[19]
port 44 nsew signal output
rlabel metal2 s 28814 542200 28870 543000 6 gfpga_pad_io_soc_dir[1]
port 45 nsew signal output
rlabel metal2 s 289358 542200 289414 543000 6 gfpga_pad_io_soc_dir[20]
port 46 nsew signal output
rlabel metal2 s 302606 542200 302662 543000 6 gfpga_pad_io_soc_dir[21]
port 47 nsew signal output
rlabel metal2 s 315854 542200 315910 543000 6 gfpga_pad_io_soc_dir[22]
port 48 nsew signal output
rlabel metal2 s 329102 542200 329158 543000 6 gfpga_pad_io_soc_dir[23]
port 49 nsew signal output
rlabel metal2 s 342350 542200 342406 543000 6 gfpga_pad_io_soc_dir[24]
port 50 nsew signal output
rlabel metal2 s 355598 542200 355654 543000 6 gfpga_pad_io_soc_dir[25]
port 51 nsew signal output
rlabel metal2 s 368846 542200 368902 543000 6 gfpga_pad_io_soc_dir[26]
port 52 nsew signal output
rlabel metal2 s 382094 542200 382150 543000 6 gfpga_pad_io_soc_dir[27]
port 53 nsew signal output
rlabel metal2 s 395342 542200 395398 543000 6 gfpga_pad_io_soc_dir[28]
port 54 nsew signal output
rlabel metal2 s 408590 542200 408646 543000 6 gfpga_pad_io_soc_dir[29]
port 55 nsew signal output
rlabel metal2 s 42062 542200 42118 543000 6 gfpga_pad_io_soc_dir[2]
port 56 nsew signal output
rlabel metal2 s 421838 542200 421894 543000 6 gfpga_pad_io_soc_dir[30]
port 57 nsew signal output
rlabel metal2 s 435086 542200 435142 543000 6 gfpga_pad_io_soc_dir[31]
port 58 nsew signal output
rlabel metal2 s 448334 542200 448390 543000 6 gfpga_pad_io_soc_dir[32]
port 59 nsew signal output
rlabel metal2 s 461582 542200 461638 543000 6 gfpga_pad_io_soc_dir[33]
port 60 nsew signal output
rlabel metal2 s 474830 542200 474886 543000 6 gfpga_pad_io_soc_dir[34]
port 61 nsew signal output
rlabel metal2 s 488078 542200 488134 543000 6 gfpga_pad_io_soc_dir[35]
port 62 nsew signal output
rlabel metal3 s 494200 518032 495000 518152 6 gfpga_pad_io_soc_dir[36]
port 63 nsew signal output
rlabel metal3 s 494200 502120 495000 502240 6 gfpga_pad_io_soc_dir[37]
port 64 nsew signal output
rlabel metal3 s 494200 486208 495000 486328 6 gfpga_pad_io_soc_dir[38]
port 65 nsew signal output
rlabel metal3 s 494200 470296 495000 470416 6 gfpga_pad_io_soc_dir[39]
port 66 nsew signal output
rlabel metal2 s 55310 542200 55366 543000 6 gfpga_pad_io_soc_dir[3]
port 67 nsew signal output
rlabel metal3 s 494200 454384 495000 454504 6 gfpga_pad_io_soc_dir[40]
port 68 nsew signal output
rlabel metal3 s 494200 438472 495000 438592 6 gfpga_pad_io_soc_dir[41]
port 69 nsew signal output
rlabel metal3 s 494200 422560 495000 422680 6 gfpga_pad_io_soc_dir[42]
port 70 nsew signal output
rlabel metal3 s 494200 406648 495000 406768 6 gfpga_pad_io_soc_dir[43]
port 71 nsew signal output
rlabel metal3 s 494200 390736 495000 390856 6 gfpga_pad_io_soc_dir[44]
port 72 nsew signal output
rlabel metal3 s 494200 374824 495000 374944 6 gfpga_pad_io_soc_dir[45]
port 73 nsew signal output
rlabel metal3 s 494200 358912 495000 359032 6 gfpga_pad_io_soc_dir[46]
port 74 nsew signal output
rlabel metal3 s 494200 343000 495000 343120 6 gfpga_pad_io_soc_dir[47]
port 75 nsew signal output
rlabel metal3 s 494200 327088 495000 327208 6 gfpga_pad_io_soc_dir[48]
port 76 nsew signal output
rlabel metal3 s 494200 311176 495000 311296 6 gfpga_pad_io_soc_dir[49]
port 77 nsew signal output
rlabel metal2 s 77390 542200 77446 543000 6 gfpga_pad_io_soc_dir[4]
port 78 nsew signal output
rlabel metal3 s 494200 295264 495000 295384 6 gfpga_pad_io_soc_dir[50]
port 79 nsew signal output
rlabel metal3 s 494200 279352 495000 279472 6 gfpga_pad_io_soc_dir[51]
port 80 nsew signal output
rlabel metal3 s 494200 263440 495000 263560 6 gfpga_pad_io_soc_dir[52]
port 81 nsew signal output
rlabel metal3 s 494200 247528 495000 247648 6 gfpga_pad_io_soc_dir[53]
port 82 nsew signal output
rlabel metal3 s 494200 221008 495000 221128 6 gfpga_pad_io_soc_dir[54]
port 83 nsew signal output
rlabel metal3 s 494200 205096 495000 205216 6 gfpga_pad_io_soc_dir[55]
port 84 nsew signal output
rlabel metal3 s 494200 189184 495000 189304 6 gfpga_pad_io_soc_dir[56]
port 85 nsew signal output
rlabel metal3 s 494200 173272 495000 173392 6 gfpga_pad_io_soc_dir[57]
port 86 nsew signal output
rlabel metal3 s 494200 157360 495000 157480 6 gfpga_pad_io_soc_dir[58]
port 87 nsew signal output
rlabel metal3 s 494200 141448 495000 141568 6 gfpga_pad_io_soc_dir[59]
port 88 nsew signal output
rlabel metal2 s 90638 542200 90694 543000 6 gfpga_pad_io_soc_dir[5]
port 89 nsew signal output
rlabel metal3 s 494200 125536 495000 125656 6 gfpga_pad_io_soc_dir[60]
port 90 nsew signal output
rlabel metal3 s 494200 109624 495000 109744 6 gfpga_pad_io_soc_dir[61]
port 91 nsew signal output
rlabel metal3 s 494200 93712 495000 93832 6 gfpga_pad_io_soc_dir[62]
port 92 nsew signal output
rlabel metal3 s 494200 77800 495000 77920 6 gfpga_pad_io_soc_dir[63]
port 93 nsew signal output
rlabel metal3 s 494200 61888 495000 62008 6 gfpga_pad_io_soc_dir[64]
port 94 nsew signal output
rlabel metal3 s 494200 45976 495000 46096 6 gfpga_pad_io_soc_dir[65]
port 95 nsew signal output
rlabel metal3 s 494200 30064 495000 30184 6 gfpga_pad_io_soc_dir[66]
port 96 nsew signal output
rlabel metal3 s 494200 14152 495000 14272 6 gfpga_pad_io_soc_dir[67]
port 97 nsew signal output
rlabel metal2 s 479246 0 479302 800 6 gfpga_pad_io_soc_dir[68]
port 98 nsew signal output
rlabel metal2 s 461858 0 461914 800 6 gfpga_pad_io_soc_dir[69]
port 99 nsew signal output
rlabel metal2 s 103886 542200 103942 543000 6 gfpga_pad_io_soc_dir[6]
port 100 nsew signal output
rlabel metal2 s 444470 0 444526 800 6 gfpga_pad_io_soc_dir[70]
port 101 nsew signal output
rlabel metal2 s 427082 0 427138 800 6 gfpga_pad_io_soc_dir[71]
port 102 nsew signal output
rlabel metal2 s 409694 0 409750 800 6 gfpga_pad_io_soc_dir[72]
port 103 nsew signal output
rlabel metal2 s 392306 0 392362 800 6 gfpga_pad_io_soc_dir[73]
port 104 nsew signal output
rlabel metal2 s 374918 0 374974 800 6 gfpga_pad_io_soc_dir[74]
port 105 nsew signal output
rlabel metal2 s 357530 0 357586 800 6 gfpga_pad_io_soc_dir[75]
port 106 nsew signal output
rlabel metal2 s 340142 0 340198 800 6 gfpga_pad_io_soc_dir[76]
port 107 nsew signal output
rlabel metal2 s 322754 0 322810 800 6 gfpga_pad_io_soc_dir[77]
port 108 nsew signal output
rlabel metal2 s 305366 0 305422 800 6 gfpga_pad_io_soc_dir[78]
port 109 nsew signal output
rlabel metal2 s 287978 0 288034 800 6 gfpga_pad_io_soc_dir[79]
port 110 nsew signal output
rlabel metal2 s 117134 542200 117190 543000 6 gfpga_pad_io_soc_dir[7]
port 111 nsew signal output
rlabel metal2 s 270590 0 270646 800 6 gfpga_pad_io_soc_dir[80]
port 112 nsew signal output
rlabel metal2 s 253202 0 253258 800 6 gfpga_pad_io_soc_dir[81]
port 113 nsew signal output
rlabel metal2 s 235814 0 235870 800 6 gfpga_pad_io_soc_dir[82]
port 114 nsew signal output
rlabel metal2 s 218426 0 218482 800 6 gfpga_pad_io_soc_dir[83]
port 115 nsew signal output
rlabel metal2 s 201038 0 201094 800 6 gfpga_pad_io_soc_dir[84]
port 116 nsew signal output
rlabel metal2 s 183650 0 183706 800 6 gfpga_pad_io_soc_dir[85]
port 117 nsew signal output
rlabel metal2 s 166262 0 166318 800 6 gfpga_pad_io_soc_dir[86]
port 118 nsew signal output
rlabel metal2 s 148874 0 148930 800 6 gfpga_pad_io_soc_dir[87]
port 119 nsew signal output
rlabel metal2 s 131486 0 131542 800 6 gfpga_pad_io_soc_dir[88]
port 120 nsew signal output
rlabel metal2 s 114098 0 114154 800 6 gfpga_pad_io_soc_dir[89]
port 121 nsew signal output
rlabel metal2 s 130382 542200 130438 543000 6 gfpga_pad_io_soc_dir[8]
port 122 nsew signal output
rlabel metal2 s 96710 0 96766 800 6 gfpga_pad_io_soc_dir[90]
port 123 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 gfpga_pad_io_soc_dir[91]
port 124 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 gfpga_pad_io_soc_dir[92]
port 125 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 gfpga_pad_io_soc_dir[93]
port 126 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 gfpga_pad_io_soc_dir[94]
port 127 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 gfpga_pad_io_soc_dir[95]
port 128 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 gfpga_pad_io_soc_dir[96]
port 129 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 gfpga_pad_io_soc_dir[97]
port 130 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 gfpga_pad_io_soc_dir[98]
port 131 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 gfpga_pad_io_soc_dir[99]
port 132 nsew signal output
rlabel metal2 s 143630 542200 143686 543000 6 gfpga_pad_io_soc_dir[9]
port 133 nsew signal output
rlabel metal2 s 6734 542200 6790 543000 6 gfpga_pad_io_soc_in[0]
port 134 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 gfpga_pad_io_soc_in[100]
port 135 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 gfpga_pad_io_soc_in[101]
port 136 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 gfpga_pad_io_soc_in[102]
port 137 nsew signal input
rlabel metal3 s 0 129888 800 130008 6 gfpga_pad_io_soc_in[103]
port 138 nsew signal input
rlabel metal3 s 0 146208 800 146328 6 gfpga_pad_io_soc_in[104]
port 139 nsew signal input
rlabel metal3 s 0 162528 800 162648 6 gfpga_pad_io_soc_in[105]
port 140 nsew signal input
rlabel metal3 s 0 178848 800 178968 6 gfpga_pad_io_soc_in[106]
port 141 nsew signal input
rlabel metal3 s 0 195168 800 195288 6 gfpga_pad_io_soc_in[107]
port 142 nsew signal input
rlabel metal3 s 0 211488 800 211608 6 gfpga_pad_io_soc_in[108]
port 143 nsew signal input
rlabel metal3 s 0 227808 800 227928 6 gfpga_pad_io_soc_in[109]
port 144 nsew signal input
rlabel metal2 s 148046 542200 148102 543000 6 gfpga_pad_io_soc_in[10]
port 145 nsew signal input
rlabel metal3 s 0 244128 800 244248 6 gfpga_pad_io_soc_in[110]
port 146 nsew signal input
rlabel metal3 s 0 265888 800 266008 6 gfpga_pad_io_soc_in[111]
port 147 nsew signal input
rlabel metal3 s 0 282208 800 282328 6 gfpga_pad_io_soc_in[112]
port 148 nsew signal input
rlabel metal3 s 0 298528 800 298648 6 gfpga_pad_io_soc_in[113]
port 149 nsew signal input
rlabel metal3 s 0 314848 800 314968 6 gfpga_pad_io_soc_in[114]
port 150 nsew signal input
rlabel metal3 s 0 331168 800 331288 6 gfpga_pad_io_soc_in[115]
port 151 nsew signal input
rlabel metal3 s 0 347488 800 347608 6 gfpga_pad_io_soc_in[116]
port 152 nsew signal input
rlabel metal3 s 0 363808 800 363928 6 gfpga_pad_io_soc_in[117]
port 153 nsew signal input
rlabel metal3 s 0 380128 800 380248 6 gfpga_pad_io_soc_in[118]
port 154 nsew signal input
rlabel metal3 s 0 396448 800 396568 6 gfpga_pad_io_soc_in[119]
port 155 nsew signal input
rlabel metal2 s 161294 542200 161350 543000 6 gfpga_pad_io_soc_in[11]
port 156 nsew signal input
rlabel metal3 s 0 412768 800 412888 6 gfpga_pad_io_soc_in[120]
port 157 nsew signal input
rlabel metal3 s 0 429088 800 429208 6 gfpga_pad_io_soc_in[121]
port 158 nsew signal input
rlabel metal3 s 0 445408 800 445528 6 gfpga_pad_io_soc_in[122]
port 159 nsew signal input
rlabel metal3 s 0 461728 800 461848 6 gfpga_pad_io_soc_in[123]
port 160 nsew signal input
rlabel metal3 s 0 478048 800 478168 6 gfpga_pad_io_soc_in[124]
port 161 nsew signal input
rlabel metal3 s 0 494368 800 494488 6 gfpga_pad_io_soc_in[125]
port 162 nsew signal input
rlabel metal3 s 0 510688 800 510808 6 gfpga_pad_io_soc_in[126]
port 163 nsew signal input
rlabel metal3 s 0 527008 800 527128 6 gfpga_pad_io_soc_in[127]
port 164 nsew signal input
rlabel metal2 s 174542 542200 174598 543000 6 gfpga_pad_io_soc_in[12]
port 165 nsew signal input
rlabel metal2 s 187790 542200 187846 543000 6 gfpga_pad_io_soc_in[13]
port 166 nsew signal input
rlabel metal2 s 201038 542200 201094 543000 6 gfpga_pad_io_soc_in[14]
port 167 nsew signal input
rlabel metal2 s 214286 542200 214342 543000 6 gfpga_pad_io_soc_in[15]
port 168 nsew signal input
rlabel metal2 s 227534 542200 227590 543000 6 gfpga_pad_io_soc_in[16]
port 169 nsew signal input
rlabel metal2 s 240782 542200 240838 543000 6 gfpga_pad_io_soc_in[17]
port 170 nsew signal input
rlabel metal2 s 254030 542200 254086 543000 6 gfpga_pad_io_soc_in[18]
port 171 nsew signal input
rlabel metal2 s 267278 542200 267334 543000 6 gfpga_pad_io_soc_in[19]
port 172 nsew signal input
rlabel metal2 s 19982 542200 20038 543000 6 gfpga_pad_io_soc_in[1]
port 173 nsew signal input
rlabel metal2 s 280526 542200 280582 543000 6 gfpga_pad_io_soc_in[20]
port 174 nsew signal input
rlabel metal2 s 293774 542200 293830 543000 6 gfpga_pad_io_soc_in[21]
port 175 nsew signal input
rlabel metal2 s 307022 542200 307078 543000 6 gfpga_pad_io_soc_in[22]
port 176 nsew signal input
rlabel metal2 s 320270 542200 320326 543000 6 gfpga_pad_io_soc_in[23]
port 177 nsew signal input
rlabel metal2 s 333518 542200 333574 543000 6 gfpga_pad_io_soc_in[24]
port 178 nsew signal input
rlabel metal2 s 346766 542200 346822 543000 6 gfpga_pad_io_soc_in[25]
port 179 nsew signal input
rlabel metal2 s 360014 542200 360070 543000 6 gfpga_pad_io_soc_in[26]
port 180 nsew signal input
rlabel metal2 s 373262 542200 373318 543000 6 gfpga_pad_io_soc_in[27]
port 181 nsew signal input
rlabel metal2 s 386510 542200 386566 543000 6 gfpga_pad_io_soc_in[28]
port 182 nsew signal input
rlabel metal2 s 399758 542200 399814 543000 6 gfpga_pad_io_soc_in[29]
port 183 nsew signal input
rlabel metal2 s 33230 542200 33286 543000 6 gfpga_pad_io_soc_in[2]
port 184 nsew signal input
rlabel metal2 s 413006 542200 413062 543000 6 gfpga_pad_io_soc_in[30]
port 185 nsew signal input
rlabel metal2 s 426254 542200 426310 543000 6 gfpga_pad_io_soc_in[31]
port 186 nsew signal input
rlabel metal2 s 439502 542200 439558 543000 6 gfpga_pad_io_soc_in[32]
port 187 nsew signal input
rlabel metal2 s 452750 542200 452806 543000 6 gfpga_pad_io_soc_in[33]
port 188 nsew signal input
rlabel metal2 s 465998 542200 466054 543000 6 gfpga_pad_io_soc_in[34]
port 189 nsew signal input
rlabel metal2 s 479246 542200 479302 543000 6 gfpga_pad_io_soc_in[35]
port 190 nsew signal input
rlabel metal3 s 494200 528640 495000 528760 6 gfpga_pad_io_soc_in[36]
port 191 nsew signal input
rlabel metal3 s 494200 512728 495000 512848 6 gfpga_pad_io_soc_in[37]
port 192 nsew signal input
rlabel metal3 s 494200 496816 495000 496936 6 gfpga_pad_io_soc_in[38]
port 193 nsew signal input
rlabel metal3 s 494200 480904 495000 481024 6 gfpga_pad_io_soc_in[39]
port 194 nsew signal input
rlabel metal2 s 46478 542200 46534 543000 6 gfpga_pad_io_soc_in[3]
port 195 nsew signal input
rlabel metal3 s 494200 464992 495000 465112 6 gfpga_pad_io_soc_in[40]
port 196 nsew signal input
rlabel metal3 s 494200 449080 495000 449200 6 gfpga_pad_io_soc_in[41]
port 197 nsew signal input
rlabel metal3 s 494200 433168 495000 433288 6 gfpga_pad_io_soc_in[42]
port 198 nsew signal input
rlabel metal3 s 494200 417256 495000 417376 6 gfpga_pad_io_soc_in[43]
port 199 nsew signal input
rlabel metal3 s 494200 401344 495000 401464 6 gfpga_pad_io_soc_in[44]
port 200 nsew signal input
rlabel metal3 s 494200 385432 495000 385552 6 gfpga_pad_io_soc_in[45]
port 201 nsew signal input
rlabel metal3 s 494200 369520 495000 369640 6 gfpga_pad_io_soc_in[46]
port 202 nsew signal input
rlabel metal3 s 494200 353608 495000 353728 6 gfpga_pad_io_soc_in[47]
port 203 nsew signal input
rlabel metal3 s 494200 337696 495000 337816 6 gfpga_pad_io_soc_in[48]
port 204 nsew signal input
rlabel metal3 s 494200 321784 495000 321904 6 gfpga_pad_io_soc_in[49]
port 205 nsew signal input
rlabel metal2 s 68558 542200 68614 543000 6 gfpga_pad_io_soc_in[4]
port 206 nsew signal input
rlabel metal3 s 494200 305872 495000 305992 6 gfpga_pad_io_soc_in[50]
port 207 nsew signal input
rlabel metal3 s 494200 289960 495000 290080 6 gfpga_pad_io_soc_in[51]
port 208 nsew signal input
rlabel metal3 s 494200 274048 495000 274168 6 gfpga_pad_io_soc_in[52]
port 209 nsew signal input
rlabel metal3 s 494200 258136 495000 258256 6 gfpga_pad_io_soc_in[53]
port 210 nsew signal input
rlabel metal3 s 494200 231616 495000 231736 6 gfpga_pad_io_soc_in[54]
port 211 nsew signal input
rlabel metal3 s 494200 215704 495000 215824 6 gfpga_pad_io_soc_in[55]
port 212 nsew signal input
rlabel metal3 s 494200 199792 495000 199912 6 gfpga_pad_io_soc_in[56]
port 213 nsew signal input
rlabel metal3 s 494200 183880 495000 184000 6 gfpga_pad_io_soc_in[57]
port 214 nsew signal input
rlabel metal3 s 494200 167968 495000 168088 6 gfpga_pad_io_soc_in[58]
port 215 nsew signal input
rlabel metal3 s 494200 152056 495000 152176 6 gfpga_pad_io_soc_in[59]
port 216 nsew signal input
rlabel metal2 s 81806 542200 81862 543000 6 gfpga_pad_io_soc_in[5]
port 217 nsew signal input
rlabel metal3 s 494200 136144 495000 136264 6 gfpga_pad_io_soc_in[60]
port 218 nsew signal input
rlabel metal3 s 494200 120232 495000 120352 6 gfpga_pad_io_soc_in[61]
port 219 nsew signal input
rlabel metal3 s 494200 104320 495000 104440 6 gfpga_pad_io_soc_in[62]
port 220 nsew signal input
rlabel metal3 s 494200 88408 495000 88528 6 gfpga_pad_io_soc_in[63]
port 221 nsew signal input
rlabel metal3 s 494200 72496 495000 72616 6 gfpga_pad_io_soc_in[64]
port 222 nsew signal input
rlabel metal3 s 494200 56584 495000 56704 6 gfpga_pad_io_soc_in[65]
port 223 nsew signal input
rlabel metal3 s 494200 40672 495000 40792 6 gfpga_pad_io_soc_in[66]
port 224 nsew signal input
rlabel metal3 s 494200 24760 495000 24880 6 gfpga_pad_io_soc_in[67]
port 225 nsew signal input
rlabel metal2 s 490838 0 490894 800 6 gfpga_pad_io_soc_in[68]
port 226 nsew signal input
rlabel metal2 s 473450 0 473506 800 6 gfpga_pad_io_soc_in[69]
port 227 nsew signal input
rlabel metal2 s 95054 542200 95110 543000 6 gfpga_pad_io_soc_in[6]
port 228 nsew signal input
rlabel metal2 s 456062 0 456118 800 6 gfpga_pad_io_soc_in[70]
port 229 nsew signal input
rlabel metal2 s 438674 0 438730 800 6 gfpga_pad_io_soc_in[71]
port 230 nsew signal input
rlabel metal2 s 421286 0 421342 800 6 gfpga_pad_io_soc_in[72]
port 231 nsew signal input
rlabel metal2 s 403898 0 403954 800 6 gfpga_pad_io_soc_in[73]
port 232 nsew signal input
rlabel metal2 s 386510 0 386566 800 6 gfpga_pad_io_soc_in[74]
port 233 nsew signal input
rlabel metal2 s 369122 0 369178 800 6 gfpga_pad_io_soc_in[75]
port 234 nsew signal input
rlabel metal2 s 351734 0 351790 800 6 gfpga_pad_io_soc_in[76]
port 235 nsew signal input
rlabel metal2 s 334346 0 334402 800 6 gfpga_pad_io_soc_in[77]
port 236 nsew signal input
rlabel metal2 s 316958 0 317014 800 6 gfpga_pad_io_soc_in[78]
port 237 nsew signal input
rlabel metal2 s 299570 0 299626 800 6 gfpga_pad_io_soc_in[79]
port 238 nsew signal input
rlabel metal2 s 108302 542200 108358 543000 6 gfpga_pad_io_soc_in[7]
port 239 nsew signal input
rlabel metal2 s 282182 0 282238 800 6 gfpga_pad_io_soc_in[80]
port 240 nsew signal input
rlabel metal2 s 264794 0 264850 800 6 gfpga_pad_io_soc_in[81]
port 241 nsew signal input
rlabel metal2 s 247406 0 247462 800 6 gfpga_pad_io_soc_in[82]
port 242 nsew signal input
rlabel metal2 s 230018 0 230074 800 6 gfpga_pad_io_soc_in[83]
port 243 nsew signal input
rlabel metal2 s 212630 0 212686 800 6 gfpga_pad_io_soc_in[84]
port 244 nsew signal input
rlabel metal2 s 195242 0 195298 800 6 gfpga_pad_io_soc_in[85]
port 245 nsew signal input
rlabel metal2 s 177854 0 177910 800 6 gfpga_pad_io_soc_in[86]
port 246 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 gfpga_pad_io_soc_in[87]
port 247 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 gfpga_pad_io_soc_in[88]
port 248 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 gfpga_pad_io_soc_in[89]
port 249 nsew signal input
rlabel metal2 s 121550 542200 121606 543000 6 gfpga_pad_io_soc_in[8]
port 250 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 gfpga_pad_io_soc_in[90]
port 251 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 gfpga_pad_io_soc_in[91]
port 252 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 gfpga_pad_io_soc_in[92]
port 253 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 gfpga_pad_io_soc_in[93]
port 254 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 gfpga_pad_io_soc_in[94]
port 255 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 gfpga_pad_io_soc_in[95]
port 256 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 gfpga_pad_io_soc_in[96]
port 257 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 gfpga_pad_io_soc_in[97]
port 258 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 gfpga_pad_io_soc_in[98]
port 259 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 gfpga_pad_io_soc_in[99]
port 260 nsew signal input
rlabel metal2 s 134798 542200 134854 543000 6 gfpga_pad_io_soc_in[9]
port 261 nsew signal input
rlabel metal2 s 11150 542200 11206 543000 6 gfpga_pad_io_soc_out[0]
port 262 nsew signal output
rlabel metal3 s 0 86368 800 86488 6 gfpga_pad_io_soc_out[100]
port 263 nsew signal output
rlabel metal3 s 0 102688 800 102808 6 gfpga_pad_io_soc_out[101]
port 264 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 gfpga_pad_io_soc_out[102]
port 265 nsew signal output
rlabel metal3 s 0 135328 800 135448 6 gfpga_pad_io_soc_out[103]
port 266 nsew signal output
rlabel metal3 s 0 151648 800 151768 6 gfpga_pad_io_soc_out[104]
port 267 nsew signal output
rlabel metal3 s 0 167968 800 168088 6 gfpga_pad_io_soc_out[105]
port 268 nsew signal output
rlabel metal3 s 0 184288 800 184408 6 gfpga_pad_io_soc_out[106]
port 269 nsew signal output
rlabel metal3 s 0 200608 800 200728 6 gfpga_pad_io_soc_out[107]
port 270 nsew signal output
rlabel metal3 s 0 216928 800 217048 6 gfpga_pad_io_soc_out[108]
port 271 nsew signal output
rlabel metal3 s 0 233248 800 233368 6 gfpga_pad_io_soc_out[109]
port 272 nsew signal output
rlabel metal2 s 152462 542200 152518 543000 6 gfpga_pad_io_soc_out[10]
port 273 nsew signal output
rlabel metal3 s 0 249568 800 249688 6 gfpga_pad_io_soc_out[110]
port 274 nsew signal output
rlabel metal3 s 0 271328 800 271448 6 gfpga_pad_io_soc_out[111]
port 275 nsew signal output
rlabel metal3 s 0 287648 800 287768 6 gfpga_pad_io_soc_out[112]
port 276 nsew signal output
rlabel metal3 s 0 303968 800 304088 6 gfpga_pad_io_soc_out[113]
port 277 nsew signal output
rlabel metal3 s 0 320288 800 320408 6 gfpga_pad_io_soc_out[114]
port 278 nsew signal output
rlabel metal3 s 0 336608 800 336728 6 gfpga_pad_io_soc_out[115]
port 279 nsew signal output
rlabel metal3 s 0 352928 800 353048 6 gfpga_pad_io_soc_out[116]
port 280 nsew signal output
rlabel metal3 s 0 369248 800 369368 6 gfpga_pad_io_soc_out[117]
port 281 nsew signal output
rlabel metal3 s 0 385568 800 385688 6 gfpga_pad_io_soc_out[118]
port 282 nsew signal output
rlabel metal3 s 0 401888 800 402008 6 gfpga_pad_io_soc_out[119]
port 283 nsew signal output
rlabel metal2 s 165710 542200 165766 543000 6 gfpga_pad_io_soc_out[11]
port 284 nsew signal output
rlabel metal3 s 0 418208 800 418328 6 gfpga_pad_io_soc_out[120]
port 285 nsew signal output
rlabel metal3 s 0 434528 800 434648 6 gfpga_pad_io_soc_out[121]
port 286 nsew signal output
rlabel metal3 s 0 450848 800 450968 6 gfpga_pad_io_soc_out[122]
port 287 nsew signal output
rlabel metal3 s 0 467168 800 467288 6 gfpga_pad_io_soc_out[123]
port 288 nsew signal output
rlabel metal3 s 0 483488 800 483608 6 gfpga_pad_io_soc_out[124]
port 289 nsew signal output
rlabel metal3 s 0 499808 800 499928 6 gfpga_pad_io_soc_out[125]
port 290 nsew signal output
rlabel metal3 s 0 516128 800 516248 6 gfpga_pad_io_soc_out[126]
port 291 nsew signal output
rlabel metal3 s 0 532448 800 532568 6 gfpga_pad_io_soc_out[127]
port 292 nsew signal output
rlabel metal2 s 178958 542200 179014 543000 6 gfpga_pad_io_soc_out[12]
port 293 nsew signal output
rlabel metal2 s 192206 542200 192262 543000 6 gfpga_pad_io_soc_out[13]
port 294 nsew signal output
rlabel metal2 s 205454 542200 205510 543000 6 gfpga_pad_io_soc_out[14]
port 295 nsew signal output
rlabel metal2 s 218702 542200 218758 543000 6 gfpga_pad_io_soc_out[15]
port 296 nsew signal output
rlabel metal2 s 231950 542200 232006 543000 6 gfpga_pad_io_soc_out[16]
port 297 nsew signal output
rlabel metal2 s 245198 542200 245254 543000 6 gfpga_pad_io_soc_out[17]
port 298 nsew signal output
rlabel metal2 s 258446 542200 258502 543000 6 gfpga_pad_io_soc_out[18]
port 299 nsew signal output
rlabel metal2 s 271694 542200 271750 543000 6 gfpga_pad_io_soc_out[19]
port 300 nsew signal output
rlabel metal2 s 24398 542200 24454 543000 6 gfpga_pad_io_soc_out[1]
port 301 nsew signal output
rlabel metal2 s 284942 542200 284998 543000 6 gfpga_pad_io_soc_out[20]
port 302 nsew signal output
rlabel metal2 s 298190 542200 298246 543000 6 gfpga_pad_io_soc_out[21]
port 303 nsew signal output
rlabel metal2 s 311438 542200 311494 543000 6 gfpga_pad_io_soc_out[22]
port 304 nsew signal output
rlabel metal2 s 324686 542200 324742 543000 6 gfpga_pad_io_soc_out[23]
port 305 nsew signal output
rlabel metal2 s 337934 542200 337990 543000 6 gfpga_pad_io_soc_out[24]
port 306 nsew signal output
rlabel metal2 s 351182 542200 351238 543000 6 gfpga_pad_io_soc_out[25]
port 307 nsew signal output
rlabel metal2 s 364430 542200 364486 543000 6 gfpga_pad_io_soc_out[26]
port 308 nsew signal output
rlabel metal2 s 377678 542200 377734 543000 6 gfpga_pad_io_soc_out[27]
port 309 nsew signal output
rlabel metal2 s 390926 542200 390982 543000 6 gfpga_pad_io_soc_out[28]
port 310 nsew signal output
rlabel metal2 s 404174 542200 404230 543000 6 gfpga_pad_io_soc_out[29]
port 311 nsew signal output
rlabel metal2 s 37646 542200 37702 543000 6 gfpga_pad_io_soc_out[2]
port 312 nsew signal output
rlabel metal2 s 417422 542200 417478 543000 6 gfpga_pad_io_soc_out[30]
port 313 nsew signal output
rlabel metal2 s 430670 542200 430726 543000 6 gfpga_pad_io_soc_out[31]
port 314 nsew signal output
rlabel metal2 s 443918 542200 443974 543000 6 gfpga_pad_io_soc_out[32]
port 315 nsew signal output
rlabel metal2 s 457166 542200 457222 543000 6 gfpga_pad_io_soc_out[33]
port 316 nsew signal output
rlabel metal2 s 470414 542200 470470 543000 6 gfpga_pad_io_soc_out[34]
port 317 nsew signal output
rlabel metal2 s 483662 542200 483718 543000 6 gfpga_pad_io_soc_out[35]
port 318 nsew signal output
rlabel metal3 s 494200 523336 495000 523456 6 gfpga_pad_io_soc_out[36]
port 319 nsew signal output
rlabel metal3 s 494200 507424 495000 507544 6 gfpga_pad_io_soc_out[37]
port 320 nsew signal output
rlabel metal3 s 494200 491512 495000 491632 6 gfpga_pad_io_soc_out[38]
port 321 nsew signal output
rlabel metal3 s 494200 475600 495000 475720 6 gfpga_pad_io_soc_out[39]
port 322 nsew signal output
rlabel metal2 s 50894 542200 50950 543000 6 gfpga_pad_io_soc_out[3]
port 323 nsew signal output
rlabel metal3 s 494200 459688 495000 459808 6 gfpga_pad_io_soc_out[40]
port 324 nsew signal output
rlabel metal3 s 494200 443776 495000 443896 6 gfpga_pad_io_soc_out[41]
port 325 nsew signal output
rlabel metal3 s 494200 427864 495000 427984 6 gfpga_pad_io_soc_out[42]
port 326 nsew signal output
rlabel metal3 s 494200 411952 495000 412072 6 gfpga_pad_io_soc_out[43]
port 327 nsew signal output
rlabel metal3 s 494200 396040 495000 396160 6 gfpga_pad_io_soc_out[44]
port 328 nsew signal output
rlabel metal3 s 494200 380128 495000 380248 6 gfpga_pad_io_soc_out[45]
port 329 nsew signal output
rlabel metal3 s 494200 364216 495000 364336 6 gfpga_pad_io_soc_out[46]
port 330 nsew signal output
rlabel metal3 s 494200 348304 495000 348424 6 gfpga_pad_io_soc_out[47]
port 331 nsew signal output
rlabel metal3 s 494200 332392 495000 332512 6 gfpga_pad_io_soc_out[48]
port 332 nsew signal output
rlabel metal3 s 494200 316480 495000 316600 6 gfpga_pad_io_soc_out[49]
port 333 nsew signal output
rlabel metal2 s 72974 542200 73030 543000 6 gfpga_pad_io_soc_out[4]
port 334 nsew signal output
rlabel metal3 s 494200 300568 495000 300688 6 gfpga_pad_io_soc_out[50]
port 335 nsew signal output
rlabel metal3 s 494200 284656 495000 284776 6 gfpga_pad_io_soc_out[51]
port 336 nsew signal output
rlabel metal3 s 494200 268744 495000 268864 6 gfpga_pad_io_soc_out[52]
port 337 nsew signal output
rlabel metal3 s 494200 252832 495000 252952 6 gfpga_pad_io_soc_out[53]
port 338 nsew signal output
rlabel metal3 s 494200 226312 495000 226432 6 gfpga_pad_io_soc_out[54]
port 339 nsew signal output
rlabel metal3 s 494200 210400 495000 210520 6 gfpga_pad_io_soc_out[55]
port 340 nsew signal output
rlabel metal3 s 494200 194488 495000 194608 6 gfpga_pad_io_soc_out[56]
port 341 nsew signal output
rlabel metal3 s 494200 178576 495000 178696 6 gfpga_pad_io_soc_out[57]
port 342 nsew signal output
rlabel metal3 s 494200 162664 495000 162784 6 gfpga_pad_io_soc_out[58]
port 343 nsew signal output
rlabel metal3 s 494200 146752 495000 146872 6 gfpga_pad_io_soc_out[59]
port 344 nsew signal output
rlabel metal2 s 86222 542200 86278 543000 6 gfpga_pad_io_soc_out[5]
port 345 nsew signal output
rlabel metal3 s 494200 130840 495000 130960 6 gfpga_pad_io_soc_out[60]
port 346 nsew signal output
rlabel metal3 s 494200 114928 495000 115048 6 gfpga_pad_io_soc_out[61]
port 347 nsew signal output
rlabel metal3 s 494200 99016 495000 99136 6 gfpga_pad_io_soc_out[62]
port 348 nsew signal output
rlabel metal3 s 494200 83104 495000 83224 6 gfpga_pad_io_soc_out[63]
port 349 nsew signal output
rlabel metal3 s 494200 67192 495000 67312 6 gfpga_pad_io_soc_out[64]
port 350 nsew signal output
rlabel metal3 s 494200 51280 495000 51400 6 gfpga_pad_io_soc_out[65]
port 351 nsew signal output
rlabel metal3 s 494200 35368 495000 35488 6 gfpga_pad_io_soc_out[66]
port 352 nsew signal output
rlabel metal3 s 494200 19456 495000 19576 6 gfpga_pad_io_soc_out[67]
port 353 nsew signal output
rlabel metal2 s 485042 0 485098 800 6 gfpga_pad_io_soc_out[68]
port 354 nsew signal output
rlabel metal2 s 467654 0 467710 800 6 gfpga_pad_io_soc_out[69]
port 355 nsew signal output
rlabel metal2 s 99470 542200 99526 543000 6 gfpga_pad_io_soc_out[6]
port 356 nsew signal output
rlabel metal2 s 450266 0 450322 800 6 gfpga_pad_io_soc_out[70]
port 357 nsew signal output
rlabel metal2 s 432878 0 432934 800 6 gfpga_pad_io_soc_out[71]
port 358 nsew signal output
rlabel metal2 s 415490 0 415546 800 6 gfpga_pad_io_soc_out[72]
port 359 nsew signal output
rlabel metal2 s 398102 0 398158 800 6 gfpga_pad_io_soc_out[73]
port 360 nsew signal output
rlabel metal2 s 380714 0 380770 800 6 gfpga_pad_io_soc_out[74]
port 361 nsew signal output
rlabel metal2 s 363326 0 363382 800 6 gfpga_pad_io_soc_out[75]
port 362 nsew signal output
rlabel metal2 s 345938 0 345994 800 6 gfpga_pad_io_soc_out[76]
port 363 nsew signal output
rlabel metal2 s 328550 0 328606 800 6 gfpga_pad_io_soc_out[77]
port 364 nsew signal output
rlabel metal2 s 311162 0 311218 800 6 gfpga_pad_io_soc_out[78]
port 365 nsew signal output
rlabel metal2 s 293774 0 293830 800 6 gfpga_pad_io_soc_out[79]
port 366 nsew signal output
rlabel metal2 s 112718 542200 112774 543000 6 gfpga_pad_io_soc_out[7]
port 367 nsew signal output
rlabel metal2 s 276386 0 276442 800 6 gfpga_pad_io_soc_out[80]
port 368 nsew signal output
rlabel metal2 s 258998 0 259054 800 6 gfpga_pad_io_soc_out[81]
port 369 nsew signal output
rlabel metal2 s 241610 0 241666 800 6 gfpga_pad_io_soc_out[82]
port 370 nsew signal output
rlabel metal2 s 224222 0 224278 800 6 gfpga_pad_io_soc_out[83]
port 371 nsew signal output
rlabel metal2 s 206834 0 206890 800 6 gfpga_pad_io_soc_out[84]
port 372 nsew signal output
rlabel metal2 s 189446 0 189502 800 6 gfpga_pad_io_soc_out[85]
port 373 nsew signal output
rlabel metal2 s 172058 0 172114 800 6 gfpga_pad_io_soc_out[86]
port 374 nsew signal output
rlabel metal2 s 154670 0 154726 800 6 gfpga_pad_io_soc_out[87]
port 375 nsew signal output
rlabel metal2 s 137282 0 137338 800 6 gfpga_pad_io_soc_out[88]
port 376 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 gfpga_pad_io_soc_out[89]
port 377 nsew signal output
rlabel metal2 s 125966 542200 126022 543000 6 gfpga_pad_io_soc_out[8]
port 378 nsew signal output
rlabel metal2 s 102506 0 102562 800 6 gfpga_pad_io_soc_out[90]
port 379 nsew signal output
rlabel metal2 s 85118 0 85174 800 6 gfpga_pad_io_soc_out[91]
port 380 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 gfpga_pad_io_soc_out[92]
port 381 nsew signal output
rlabel metal2 s 44546 0 44602 800 6 gfpga_pad_io_soc_out[93]
port 382 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 gfpga_pad_io_soc_out[94]
port 383 nsew signal output
rlabel metal2 s 9770 0 9826 800 6 gfpga_pad_io_soc_out[95]
port 384 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 gfpga_pad_io_soc_out[96]
port 385 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 gfpga_pad_io_soc_out[97]
port 386 nsew signal output
rlabel metal3 s 0 53728 800 53848 6 gfpga_pad_io_soc_out[98]
port 387 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 gfpga_pad_io_soc_out[99]
port 388 nsew signal output
rlabel metal2 s 139214 542200 139270 543000 6 gfpga_pad_io_soc_out[9]
port 389 nsew signal output
rlabel metal3 s 494200 8848 495000 8968 6 isol_n
port 390 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 prog_clk
port 391 nsew signal input
rlabel metal3 s 0 260448 800 260568 6 prog_reset
port 392 nsew signal input
rlabel metal3 s 494200 236920 495000 237040 6 reset
port 393 nsew signal input
rlabel metal2 s 64142 542200 64198 543000 6 sc_head
port 394 nsew signal input
rlabel metal3 s 494200 533944 495000 534064 6 sc_tail
port 395 nsew signal output
rlabel metal3 s 494200 242224 495000 242344 6 test_enable
port 396 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 495000 543000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 79861408
string GDS_FILE /home/hosni/OpenFPGA/erc-fixes/clear/openlane/fpga_core/runs/23_04_16_15_53/results/signoff/fpga_core.magic.gds
string GDS_START 44272806
<< end >>

