//Generated from netlist by SpyDrNet
//netlist name: FPGA88_SOFA_A
module const1
(
    const1
);

    output const1;

    wire \<const1> = 1 ;
    wire const1;

assign const1 = \<const1> ;
endmodule

