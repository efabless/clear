magic
tech sky130A
magscale 1 2
timestamp 1679346777
<< obsli1 >>
rect 1104 2159 25852 54417
<< obsm1 >>
rect 934 2128 26114 54448
<< metal2 >>
rect 938 56200 994 57000
rect 1306 56200 1362 57000
rect 1674 56200 1730 57000
rect 2042 56200 2098 57000
rect 2410 56200 2466 57000
rect 2778 56200 2834 57000
rect 3146 56200 3202 57000
rect 3514 56200 3570 57000
rect 3882 56200 3938 57000
rect 4250 56200 4306 57000
rect 4618 56200 4674 57000
rect 4986 56200 5042 57000
rect 5354 56200 5410 57000
rect 5722 56200 5778 57000
rect 6090 56200 6146 57000
rect 6458 56200 6514 57000
rect 6826 56200 6882 57000
rect 7194 56200 7250 57000
rect 7562 56200 7618 57000
rect 7930 56200 7986 57000
rect 8298 56200 8354 57000
rect 8666 56200 8722 57000
rect 9034 56200 9090 57000
rect 9402 56200 9458 57000
rect 9770 56200 9826 57000
rect 10138 56200 10194 57000
rect 10506 56200 10562 57000
rect 10874 56200 10930 57000
rect 11242 56200 11298 57000
rect 11610 56200 11666 57000
rect 11978 56200 12034 57000
rect 12346 56200 12402 57000
rect 12714 56200 12770 57000
rect 13082 56200 13138 57000
rect 13450 56200 13506 57000
rect 13818 56200 13874 57000
rect 14186 56200 14242 57000
rect 14554 56200 14610 57000
rect 14922 56200 14978 57000
rect 15290 56200 15346 57000
rect 15658 56200 15714 57000
rect 16026 56200 16082 57000
rect 16394 56200 16450 57000
rect 16762 56200 16818 57000
rect 17130 56200 17186 57000
rect 17498 56200 17554 57000
rect 17866 56200 17922 57000
rect 18234 56200 18290 57000
rect 18602 56200 18658 57000
rect 18970 56200 19026 57000
rect 19338 56200 19394 57000
rect 19706 56200 19762 57000
rect 20074 56200 20130 57000
rect 20442 56200 20498 57000
rect 20810 56200 20866 57000
rect 21178 56200 21234 57000
rect 21546 56200 21602 57000
rect 21914 56200 21970 57000
rect 22282 56200 22338 57000
rect 22650 56200 22706 57000
rect 23018 56200 23074 57000
rect 24122 56200 24178 57000
rect 24490 56200 24546 57000
rect 24858 56200 24914 57000
rect 25226 56200 25282 57000
rect 25594 56200 25650 57000
rect 25962 56200 26018 57000
rect 1122 0 1178 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21730 0 21786 800
rect 22098 0 22154 800
rect 22466 0 22522 800
rect 22834 0 22890 800
rect 23202 0 23258 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 25042 0 25098 800
rect 25410 0 25466 800
<< obsm2 >>
rect 1050 56144 1250 56250
rect 1418 56144 1618 56250
rect 1786 56144 1986 56250
rect 2154 56144 2354 56250
rect 2522 56144 2722 56250
rect 2890 56144 3090 56250
rect 3258 56144 3458 56250
rect 3626 56144 3826 56250
rect 3994 56144 4194 56250
rect 4362 56144 4562 56250
rect 4730 56144 4930 56250
rect 5098 56144 5298 56250
rect 5466 56144 5666 56250
rect 5834 56144 6034 56250
rect 6202 56144 6402 56250
rect 6570 56144 6770 56250
rect 6938 56144 7138 56250
rect 7306 56144 7506 56250
rect 7674 56144 7874 56250
rect 8042 56144 8242 56250
rect 8410 56144 8610 56250
rect 8778 56144 8978 56250
rect 9146 56144 9346 56250
rect 9514 56144 9714 56250
rect 9882 56144 10082 56250
rect 10250 56144 10450 56250
rect 10618 56144 10818 56250
rect 10986 56144 11186 56250
rect 11354 56144 11554 56250
rect 11722 56144 11922 56250
rect 12090 56144 12290 56250
rect 12458 56144 12658 56250
rect 12826 56144 13026 56250
rect 13194 56144 13394 56250
rect 13562 56144 13762 56250
rect 13930 56144 14130 56250
rect 14298 56144 14498 56250
rect 14666 56144 14866 56250
rect 15034 56144 15234 56250
rect 15402 56144 15602 56250
rect 15770 56144 15970 56250
rect 16138 56144 16338 56250
rect 16506 56144 16706 56250
rect 16874 56144 17074 56250
rect 17242 56144 17442 56250
rect 17610 56144 17810 56250
rect 17978 56144 18178 56250
rect 18346 56144 18546 56250
rect 18714 56144 18914 56250
rect 19082 56144 19282 56250
rect 19450 56144 19650 56250
rect 19818 56144 20018 56250
rect 20186 56144 20386 56250
rect 20554 56144 20754 56250
rect 20922 56144 21122 56250
rect 21290 56144 21490 56250
rect 21658 56144 21858 56250
rect 22026 56144 22226 56250
rect 22394 56144 22594 56250
rect 22762 56144 22962 56250
rect 23130 56144 24066 56250
rect 24234 56144 24434 56250
rect 24602 56144 24802 56250
rect 24970 56144 25170 56250
rect 25338 56144 25538 56250
rect 25706 56144 25906 56250
rect 26074 56144 26110 56250
rect 938 856 26110 56144
rect 938 734 1066 856
rect 1234 734 1434 856
rect 1602 734 1802 856
rect 1970 734 2170 856
rect 2338 734 2538 856
rect 2706 734 2906 856
rect 3074 734 3274 856
rect 3442 734 3642 856
rect 3810 734 4010 856
rect 4178 734 4378 856
rect 4546 734 4746 856
rect 4914 734 5114 856
rect 5282 734 5482 856
rect 5650 734 5850 856
rect 6018 734 6218 856
rect 6386 734 6586 856
rect 6754 734 6954 856
rect 7122 734 7322 856
rect 7490 734 7690 856
rect 7858 734 8058 856
rect 8226 734 8426 856
rect 8594 734 8794 856
rect 8962 734 9162 856
rect 9330 734 9530 856
rect 9698 734 9898 856
rect 10066 734 10266 856
rect 10434 734 10634 856
rect 10802 734 11002 856
rect 11170 734 11370 856
rect 11538 734 11738 856
rect 11906 734 12106 856
rect 12274 734 12474 856
rect 12642 734 12842 856
rect 13010 734 13210 856
rect 13378 734 13578 856
rect 13746 734 13946 856
rect 14114 734 14314 856
rect 14482 734 14682 856
rect 14850 734 15050 856
rect 15218 734 15418 856
rect 15586 734 15786 856
rect 15954 734 16154 856
rect 16322 734 16522 856
rect 16690 734 16890 856
rect 17058 734 17258 856
rect 17426 734 17626 856
rect 17794 734 17994 856
rect 18162 734 18362 856
rect 18530 734 18730 856
rect 18898 734 19098 856
rect 19266 734 19466 856
rect 19634 734 19834 856
rect 20002 734 20202 856
rect 20370 734 20570 856
rect 20738 734 20938 856
rect 21106 734 21306 856
rect 21474 734 21674 856
rect 21842 734 22042 856
rect 22210 734 22410 856
rect 22578 734 22778 856
rect 22946 734 23146 856
rect 23314 734 23514 856
rect 23682 734 23882 856
rect 24050 734 24250 856
rect 24418 734 24618 856
rect 24786 734 24986 856
rect 25154 734 25354 856
rect 25522 734 26110 856
<< metal3 >>
rect 0 54952 800 55072
rect 0 52640 800 52760
rect 26200 52504 27000 52624
rect 26200 51824 27000 51944
rect 26200 51144 27000 51264
rect 0 50328 800 50448
rect 26200 50464 27000 50584
rect 26200 49784 27000 49904
rect 26200 49104 27000 49224
rect 26200 48424 27000 48544
rect 0 48016 800 48136
rect 26200 47744 27000 47864
rect 26200 47064 27000 47184
rect 26200 46384 27000 46504
rect 0 45704 800 45824
rect 26200 45704 27000 45824
rect 26200 45024 27000 45144
rect 26200 44344 27000 44464
rect 26200 43664 27000 43784
rect 0 43392 800 43512
rect 26200 42984 27000 43104
rect 26200 42304 27000 42424
rect 26200 41624 27000 41744
rect 0 41080 800 41200
rect 26200 40944 27000 41064
rect 26200 40264 27000 40384
rect 26200 39584 27000 39704
rect 0 38768 800 38888
rect 26200 38904 27000 39024
rect 26200 38224 27000 38344
rect 26200 37544 27000 37664
rect 26200 36864 27000 36984
rect 0 36456 800 36576
rect 26200 36184 27000 36304
rect 26200 35504 27000 35624
rect 26200 34824 27000 34944
rect 0 34144 800 34264
rect 26200 34144 27000 34264
rect 26200 33464 27000 33584
rect 26200 32784 27000 32904
rect 26200 32104 27000 32224
rect 0 31832 800 31952
rect 26200 31424 27000 31544
rect 26200 30744 27000 30864
rect 26200 30064 27000 30184
rect 0 29520 800 29640
rect 26200 29384 27000 29504
rect 26200 28704 27000 28824
rect 26200 28024 27000 28144
rect 0 27208 800 27328
rect 26200 27344 27000 27464
rect 26200 26664 27000 26784
rect 26200 25984 27000 26104
rect 26200 25304 27000 25424
rect 0 24896 800 25016
rect 26200 24624 27000 24744
rect 26200 23944 27000 24064
rect 26200 23264 27000 23384
rect 0 22584 800 22704
rect 26200 22584 27000 22704
rect 26200 21904 27000 22024
rect 26200 21224 27000 21344
rect 26200 20544 27000 20664
rect 0 20272 800 20392
rect 26200 19864 27000 19984
rect 26200 19184 27000 19304
rect 26200 18504 27000 18624
rect 0 17960 800 18080
rect 26200 17824 27000 17944
rect 26200 17144 27000 17264
rect 26200 16464 27000 16584
rect 0 15648 800 15768
rect 26200 15784 27000 15904
rect 26200 15104 27000 15224
rect 26200 14424 27000 14544
rect 26200 13744 27000 13864
rect 0 13336 800 13456
rect 26200 13064 27000 13184
rect 26200 12384 27000 12504
rect 26200 11704 27000 11824
rect 0 11024 800 11144
rect 26200 11024 27000 11144
rect 26200 10344 27000 10464
rect 26200 9664 27000 9784
rect 26200 8984 27000 9104
rect 0 8712 800 8832
rect 26200 8304 27000 8424
rect 26200 7624 27000 7744
rect 26200 6944 27000 7064
rect 0 6400 800 6520
rect 26200 6264 27000 6384
rect 26200 5584 27000 5704
rect 26200 4904 27000 5024
rect 0 4088 800 4208
rect 26200 4224 27000 4344
rect 0 1776 800 1896
<< obsm3 >>
rect 880 54872 26200 55045
rect 800 52840 26200 54872
rect 880 52704 26200 52840
rect 880 52560 26120 52704
rect 800 52424 26120 52560
rect 800 52024 26200 52424
rect 800 51744 26120 52024
rect 800 51344 26200 51744
rect 800 51064 26120 51344
rect 800 50664 26200 51064
rect 800 50528 26120 50664
rect 880 50384 26120 50528
rect 880 50248 26200 50384
rect 800 49984 26200 50248
rect 800 49704 26120 49984
rect 800 49304 26200 49704
rect 800 49024 26120 49304
rect 800 48624 26200 49024
rect 800 48344 26120 48624
rect 800 48216 26200 48344
rect 880 47944 26200 48216
rect 880 47936 26120 47944
rect 800 47664 26120 47936
rect 800 47264 26200 47664
rect 800 46984 26120 47264
rect 800 46584 26200 46984
rect 800 46304 26120 46584
rect 800 45904 26200 46304
rect 880 45624 26120 45904
rect 800 45224 26200 45624
rect 800 44944 26120 45224
rect 800 44544 26200 44944
rect 800 44264 26120 44544
rect 800 43864 26200 44264
rect 800 43592 26120 43864
rect 880 43584 26120 43592
rect 880 43312 26200 43584
rect 800 43184 26200 43312
rect 800 42904 26120 43184
rect 800 42504 26200 42904
rect 800 42224 26120 42504
rect 800 41824 26200 42224
rect 800 41544 26120 41824
rect 800 41280 26200 41544
rect 880 41144 26200 41280
rect 880 41000 26120 41144
rect 800 40864 26120 41000
rect 800 40464 26200 40864
rect 800 40184 26120 40464
rect 800 39784 26200 40184
rect 800 39504 26120 39784
rect 800 39104 26200 39504
rect 800 38968 26120 39104
rect 880 38824 26120 38968
rect 880 38688 26200 38824
rect 800 38424 26200 38688
rect 800 38144 26120 38424
rect 800 37744 26200 38144
rect 800 37464 26120 37744
rect 800 37064 26200 37464
rect 800 36784 26120 37064
rect 800 36656 26200 36784
rect 880 36384 26200 36656
rect 880 36376 26120 36384
rect 800 36104 26120 36376
rect 800 35704 26200 36104
rect 800 35424 26120 35704
rect 800 35024 26200 35424
rect 800 34744 26120 35024
rect 800 34344 26200 34744
rect 880 34064 26120 34344
rect 800 33664 26200 34064
rect 800 33384 26120 33664
rect 800 32984 26200 33384
rect 800 32704 26120 32984
rect 800 32304 26200 32704
rect 800 32032 26120 32304
rect 880 32024 26120 32032
rect 880 31752 26200 32024
rect 800 31624 26200 31752
rect 800 31344 26120 31624
rect 800 30944 26200 31344
rect 800 30664 26120 30944
rect 800 30264 26200 30664
rect 800 29984 26120 30264
rect 800 29720 26200 29984
rect 880 29584 26200 29720
rect 880 29440 26120 29584
rect 800 29304 26120 29440
rect 800 28904 26200 29304
rect 800 28624 26120 28904
rect 800 28224 26200 28624
rect 800 27944 26120 28224
rect 800 27544 26200 27944
rect 800 27408 26120 27544
rect 880 27264 26120 27408
rect 880 27128 26200 27264
rect 800 26864 26200 27128
rect 800 26584 26120 26864
rect 800 26184 26200 26584
rect 800 25904 26120 26184
rect 800 25504 26200 25904
rect 800 25224 26120 25504
rect 800 25096 26200 25224
rect 880 24824 26200 25096
rect 880 24816 26120 24824
rect 800 24544 26120 24816
rect 800 24144 26200 24544
rect 800 23864 26120 24144
rect 800 23464 26200 23864
rect 800 23184 26120 23464
rect 800 22784 26200 23184
rect 880 22504 26120 22784
rect 800 22104 26200 22504
rect 800 21824 26120 22104
rect 800 21424 26200 21824
rect 800 21144 26120 21424
rect 800 20744 26200 21144
rect 800 20472 26120 20744
rect 880 20464 26120 20472
rect 880 20192 26200 20464
rect 800 20064 26200 20192
rect 800 19784 26120 20064
rect 800 19384 26200 19784
rect 800 19104 26120 19384
rect 800 18704 26200 19104
rect 800 18424 26120 18704
rect 800 18160 26200 18424
rect 880 18024 26200 18160
rect 880 17880 26120 18024
rect 800 17744 26120 17880
rect 800 17344 26200 17744
rect 800 17064 26120 17344
rect 800 16664 26200 17064
rect 800 16384 26120 16664
rect 800 15984 26200 16384
rect 800 15848 26120 15984
rect 880 15704 26120 15848
rect 880 15568 26200 15704
rect 800 15304 26200 15568
rect 800 15024 26120 15304
rect 800 14624 26200 15024
rect 800 14344 26120 14624
rect 800 13944 26200 14344
rect 800 13664 26120 13944
rect 800 13536 26200 13664
rect 880 13264 26200 13536
rect 880 13256 26120 13264
rect 800 12984 26120 13256
rect 800 12584 26200 12984
rect 800 12304 26120 12584
rect 800 11904 26200 12304
rect 800 11624 26120 11904
rect 800 11224 26200 11624
rect 880 10944 26120 11224
rect 800 10544 26200 10944
rect 800 10264 26120 10544
rect 800 9864 26200 10264
rect 800 9584 26120 9864
rect 800 9184 26200 9584
rect 800 8912 26120 9184
rect 880 8904 26120 8912
rect 880 8632 26200 8904
rect 800 8504 26200 8632
rect 800 8224 26120 8504
rect 800 7824 26200 8224
rect 800 7544 26120 7824
rect 800 7144 26200 7544
rect 800 6864 26120 7144
rect 800 6600 26200 6864
rect 880 6464 26200 6600
rect 880 6320 26120 6464
rect 800 6184 26120 6320
rect 800 5784 26200 6184
rect 800 5504 26120 5784
rect 800 5104 26200 5504
rect 800 4824 26120 5104
rect 800 4424 26200 4824
rect 800 4288 26120 4424
rect 880 4144 26120 4288
rect 880 4008 26200 4144
rect 800 1976 26200 4008
rect 880 1803 26200 1976
<< metal4 >>
rect 2944 2128 3264 54448
rect 7944 2128 8264 54448
rect 12944 2128 13264 54448
rect 17944 2128 18264 54448
rect 22944 2128 23264 54448
<< obsm4 >>
rect 10547 2891 12864 53957
rect 13344 2891 17864 53957
rect 18344 2891 22864 53957
rect 23344 2891 24597 53957
<< labels >>
rlabel metal4 s 7944 2128 8264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17944 2128 18264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2944 2128 3264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12944 2128 13264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 22944 2128 23264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 54952 800 55072 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 ccff_head_0
port 4 nsew signal input
rlabel metal3 s 26200 4224 27000 4344 6 ccff_tail
port 5 nsew signal output
rlabel metal2 s 938 56200 994 57000 6 ccff_tail_0
port 6 nsew signal output
rlabel metal3 s 26200 25304 27000 25424 6 chanx_right_in[0]
port 7 nsew signal input
rlabel metal3 s 26200 32104 27000 32224 6 chanx_right_in[10]
port 8 nsew signal input
rlabel metal3 s 26200 32784 27000 32904 6 chanx_right_in[11]
port 9 nsew signal input
rlabel metal3 s 26200 33464 27000 33584 6 chanx_right_in[12]
port 10 nsew signal input
rlabel metal3 s 26200 34144 27000 34264 6 chanx_right_in[13]
port 11 nsew signal input
rlabel metal3 s 26200 34824 27000 34944 6 chanx_right_in[14]
port 12 nsew signal input
rlabel metal3 s 26200 35504 27000 35624 6 chanx_right_in[15]
port 13 nsew signal input
rlabel metal3 s 26200 36184 27000 36304 6 chanx_right_in[16]
port 14 nsew signal input
rlabel metal3 s 26200 36864 27000 36984 6 chanx_right_in[17]
port 15 nsew signal input
rlabel metal3 s 26200 37544 27000 37664 6 chanx_right_in[18]
port 16 nsew signal input
rlabel metal3 s 26200 38224 27000 38344 6 chanx_right_in[19]
port 17 nsew signal input
rlabel metal3 s 26200 25984 27000 26104 6 chanx_right_in[1]
port 18 nsew signal input
rlabel metal3 s 26200 38904 27000 39024 6 chanx_right_in[20]
port 19 nsew signal input
rlabel metal3 s 26200 39584 27000 39704 6 chanx_right_in[21]
port 20 nsew signal input
rlabel metal3 s 26200 40264 27000 40384 6 chanx_right_in[22]
port 21 nsew signal input
rlabel metal3 s 26200 40944 27000 41064 6 chanx_right_in[23]
port 22 nsew signal input
rlabel metal3 s 26200 41624 27000 41744 6 chanx_right_in[24]
port 23 nsew signal input
rlabel metal3 s 26200 42304 27000 42424 6 chanx_right_in[25]
port 24 nsew signal input
rlabel metal3 s 26200 42984 27000 43104 6 chanx_right_in[26]
port 25 nsew signal input
rlabel metal3 s 26200 43664 27000 43784 6 chanx_right_in[27]
port 26 nsew signal input
rlabel metal3 s 26200 44344 27000 44464 6 chanx_right_in[28]
port 27 nsew signal input
rlabel metal3 s 26200 45024 27000 45144 6 chanx_right_in[29]
port 28 nsew signal input
rlabel metal3 s 26200 26664 27000 26784 6 chanx_right_in[2]
port 29 nsew signal input
rlabel metal3 s 26200 27344 27000 27464 6 chanx_right_in[3]
port 30 nsew signal input
rlabel metal3 s 26200 28024 27000 28144 6 chanx_right_in[4]
port 31 nsew signal input
rlabel metal3 s 26200 28704 27000 28824 6 chanx_right_in[5]
port 32 nsew signal input
rlabel metal3 s 26200 29384 27000 29504 6 chanx_right_in[6]
port 33 nsew signal input
rlabel metal3 s 26200 30064 27000 30184 6 chanx_right_in[7]
port 34 nsew signal input
rlabel metal3 s 26200 30744 27000 30864 6 chanx_right_in[8]
port 35 nsew signal input
rlabel metal3 s 26200 31424 27000 31544 6 chanx_right_in[9]
port 36 nsew signal input
rlabel metal3 s 26200 4904 27000 5024 6 chanx_right_out[0]
port 37 nsew signal output
rlabel metal3 s 26200 11704 27000 11824 6 chanx_right_out[10]
port 38 nsew signal output
rlabel metal3 s 26200 12384 27000 12504 6 chanx_right_out[11]
port 39 nsew signal output
rlabel metal3 s 26200 13064 27000 13184 6 chanx_right_out[12]
port 40 nsew signal output
rlabel metal3 s 26200 13744 27000 13864 6 chanx_right_out[13]
port 41 nsew signal output
rlabel metal3 s 26200 14424 27000 14544 6 chanx_right_out[14]
port 42 nsew signal output
rlabel metal3 s 26200 15104 27000 15224 6 chanx_right_out[15]
port 43 nsew signal output
rlabel metal3 s 26200 15784 27000 15904 6 chanx_right_out[16]
port 44 nsew signal output
rlabel metal3 s 26200 16464 27000 16584 6 chanx_right_out[17]
port 45 nsew signal output
rlabel metal3 s 26200 17144 27000 17264 6 chanx_right_out[18]
port 46 nsew signal output
rlabel metal3 s 26200 17824 27000 17944 6 chanx_right_out[19]
port 47 nsew signal output
rlabel metal3 s 26200 5584 27000 5704 6 chanx_right_out[1]
port 48 nsew signal output
rlabel metal3 s 26200 18504 27000 18624 6 chanx_right_out[20]
port 49 nsew signal output
rlabel metal3 s 26200 19184 27000 19304 6 chanx_right_out[21]
port 50 nsew signal output
rlabel metal3 s 26200 19864 27000 19984 6 chanx_right_out[22]
port 51 nsew signal output
rlabel metal3 s 26200 20544 27000 20664 6 chanx_right_out[23]
port 52 nsew signal output
rlabel metal3 s 26200 21224 27000 21344 6 chanx_right_out[24]
port 53 nsew signal output
rlabel metal3 s 26200 21904 27000 22024 6 chanx_right_out[25]
port 54 nsew signal output
rlabel metal3 s 26200 22584 27000 22704 6 chanx_right_out[26]
port 55 nsew signal output
rlabel metal3 s 26200 23264 27000 23384 6 chanx_right_out[27]
port 56 nsew signal output
rlabel metal3 s 26200 23944 27000 24064 6 chanx_right_out[28]
port 57 nsew signal output
rlabel metal3 s 26200 24624 27000 24744 6 chanx_right_out[29]
port 58 nsew signal output
rlabel metal3 s 26200 6264 27000 6384 6 chanx_right_out[2]
port 59 nsew signal output
rlabel metal3 s 26200 6944 27000 7064 6 chanx_right_out[3]
port 60 nsew signal output
rlabel metal3 s 26200 7624 27000 7744 6 chanx_right_out[4]
port 61 nsew signal output
rlabel metal3 s 26200 8304 27000 8424 6 chanx_right_out[5]
port 62 nsew signal output
rlabel metal3 s 26200 8984 27000 9104 6 chanx_right_out[6]
port 63 nsew signal output
rlabel metal3 s 26200 9664 27000 9784 6 chanx_right_out[7]
port 64 nsew signal output
rlabel metal3 s 26200 10344 27000 10464 6 chanx_right_out[8]
port 65 nsew signal output
rlabel metal3 s 26200 11024 27000 11144 6 chanx_right_out[9]
port 66 nsew signal output
rlabel metal2 s 1122 0 1178 800 6 chany_bottom_in[0]
port 67 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 chany_bottom_in[10]
port 68 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 chany_bottom_in[11]
port 69 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 chany_bottom_in[12]
port 70 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 chany_bottom_in[13]
port 71 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 chany_bottom_in[14]
port 72 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 chany_bottom_in[15]
port 73 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 chany_bottom_in[16]
port 74 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 chany_bottom_in[17]
port 75 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 chany_bottom_in[18]
port 76 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[19]
port 77 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 chany_bottom_in[1]
port 78 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 chany_bottom_in[20]
port 79 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 chany_bottom_in[21]
port 80 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[22]
port 81 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[23]
port 82 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 chany_bottom_in[24]
port 83 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 chany_bottom_in[25]
port 84 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 chany_bottom_in[26]
port 85 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 chany_bottom_in[27]
port 86 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[28]
port 87 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 chany_bottom_in[29]
port 88 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 chany_bottom_in[2]
port 89 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 chany_bottom_in[3]
port 90 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 chany_bottom_in[4]
port 91 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 chany_bottom_in[5]
port 92 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 chany_bottom_in[6]
port 93 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 chany_bottom_in[7]
port 94 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 chany_bottom_in[8]
port 95 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 chany_bottom_in[9]
port 96 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 chany_bottom_out[0]
port 97 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 chany_bottom_out[10]
port 98 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 chany_bottom_out[11]
port 99 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 chany_bottom_out[12]
port 100 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_out[13]
port 101 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 chany_bottom_out[14]
port 102 nsew signal output
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_out[15]
port 103 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 chany_bottom_out[16]
port 104 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 chany_bottom_out[17]
port 105 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 chany_bottom_out[18]
port 106 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 chany_bottom_out[19]
port 107 nsew signal output
rlabel metal2 s 12530 0 12586 800 6 chany_bottom_out[1]
port 108 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 chany_bottom_out[20]
port 109 nsew signal output
rlabel metal2 s 19890 0 19946 800 6 chany_bottom_out[21]
port 110 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 chany_bottom_out[22]
port 111 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 chany_bottom_out[23]
port 112 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 chany_bottom_out[24]
port 113 nsew signal output
rlabel metal2 s 21362 0 21418 800 6 chany_bottom_out[25]
port 114 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 chany_bottom_out[26]
port 115 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 chany_bottom_out[27]
port 116 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 chany_bottom_out[28]
port 117 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 chany_bottom_out[29]
port 118 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 chany_bottom_out[2]
port 119 nsew signal output
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_out[3]
port 120 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 chany_bottom_out[4]
port 121 nsew signal output
rlabel metal2 s 14002 0 14058 800 6 chany_bottom_out[5]
port 122 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 chany_bottom_out[6]
port 123 nsew signal output
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_out[7]
port 124 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 chany_bottom_out[8]
port 125 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_out[9]
port 126 nsew signal output
rlabel metal2 s 12346 56200 12402 57000 6 chany_top_in_0[0]
port 127 nsew signal input
rlabel metal2 s 16026 56200 16082 57000 6 chany_top_in_0[10]
port 128 nsew signal input
rlabel metal2 s 16394 56200 16450 57000 6 chany_top_in_0[11]
port 129 nsew signal input
rlabel metal2 s 16762 56200 16818 57000 6 chany_top_in_0[12]
port 130 nsew signal input
rlabel metal2 s 17130 56200 17186 57000 6 chany_top_in_0[13]
port 131 nsew signal input
rlabel metal2 s 17498 56200 17554 57000 6 chany_top_in_0[14]
port 132 nsew signal input
rlabel metal2 s 17866 56200 17922 57000 6 chany_top_in_0[15]
port 133 nsew signal input
rlabel metal2 s 18234 56200 18290 57000 6 chany_top_in_0[16]
port 134 nsew signal input
rlabel metal2 s 18602 56200 18658 57000 6 chany_top_in_0[17]
port 135 nsew signal input
rlabel metal2 s 18970 56200 19026 57000 6 chany_top_in_0[18]
port 136 nsew signal input
rlabel metal2 s 19338 56200 19394 57000 6 chany_top_in_0[19]
port 137 nsew signal input
rlabel metal2 s 12714 56200 12770 57000 6 chany_top_in_0[1]
port 138 nsew signal input
rlabel metal2 s 19706 56200 19762 57000 6 chany_top_in_0[20]
port 139 nsew signal input
rlabel metal2 s 20074 56200 20130 57000 6 chany_top_in_0[21]
port 140 nsew signal input
rlabel metal2 s 20442 56200 20498 57000 6 chany_top_in_0[22]
port 141 nsew signal input
rlabel metal2 s 20810 56200 20866 57000 6 chany_top_in_0[23]
port 142 nsew signal input
rlabel metal2 s 21178 56200 21234 57000 6 chany_top_in_0[24]
port 143 nsew signal input
rlabel metal2 s 21546 56200 21602 57000 6 chany_top_in_0[25]
port 144 nsew signal input
rlabel metal2 s 21914 56200 21970 57000 6 chany_top_in_0[26]
port 145 nsew signal input
rlabel metal2 s 22282 56200 22338 57000 6 chany_top_in_0[27]
port 146 nsew signal input
rlabel metal2 s 22650 56200 22706 57000 6 chany_top_in_0[28]
port 147 nsew signal input
rlabel metal2 s 23018 56200 23074 57000 6 chany_top_in_0[29]
port 148 nsew signal input
rlabel metal2 s 13082 56200 13138 57000 6 chany_top_in_0[2]
port 149 nsew signal input
rlabel metal2 s 13450 56200 13506 57000 6 chany_top_in_0[3]
port 150 nsew signal input
rlabel metal2 s 13818 56200 13874 57000 6 chany_top_in_0[4]
port 151 nsew signal input
rlabel metal2 s 14186 56200 14242 57000 6 chany_top_in_0[5]
port 152 nsew signal input
rlabel metal2 s 14554 56200 14610 57000 6 chany_top_in_0[6]
port 153 nsew signal input
rlabel metal2 s 14922 56200 14978 57000 6 chany_top_in_0[7]
port 154 nsew signal input
rlabel metal2 s 15290 56200 15346 57000 6 chany_top_in_0[8]
port 155 nsew signal input
rlabel metal2 s 15658 56200 15714 57000 6 chany_top_in_0[9]
port 156 nsew signal input
rlabel metal2 s 1306 56200 1362 57000 6 chany_top_out_0[0]
port 157 nsew signal output
rlabel metal2 s 4986 56200 5042 57000 6 chany_top_out_0[10]
port 158 nsew signal output
rlabel metal2 s 5354 56200 5410 57000 6 chany_top_out_0[11]
port 159 nsew signal output
rlabel metal2 s 5722 56200 5778 57000 6 chany_top_out_0[12]
port 160 nsew signal output
rlabel metal2 s 6090 56200 6146 57000 6 chany_top_out_0[13]
port 161 nsew signal output
rlabel metal2 s 6458 56200 6514 57000 6 chany_top_out_0[14]
port 162 nsew signal output
rlabel metal2 s 6826 56200 6882 57000 6 chany_top_out_0[15]
port 163 nsew signal output
rlabel metal2 s 7194 56200 7250 57000 6 chany_top_out_0[16]
port 164 nsew signal output
rlabel metal2 s 7562 56200 7618 57000 6 chany_top_out_0[17]
port 165 nsew signal output
rlabel metal2 s 7930 56200 7986 57000 6 chany_top_out_0[18]
port 166 nsew signal output
rlabel metal2 s 8298 56200 8354 57000 6 chany_top_out_0[19]
port 167 nsew signal output
rlabel metal2 s 1674 56200 1730 57000 6 chany_top_out_0[1]
port 168 nsew signal output
rlabel metal2 s 8666 56200 8722 57000 6 chany_top_out_0[20]
port 169 nsew signal output
rlabel metal2 s 9034 56200 9090 57000 6 chany_top_out_0[21]
port 170 nsew signal output
rlabel metal2 s 9402 56200 9458 57000 6 chany_top_out_0[22]
port 171 nsew signal output
rlabel metal2 s 9770 56200 9826 57000 6 chany_top_out_0[23]
port 172 nsew signal output
rlabel metal2 s 10138 56200 10194 57000 6 chany_top_out_0[24]
port 173 nsew signal output
rlabel metal2 s 10506 56200 10562 57000 6 chany_top_out_0[25]
port 174 nsew signal output
rlabel metal2 s 10874 56200 10930 57000 6 chany_top_out_0[26]
port 175 nsew signal output
rlabel metal2 s 11242 56200 11298 57000 6 chany_top_out_0[27]
port 176 nsew signal output
rlabel metal2 s 11610 56200 11666 57000 6 chany_top_out_0[28]
port 177 nsew signal output
rlabel metal2 s 11978 56200 12034 57000 6 chany_top_out_0[29]
port 178 nsew signal output
rlabel metal2 s 2042 56200 2098 57000 6 chany_top_out_0[2]
port 179 nsew signal output
rlabel metal2 s 2410 56200 2466 57000 6 chany_top_out_0[3]
port 180 nsew signal output
rlabel metal2 s 2778 56200 2834 57000 6 chany_top_out_0[4]
port 181 nsew signal output
rlabel metal2 s 3146 56200 3202 57000 6 chany_top_out_0[5]
port 182 nsew signal output
rlabel metal2 s 3514 56200 3570 57000 6 chany_top_out_0[6]
port 183 nsew signal output
rlabel metal2 s 3882 56200 3938 57000 6 chany_top_out_0[7]
port 184 nsew signal output
rlabel metal2 s 4250 56200 4306 57000 6 chany_top_out_0[8]
port 185 nsew signal output
rlabel metal2 s 4618 56200 4674 57000 6 chany_top_out_0[9]
port 186 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 gfpga_pad_io_soc_dir[0]
port 187 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 gfpga_pad_io_soc_dir[1]
port 188 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 gfpga_pad_io_soc_dir[2]
port 189 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 gfpga_pad_io_soc_dir[3]
port 190 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 gfpga_pad_io_soc_in[0]
port 191 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 gfpga_pad_io_soc_in[1]
port 192 nsew signal input
rlabel metal3 s 0 36456 800 36576 6 gfpga_pad_io_soc_in[2]
port 193 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 gfpga_pad_io_soc_in[3]
port 194 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 gfpga_pad_io_soc_out[0]
port 195 nsew signal output
rlabel metal3 s 0 24896 800 25016 6 gfpga_pad_io_soc_out[1]
port 196 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 gfpga_pad_io_soc_out[2]
port 197 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 gfpga_pad_io_soc_out[3]
port 198 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 isol_n
port 199 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 prog_clk
port 200 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 prog_reset_bottom_in
port 201 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 prog_reset_bottom_out
port 202 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 prog_reset_left_in
port 203 nsew signal input
rlabel metal3 s 26200 45704 27000 45824 6 prog_reset_right_out
port 204 nsew signal output
rlabel metal2 s 24490 56200 24546 57000 6 prog_reset_top_in
port 205 nsew signal input
rlabel metal2 s 24122 56200 24178 57000 6 prog_reset_top_out
port 206 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 reset_bottom_in
port 207 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 reset_bottom_out
port 208 nsew signal output
rlabel metal3 s 26200 46384 27000 46504 6 reset_right_in
port 209 nsew signal input
rlabel metal2 s 25226 56200 25282 57000 6 reset_top_in
port 210 nsew signal input
rlabel metal2 s 24858 56200 24914 57000 6 reset_top_out
port 211 nsew signal output
rlabel metal3 s 26200 47064 27000 47184 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 212 nsew signal input
rlabel metal3 s 26200 47744 27000 47864 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 213 nsew signal input
rlabel metal3 s 26200 48424 27000 48544 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 214 nsew signal input
rlabel metal3 s 26200 49104 27000 49224 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 215 nsew signal input
rlabel metal3 s 26200 49784 27000 49904 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 216 nsew signal input
rlabel metal3 s 26200 50464 27000 50584 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 217 nsew signal input
rlabel metal3 s 26200 51144 27000 51264 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 218 nsew signal input
rlabel metal3 s 26200 51824 27000 51944 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 219 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 right_width_0_height_0_subtile_0__pin_inpad_0_
port 220 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 right_width_0_height_0_subtile_1__pin_inpad_0_
port 221 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 right_width_0_height_0_subtile_2__pin_inpad_0_
port 222 nsew signal output
rlabel metal3 s 0 11024 800 11144 6 right_width_0_height_0_subtile_3__pin_inpad_0_
port 223 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 test_enable_bottom_in
port 224 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 test_enable_bottom_out
port 225 nsew signal output
rlabel metal3 s 26200 52504 27000 52624 6 test_enable_right_in
port 226 nsew signal input
rlabel metal2 s 25962 56200 26018 57000 6 test_enable_top_in
port 227 nsew signal input
rlabel metal2 s 25594 56200 25650 57000 6 test_enable_top_out
port 228 nsew signal output
rlabel metal3 s 0 45704 800 45824 6 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 229 nsew signal input
rlabel metal3 s 0 48016 800 48136 6 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 230 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 231 nsew signal input
rlabel metal3 s 0 52640 800 52760 6 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 232 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 27000 57000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2592300
string GDS_FILE /home/hosni/OpenFPGA/clear/openlane/left_tile/runs/23_03_20_14_11/results/signoff/left_tile.magic.gds
string GDS_START 165166
<< end >>

