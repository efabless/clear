magic
tech sky130A
magscale 1 2
timestamp 1656242847
<< viali >>
rect 1869 20553 1903 20587
rect 2237 20553 2271 20587
rect 2973 20553 3007 20587
rect 3617 20553 3651 20587
rect 6653 20553 6687 20587
rect 9413 20553 9447 20587
rect 15025 20553 15059 20587
rect 15761 20553 15795 20587
rect 16129 20553 16163 20587
rect 16865 20553 16899 20587
rect 17601 20553 17635 20587
rect 17969 20553 18003 20587
rect 18429 20553 18463 20587
rect 18889 20553 18923 20587
rect 8769 20485 8803 20519
rect 12642 20485 12676 20519
rect 19441 20485 19475 20519
rect 1685 20417 1719 20451
rect 2053 20417 2087 20451
rect 2421 20417 2455 20451
rect 2605 20417 2639 20451
rect 3065 20417 3099 20451
rect 3433 20417 3467 20451
rect 3893 20417 3927 20451
rect 4169 20417 4203 20451
rect 5273 20417 5307 20451
rect 6193 20417 6227 20451
rect 6469 20417 6503 20451
rect 7665 20417 7699 20451
rect 8953 20417 8987 20451
rect 9321 20417 9355 20451
rect 10425 20417 10459 20451
rect 11345 20417 11379 20451
rect 14105 20417 14139 20451
rect 14473 20417 14507 20451
rect 14841 20417 14875 20451
rect 15209 20417 15243 20451
rect 15577 20417 15611 20451
rect 15945 20417 15979 20451
rect 16681 20417 16715 20451
rect 17049 20417 17083 20451
rect 17417 20417 17451 20451
rect 17785 20417 17819 20451
rect 18245 20417 18279 20451
rect 18705 20417 18739 20451
rect 19533 20417 19567 20451
rect 20637 20417 20671 20451
rect 4997 20349 5031 20383
rect 5917 20349 5951 20383
rect 6745 20349 6779 20383
rect 7021 20349 7055 20383
rect 7941 20349 7975 20383
rect 10149 20349 10183 20383
rect 11069 20349 11103 20383
rect 12909 20349 12943 20383
rect 13553 20349 13587 20383
rect 13829 20349 13863 20383
rect 19809 20349 19843 20383
rect 20821 20349 20855 20383
rect 2789 20281 2823 20315
rect 3249 20281 3283 20315
rect 9137 20281 9171 20315
rect 14657 20281 14691 20315
rect 15393 20281 15427 20315
rect 17233 20281 17267 20315
rect 1501 20213 1535 20247
rect 4077 20213 4111 20247
rect 4353 20213 4387 20247
rect 11529 20213 11563 20247
rect 14289 20213 14323 20247
rect 2697 20009 2731 20043
rect 3801 20009 3835 20043
rect 4169 20009 4203 20043
rect 4445 20009 4479 20043
rect 4997 20009 5031 20043
rect 5273 20009 5307 20043
rect 6009 20009 6043 20043
rect 6193 20009 6227 20043
rect 7481 20009 7515 20043
rect 8769 20009 8803 20043
rect 9597 20009 9631 20043
rect 13001 20009 13035 20043
rect 13369 20009 13403 20043
rect 13829 20009 13863 20043
rect 18705 20009 18739 20043
rect 3157 19941 3191 19975
rect 7757 19941 7791 19975
rect 14289 19941 14323 19975
rect 14565 19941 14599 19975
rect 18981 19941 19015 19975
rect 19441 19941 19475 19975
rect 19809 19941 19843 19975
rect 2973 19873 3007 19907
rect 6285 19873 6319 19907
rect 10517 19873 10551 19907
rect 11437 19873 11471 19907
rect 1685 19805 1719 19839
rect 2053 19805 2087 19839
rect 2145 19805 2179 19839
rect 2421 19805 2455 19839
rect 2881 19805 2915 19839
rect 5365 19805 5399 19839
rect 6561 19805 6595 19839
rect 7297 19805 7331 19839
rect 7573 19805 7607 19839
rect 8033 19805 8067 19839
rect 8217 19805 8251 19839
rect 8585 19805 8619 19839
rect 9413 19805 9447 19839
rect 10241 19805 10275 19839
rect 11161 19805 11195 19839
rect 12909 19805 12943 19839
rect 13185 19805 13219 19839
rect 13737 19805 13771 19839
rect 14105 19805 14139 19839
rect 14381 19805 14415 19839
rect 14841 19805 14875 19839
rect 16313 19805 16347 19839
rect 18797 19805 18831 19839
rect 19257 19805 19291 19839
rect 19625 19805 19659 19839
rect 21557 19805 21591 19839
rect 5825 19737 5859 19771
rect 9045 19737 9079 19771
rect 9229 19737 9263 19771
rect 12642 19737 12676 19771
rect 21290 19737 21324 19771
rect 1501 19669 1535 19703
rect 1869 19669 1903 19703
rect 2329 19669 2363 19703
rect 2605 19669 2639 19703
rect 5549 19669 5583 19703
rect 7849 19669 7883 19703
rect 8309 19669 8343 19703
rect 11529 19669 11563 19703
rect 13553 19669 13587 19703
rect 14657 19669 14691 19703
rect 16221 19669 16255 19703
rect 16497 19669 16531 19703
rect 19993 19669 20027 19703
rect 20177 19669 20211 19703
rect 1961 19465 1995 19499
rect 2697 19465 2731 19499
rect 6377 19465 6411 19499
rect 7113 19465 7147 19499
rect 8309 19465 8343 19499
rect 9781 19465 9815 19499
rect 10057 19465 10091 19499
rect 10701 19465 10735 19499
rect 11253 19465 11287 19499
rect 21005 19465 21039 19499
rect 21373 19465 21407 19499
rect 1685 19329 1719 19363
rect 1777 19329 1811 19363
rect 2053 19329 2087 19363
rect 2329 19329 2363 19363
rect 7205 19329 7239 19363
rect 8125 19329 8159 19363
rect 8401 19329 8435 19363
rect 9045 19329 9079 19363
rect 9321 19329 9355 19363
rect 9597 19329 9631 19363
rect 9873 19329 9907 19363
rect 10241 19329 10275 19363
rect 10517 19329 10551 19363
rect 11069 19329 11103 19363
rect 11713 19329 11747 19363
rect 11897 19329 11931 19363
rect 12164 19329 12198 19363
rect 19616 19329 19650 19363
rect 20821 19329 20855 19363
rect 21189 19329 21223 19363
rect 7665 19261 7699 19295
rect 8861 19261 8895 19295
rect 13553 19261 13587 19295
rect 19349 19261 19383 19295
rect 2513 19193 2547 19227
rect 6929 19193 6963 19227
rect 7757 19193 7791 19227
rect 8033 19193 8067 19227
rect 9505 19193 9539 19227
rect 10425 19193 10459 19227
rect 13277 19193 13311 19227
rect 13461 19193 13495 19227
rect 13829 19193 13863 19227
rect 1501 19125 1535 19159
rect 2237 19125 2271 19159
rect 6745 19125 6779 19159
rect 7389 19125 7423 19159
rect 8585 19125 8619 19159
rect 8769 19125 8803 19159
rect 9229 19125 9263 19159
rect 10885 19125 10919 19159
rect 11621 19125 11655 19159
rect 19165 19125 19199 19159
rect 20729 19125 20763 19159
rect 7573 18921 7607 18955
rect 8217 18921 8251 18955
rect 9689 18921 9723 18955
rect 21189 18921 21223 18955
rect 9413 18853 9447 18887
rect 2053 18785 2087 18819
rect 8033 18785 8067 18819
rect 13185 18785 13219 18819
rect 13369 18785 13403 18819
rect 1685 18717 1719 18751
rect 1777 18717 1811 18751
rect 8309 18717 8343 18751
rect 8677 18717 8711 18751
rect 8953 18717 8987 18751
rect 9505 18717 9539 18751
rect 9781 18717 9815 18751
rect 10057 18717 10091 18751
rect 11529 18717 11563 18751
rect 14749 18717 14783 18751
rect 16313 18717 16347 18751
rect 16681 18717 16715 18751
rect 18245 18717 18279 18751
rect 18337 18717 18371 18751
rect 20646 18717 20680 18751
rect 20913 18717 20947 18751
rect 21005 18717 21039 18751
rect 7481 18649 7515 18683
rect 10324 18649 10358 18683
rect 11796 18649 11830 18683
rect 14994 18649 15028 18683
rect 18000 18649 18034 18683
rect 21373 18649 21407 18683
rect 1501 18581 1535 18615
rect 1961 18581 1995 18615
rect 8493 18581 8527 18615
rect 9137 18581 9171 18615
rect 9965 18581 9999 18615
rect 11437 18581 11471 18615
rect 12909 18581 12943 18615
rect 16129 18581 16163 18615
rect 16865 18581 16899 18615
rect 19533 18581 19567 18615
rect 2145 18377 2179 18411
rect 5549 18377 5583 18411
rect 8677 18377 8711 18411
rect 9781 18377 9815 18411
rect 10517 18377 10551 18411
rect 21097 18377 21131 18411
rect 21465 18377 21499 18411
rect 5641 18309 5675 18343
rect 6561 18309 6595 18343
rect 10793 18309 10827 18343
rect 11345 18309 11379 18343
rect 14657 18309 14691 18343
rect 1685 18241 1719 18275
rect 2053 18241 2087 18275
rect 2329 18241 2363 18275
rect 8585 18241 8619 18275
rect 9229 18225 9263 18259
rect 9505 18241 9539 18275
rect 9965 18241 9999 18275
rect 10885 18241 10919 18275
rect 12653 18241 12687 18275
rect 12920 18241 12954 18275
rect 14206 18241 14240 18275
rect 14473 18241 14507 18275
rect 16230 18241 16264 18275
rect 16497 18241 16531 18275
rect 17794 18241 17828 18275
rect 19266 18241 19300 18275
rect 19533 18241 19567 18275
rect 20738 18241 20772 18275
rect 21005 18241 21039 18275
rect 21281 18241 21315 18275
rect 5733 18173 5767 18207
rect 6377 18173 6411 18207
rect 7941 18173 7975 18207
rect 8861 18173 8895 18207
rect 18061 18173 18095 18207
rect 1869 18105 1903 18139
rect 9689 18105 9723 18139
rect 15117 18105 15151 18139
rect 19625 18105 19659 18139
rect 1501 18037 1535 18071
rect 5181 18037 5215 18071
rect 7757 18037 7791 18071
rect 8217 18037 8251 18071
rect 9413 18037 9447 18071
rect 10149 18037 10183 18071
rect 11529 18037 11563 18071
rect 13093 18037 13127 18071
rect 16681 18037 16715 18071
rect 18153 18037 18187 18071
rect 8585 17833 8619 17867
rect 13185 17833 13219 17867
rect 13553 17833 13587 17867
rect 13461 17765 13495 17799
rect 17877 17765 17911 17799
rect 5181 17697 5215 17731
rect 5365 17697 5399 17731
rect 6377 17697 6411 17731
rect 6469 17697 6503 17731
rect 8033 17697 8067 17731
rect 13093 17697 13127 17731
rect 1685 17629 1719 17663
rect 6285 17629 6319 17663
rect 16497 17629 16531 17663
rect 17969 17629 18003 17663
rect 18153 17629 18187 17663
rect 19625 17629 19659 17663
rect 19809 17629 19843 17663
rect 21281 17629 21315 17663
rect 8217 17561 8251 17595
rect 12826 17561 12860 17595
rect 16764 17561 16798 17595
rect 20076 17561 20110 17595
rect 1501 17493 1535 17527
rect 5457 17493 5491 17527
rect 5825 17493 5859 17527
rect 5917 17493 5951 17527
rect 8125 17493 8159 17527
rect 9505 17493 9539 17527
rect 9873 17493 9907 17527
rect 11713 17493 11747 17527
rect 21189 17493 21223 17527
rect 21465 17493 21499 17527
rect 2145 17289 2179 17323
rect 2605 17289 2639 17323
rect 2881 17289 2915 17323
rect 3249 17289 3283 17323
rect 4445 17289 4479 17323
rect 4905 17289 4939 17323
rect 5457 17289 5491 17323
rect 5917 17289 5951 17323
rect 6929 17289 6963 17323
rect 7389 17289 7423 17323
rect 7941 17289 7975 17323
rect 8309 17289 8343 17323
rect 8677 17289 8711 17323
rect 9137 17289 9171 17323
rect 9229 17289 9263 17323
rect 9597 17289 9631 17323
rect 10057 17289 10091 17323
rect 15117 17289 15151 17323
rect 18153 17289 18187 17323
rect 4537 17221 4571 17255
rect 7021 17221 7055 17255
rect 7849 17221 7883 17255
rect 12664 17221 12698 17255
rect 13268 17221 13302 17255
rect 14473 17221 14507 17255
rect 16230 17221 16264 17255
rect 20453 17221 20487 17255
rect 21281 17221 21315 17255
rect 1685 17153 1719 17187
rect 2329 17153 2363 17187
rect 2789 17153 2823 17187
rect 3065 17153 3099 17187
rect 3433 17153 3467 17187
rect 3709 17153 3743 17187
rect 5549 17153 5583 17187
rect 8493 17153 8527 17187
rect 9965 17153 9999 17187
rect 12909 17153 12943 17187
rect 13001 17153 13035 17187
rect 17805 17153 17839 17187
rect 18061 17153 18095 17187
rect 18981 17153 19015 17187
rect 19237 17153 19271 17187
rect 4353 17085 4387 17119
rect 5273 17085 5307 17119
rect 6837 17085 6871 17119
rect 7757 17085 7791 17119
rect 9413 17085 9447 17119
rect 10241 17085 10275 17119
rect 16497 17085 16531 17119
rect 3525 17017 3559 17051
rect 8769 17017 8803 17051
rect 11529 17017 11563 17051
rect 1501 16949 1535 16983
rect 10425 16949 10459 16983
rect 14381 16949 14415 16983
rect 16681 16949 16715 16983
rect 20361 16949 20395 16983
rect 2973 16745 3007 16779
rect 3433 16745 3467 16779
rect 4721 16745 4755 16779
rect 16037 16745 16071 16779
rect 18429 16745 18463 16779
rect 4077 16609 4111 16643
rect 4261 16609 4295 16643
rect 6193 16609 6227 16643
rect 7573 16609 7607 16643
rect 7757 16609 7791 16643
rect 8125 16609 8159 16643
rect 9689 16609 9723 16643
rect 10977 16609 11011 16643
rect 13277 16609 13311 16643
rect 18337 16609 18371 16643
rect 1685 16541 1719 16575
rect 2053 16541 2087 16575
rect 3157 16541 3191 16575
rect 3249 16541 3283 16575
rect 4353 16541 4387 16575
rect 8309 16541 8343 16575
rect 9229 16541 9263 16575
rect 9505 16541 9539 16575
rect 9965 16541 9999 16575
rect 11253 16541 11287 16575
rect 13021 16541 13055 16575
rect 13553 16541 13587 16575
rect 15761 16541 15795 16575
rect 16589 16541 16623 16575
rect 20637 16541 20671 16575
rect 20729 16541 20763 16575
rect 21465 16541 21499 16575
rect 7021 16473 7055 16507
rect 7481 16473 7515 16507
rect 15494 16473 15528 16507
rect 18070 16473 18104 16507
rect 20370 16473 20404 16507
rect 1501 16405 1535 16439
rect 1869 16405 1903 16439
rect 5549 16405 5583 16439
rect 5917 16405 5951 16439
rect 6009 16405 6043 16439
rect 7113 16405 7147 16439
rect 8217 16405 8251 16439
rect 8677 16405 8711 16439
rect 9045 16405 9079 16439
rect 9321 16405 9355 16439
rect 9873 16405 9907 16439
rect 10333 16405 10367 16439
rect 10425 16405 10459 16439
rect 10793 16405 10827 16439
rect 10885 16405 10919 16439
rect 11897 16405 11931 16439
rect 13461 16405 13495 16439
rect 14381 16405 14415 16439
rect 15853 16405 15887 16439
rect 16957 16405 16991 16439
rect 19257 16405 19291 16439
rect 2973 16201 3007 16235
rect 3433 16201 3467 16235
rect 5273 16201 5307 16235
rect 6101 16201 6135 16235
rect 7757 16201 7791 16235
rect 8401 16201 8435 16235
rect 9781 16201 9815 16235
rect 10609 16201 10643 16235
rect 11069 16201 11103 16235
rect 17969 16201 18003 16235
rect 6837 16133 6871 16167
rect 8861 16133 8895 16167
rect 10701 16133 10735 16167
rect 11529 16133 11563 16167
rect 13286 16133 13320 16167
rect 15301 16133 15335 16167
rect 1685 16065 1719 16099
rect 3157 16065 3191 16099
rect 3617 16065 3651 16099
rect 5733 16065 5767 16099
rect 6929 16065 6963 16099
rect 7849 16065 7883 16099
rect 9597 16065 9631 16099
rect 13553 16065 13587 16099
rect 13645 16065 13679 16099
rect 14953 16065 14987 16099
rect 19082 16065 19116 16099
rect 19349 16065 19383 16099
rect 19441 16065 19475 16099
rect 21198 16065 21232 16099
rect 21465 16065 21499 16099
rect 5457 15997 5491 16031
rect 5641 15997 5675 16031
rect 6745 15997 6779 16031
rect 7665 15997 7699 16031
rect 9965 15997 9999 16031
rect 10517 15997 10551 16031
rect 11161 15997 11195 16031
rect 15209 15997 15243 16031
rect 7297 15929 7331 15963
rect 12173 15929 12207 15963
rect 13829 15929 13863 15963
rect 1501 15861 1535 15895
rect 6377 15861 6411 15895
rect 8217 15861 8251 15895
rect 9229 15861 9263 15895
rect 9413 15861 9447 15895
rect 10149 15861 10183 15895
rect 15577 15861 15611 15895
rect 20085 15861 20119 15895
rect 1869 15657 1903 15691
rect 2237 15657 2271 15691
rect 2513 15657 2547 15691
rect 5181 15657 5215 15691
rect 6009 15657 6043 15691
rect 6101 15657 6135 15691
rect 8953 15657 8987 15691
rect 9873 15657 9907 15691
rect 16313 15657 16347 15691
rect 8401 15589 8435 15623
rect 10241 15589 10275 15623
rect 4537 15521 4571 15555
rect 4721 15521 4755 15555
rect 5365 15521 5399 15555
rect 6561 15521 6595 15555
rect 6745 15521 6779 15555
rect 7757 15521 7791 15555
rect 7941 15521 7975 15555
rect 9505 15521 9539 15555
rect 10885 15521 10919 15555
rect 13369 15521 13403 15555
rect 1685 15453 1719 15487
rect 2053 15453 2087 15487
rect 2421 15453 2455 15487
rect 2697 15453 2731 15487
rect 9321 15453 9355 15487
rect 10609 15453 10643 15487
rect 15485 15453 15519 15487
rect 15577 15453 15611 15487
rect 17693 15453 17727 15487
rect 17785 15453 17819 15487
rect 21557 15453 21591 15487
rect 4813 15385 4847 15419
rect 5641 15385 5675 15419
rect 13124 15385 13158 15419
rect 15218 15385 15252 15419
rect 15761 15385 15795 15419
rect 17426 15385 17460 15419
rect 21290 15385 21324 15419
rect 1501 15317 1535 15351
rect 3801 15317 3835 15351
rect 5549 15317 5583 15351
rect 6469 15317 6503 15351
rect 8033 15317 8067 15351
rect 9413 15317 9447 15351
rect 9965 15317 9999 15351
rect 10701 15317 10735 15351
rect 11989 15317 12023 15351
rect 13553 15317 13587 15351
rect 14105 15317 14139 15351
rect 19809 15317 19843 15351
rect 19993 15317 20027 15351
rect 20177 15317 20211 15351
rect 2145 15113 2179 15147
rect 2605 15113 2639 15147
rect 3341 15113 3375 15147
rect 4997 15113 5031 15147
rect 7481 15113 7515 15147
rect 7849 15113 7883 15147
rect 8953 15113 8987 15147
rect 9045 15113 9079 15147
rect 9505 15113 9539 15147
rect 10609 15113 10643 15147
rect 11069 15113 11103 15147
rect 8309 15045 8343 15079
rect 16948 15045 16982 15079
rect 1685 14977 1719 15011
rect 2053 14977 2087 15011
rect 2329 14977 2363 15011
rect 2789 14977 2823 15011
rect 4169 14977 4203 15011
rect 7113 14977 7147 15011
rect 7757 14977 7791 15011
rect 8217 14977 8251 15011
rect 9873 14977 9907 15011
rect 10977 14977 11011 15011
rect 13194 14977 13228 15011
rect 15034 14977 15068 15011
rect 15301 14977 15335 15011
rect 15393 14977 15427 15011
rect 16681 14977 16715 15011
rect 18153 14977 18187 15011
rect 19461 14977 19495 15011
rect 19717 14977 19751 15011
rect 21014 14977 21048 15011
rect 3065 14909 3099 14943
rect 3249 14909 3283 14943
rect 3893 14909 3927 14943
rect 4077 14909 4111 14943
rect 4721 14909 4755 14943
rect 4905 14909 4939 14943
rect 5457 14909 5491 14943
rect 6929 14909 6963 14943
rect 7021 14909 7055 14943
rect 8401 14909 8435 14943
rect 8861 14909 8895 14943
rect 9965 14909 9999 14943
rect 10149 14909 10183 14943
rect 11253 14909 11287 14943
rect 13461 14909 13495 14943
rect 21281 14909 21315 14943
rect 1869 14841 1903 14875
rect 12081 14841 12115 14875
rect 13645 14841 13679 14875
rect 1501 14773 1535 14807
rect 3709 14773 3743 14807
rect 4537 14773 4571 14807
rect 5365 14773 5399 14807
rect 6009 14773 6043 14807
rect 9413 14773 9447 14807
rect 10425 14773 10459 14807
rect 13921 14773 13955 14807
rect 16129 14773 16163 14807
rect 18061 14773 18095 14807
rect 18337 14773 18371 14807
rect 19901 14773 19935 14807
rect 21373 14773 21407 14807
rect 4629 14569 4663 14603
rect 6653 14569 6687 14603
rect 9873 14569 9907 14603
rect 15945 14569 15979 14603
rect 16221 14569 16255 14603
rect 8401 14501 8435 14535
rect 4077 14433 4111 14467
rect 5089 14433 5123 14467
rect 6101 14433 6135 14467
rect 6193 14433 6227 14467
rect 7481 14433 7515 14467
rect 8033 14433 8067 14467
rect 8125 14433 8159 14467
rect 9321 14433 9355 14467
rect 10425 14433 10459 14467
rect 10517 14433 10551 14467
rect 13553 14433 13587 14467
rect 13737 14433 13771 14467
rect 15853 14433 15887 14467
rect 1685 14365 1719 14399
rect 4261 14365 4295 14399
rect 5181 14365 5215 14399
rect 5273 14365 5307 14399
rect 9505 14365 9539 14399
rect 10333 14365 10367 14399
rect 15586 14365 15620 14399
rect 17601 14365 17635 14399
rect 17693 14365 17727 14399
rect 18153 14365 18187 14399
rect 21097 14365 21131 14399
rect 21189 14365 21223 14399
rect 4813 14297 4847 14331
rect 7941 14297 7975 14331
rect 9413 14297 9447 14331
rect 13286 14297 13320 14331
rect 17356 14297 17390 14331
rect 20852 14297 20886 14331
rect 1501 14229 1535 14263
rect 4169 14229 4203 14263
rect 5641 14229 5675 14263
rect 6285 14229 6319 14263
rect 7573 14229 7607 14263
rect 9965 14229 9999 14263
rect 12173 14229 12207 14263
rect 14473 14229 14507 14263
rect 19717 14229 19751 14263
rect 5365 14025 5399 14059
rect 5733 14025 5767 14059
rect 6377 14025 6411 14059
rect 7297 14025 7331 14059
rect 9321 14025 9355 14059
rect 10517 14025 10551 14059
rect 11253 14025 11287 14059
rect 18153 14025 18187 14059
rect 21557 14025 21591 14059
rect 6837 13957 6871 13991
rect 7665 13957 7699 13991
rect 9229 13957 9263 13991
rect 16926 13957 16960 13991
rect 1685 13889 1719 13923
rect 6745 13889 6779 13923
rect 7757 13889 7791 13923
rect 9689 13889 9723 13923
rect 11069 13889 11103 13923
rect 12532 13889 12566 13923
rect 15025 13889 15059 13923
rect 15281 13889 15315 13923
rect 16681 13889 16715 13923
rect 19266 13889 19300 13923
rect 20433 13889 20467 13923
rect 5089 13821 5123 13855
rect 5273 13821 5307 13855
rect 6101 13821 6135 13855
rect 6929 13821 6963 13855
rect 7849 13821 7883 13855
rect 9781 13821 9815 13855
rect 9965 13821 9999 13855
rect 10241 13821 10275 13855
rect 10425 13821 10459 13855
rect 12265 13821 12299 13855
rect 19533 13821 19567 13855
rect 19625 13821 19659 13855
rect 20177 13821 20211 13855
rect 13645 13753 13679 13787
rect 13829 13753 13863 13787
rect 16405 13753 16439 13787
rect 18061 13753 18095 13787
rect 1501 13685 1535 13719
rect 10885 13685 10919 13719
rect 4537 13481 4571 13515
rect 7941 13481 7975 13515
rect 9413 13481 9447 13515
rect 19257 13481 19291 13515
rect 7113 13413 7147 13447
rect 8033 13413 8067 13447
rect 16129 13413 16163 13447
rect 18981 13413 19015 13447
rect 6193 13345 6227 13379
rect 6469 13345 6503 13379
rect 6653 13345 6687 13379
rect 7389 13345 7423 13379
rect 7481 13345 7515 13379
rect 8677 13345 8711 13379
rect 10057 13345 10091 13379
rect 10793 13345 10827 13379
rect 11713 13345 11747 13379
rect 17509 13345 17543 13379
rect 17601 13345 17635 13379
rect 1685 13277 1719 13311
rect 2053 13277 2087 13311
rect 4721 13277 4755 13311
rect 9781 13277 9815 13311
rect 10701 13277 10735 13311
rect 11529 13277 11563 13311
rect 12541 13277 12575 13311
rect 12808 13277 12842 13311
rect 17242 13277 17276 13311
rect 21281 13277 21315 13311
rect 21465 13277 21499 13311
rect 6745 13209 6779 13243
rect 8493 13209 8527 13243
rect 10609 13209 10643 13243
rect 17846 13209 17880 13243
rect 21014 13209 21048 13243
rect 1501 13141 1535 13175
rect 1869 13141 1903 13175
rect 7573 13141 7607 13175
rect 8401 13141 8435 13175
rect 9873 13141 9907 13175
rect 10241 13141 10275 13175
rect 11069 13141 11103 13175
rect 11437 13141 11471 13175
rect 13921 13141 13955 13175
rect 14105 13141 14139 13175
rect 15945 13141 15979 13175
rect 19901 13141 19935 13175
rect 1869 12937 1903 12971
rect 3157 12937 3191 12971
rect 4261 12937 4295 12971
rect 5089 12937 5123 12971
rect 5457 12937 5491 12971
rect 5917 12937 5951 12971
rect 6377 12937 6411 12971
rect 6745 12937 6779 12971
rect 7297 12937 7331 12971
rect 8585 12937 8619 12971
rect 9965 12937 9999 12971
rect 10425 12937 10459 12971
rect 18153 12937 18187 12971
rect 18337 12937 18371 12971
rect 20821 12937 20855 12971
rect 21373 12937 21407 12971
rect 6837 12869 6871 12903
rect 7941 12869 7975 12903
rect 13849 12869 13883 12903
rect 15669 12869 15703 12903
rect 16926 12869 16960 12903
rect 20462 12869 20496 12903
rect 1409 12801 1443 12835
rect 1685 12801 1719 12835
rect 1961 12801 1995 12835
rect 3341 12801 3375 12835
rect 4445 12801 4479 12835
rect 4997 12801 5031 12835
rect 5825 12801 5859 12835
rect 7573 12801 7607 12835
rect 8033 12801 8067 12835
rect 8953 12801 8987 12835
rect 10333 12801 10367 12835
rect 14105 12801 14139 12835
rect 15310 12801 15344 12835
rect 15577 12801 15611 12835
rect 16681 12801 16715 12835
rect 20729 12801 20763 12835
rect 2145 12733 2179 12767
rect 5273 12733 5307 12767
rect 6101 12733 6135 12767
rect 7021 12733 7055 12767
rect 7757 12733 7791 12767
rect 9045 12733 9079 12767
rect 9229 12733 9263 12767
rect 10609 12733 10643 12767
rect 1593 12665 1627 12699
rect 4629 12665 4663 12699
rect 8401 12665 8435 12699
rect 18061 12665 18095 12699
rect 12633 12597 12667 12631
rect 12725 12597 12759 12631
rect 14197 12597 14231 12631
rect 19349 12597 19383 12631
rect 1869 12393 1903 12427
rect 4905 12393 4939 12427
rect 5641 12393 5675 12427
rect 7481 12393 7515 12427
rect 8953 12393 8987 12427
rect 10241 12393 10275 12427
rect 18245 12393 18279 12427
rect 8401 12325 8435 12359
rect 15301 12325 15335 12359
rect 18153 12325 18187 12359
rect 19809 12325 19843 12359
rect 6285 12257 6319 12291
rect 8125 12257 8159 12291
rect 9597 12257 9631 12291
rect 9781 12257 9815 12291
rect 10885 12257 10919 12291
rect 16681 12257 16715 12291
rect 16773 12257 16807 12291
rect 1409 12189 1443 12223
rect 1685 12189 1719 12223
rect 2053 12189 2087 12223
rect 5089 12189 5123 12223
rect 10701 12189 10735 12223
rect 12182 12189 12216 12223
rect 12449 12189 12483 12223
rect 12541 12189 12575 12223
rect 17040 12189 17074 12223
rect 20922 12189 20956 12223
rect 21189 12189 21223 12223
rect 7941 12121 7975 12155
rect 8677 12121 8711 12155
rect 12808 12121 12842 12155
rect 16436 12121 16470 12155
rect 1593 12053 1627 12087
rect 6009 12053 6043 12087
rect 6101 12053 6135 12087
rect 7849 12053 7883 12087
rect 9321 12053 9355 12087
rect 9413 12053 9447 12087
rect 10609 12053 10643 12087
rect 11069 12053 11103 12087
rect 13921 12053 13955 12087
rect 14197 12053 14231 12087
rect 14381 12053 14415 12087
rect 21281 12053 21315 12087
rect 3985 11849 4019 11883
rect 6377 11849 6411 11883
rect 7297 11849 7331 11883
rect 8401 11849 8435 11883
rect 9781 11849 9815 11883
rect 10149 11849 10183 11883
rect 10517 11849 10551 11883
rect 11529 11849 11563 11883
rect 12541 11849 12575 11883
rect 5549 11781 5583 11815
rect 20821 11781 20855 11815
rect 1409 11713 1443 11747
rect 1685 11713 1719 11747
rect 1961 11713 1995 11747
rect 4169 11713 4203 11747
rect 6745 11713 6779 11747
rect 8033 11713 8067 11747
rect 9689 11713 9723 11747
rect 10609 11713 10643 11747
rect 11897 11713 11931 11747
rect 12449 11713 12483 11747
rect 13654 11713 13688 11747
rect 16241 11713 16275 11747
rect 16497 11713 16531 11747
rect 16773 11713 16807 11747
rect 16957 11713 16991 11747
rect 17141 11713 17175 11747
rect 17509 11713 17543 11747
rect 17765 11713 17799 11747
rect 19616 11713 19650 11747
rect 2145 11645 2179 11679
rect 5089 11645 5123 11679
rect 6837 11645 6871 11679
rect 7021 11645 7055 11679
rect 7757 11645 7791 11679
rect 7941 11645 7975 11679
rect 9965 11645 9999 11679
rect 10793 11645 10827 11679
rect 11161 11645 11195 11679
rect 11989 11645 12023 11679
rect 12081 11645 12115 11679
rect 13921 11645 13955 11679
rect 19349 11645 19383 11679
rect 9321 11577 9355 11611
rect 18981 11577 19015 11611
rect 1593 11509 1627 11543
rect 1869 11509 1903 11543
rect 6009 11509 6043 11543
rect 6193 11509 6227 11543
rect 11345 11509 11379 11543
rect 14013 11509 14047 11543
rect 15117 11509 15151 11543
rect 18889 11509 18923 11543
rect 20729 11509 20763 11543
rect 1869 11305 1903 11339
rect 2145 11305 2179 11339
rect 5365 11305 5399 11339
rect 6193 11305 6227 11339
rect 7021 11305 7055 11339
rect 7389 11305 7423 11339
rect 16589 11305 16623 11339
rect 19625 11305 19659 11339
rect 1593 11237 1627 11271
rect 8953 11237 8987 11271
rect 10057 11237 10091 11271
rect 10977 11237 11011 11271
rect 11253 11237 11287 11271
rect 13001 11237 13035 11271
rect 16681 11237 16715 11271
rect 4813 11169 4847 11203
rect 5641 11169 5675 11203
rect 6377 11169 6411 11203
rect 9597 11169 9631 11203
rect 9965 11169 9999 11203
rect 10517 11169 10551 11203
rect 10609 11169 10643 11203
rect 15209 11169 15243 11203
rect 18337 11169 18371 11203
rect 21005 11169 21039 11203
rect 21097 11169 21131 11203
rect 1409 11101 1443 11135
rect 1685 11101 1719 11135
rect 2053 11101 2087 11135
rect 2329 11101 2363 11135
rect 4997 11101 5031 11135
rect 10425 11101 10459 11135
rect 11529 11101 11563 11135
rect 18061 11101 18095 11135
rect 4445 11033 4479 11067
rect 4905 11033 4939 11067
rect 5733 11033 5767 11067
rect 5825 11033 5859 11067
rect 7113 11033 7147 11067
rect 9321 11033 9355 11067
rect 11437 11033 11471 11067
rect 11796 11033 11830 11067
rect 15476 11033 15510 11067
rect 17816 11033 17850 11067
rect 20738 11033 20772 11067
rect 6561 10965 6595 10999
rect 6653 10965 6687 10999
rect 8585 10965 8619 10999
rect 9413 10965 9447 10999
rect 12909 10965 12943 10999
rect 13277 10965 13311 10999
rect 13461 10965 13495 10999
rect 18153 10965 18187 10999
rect 18613 10965 18647 10999
rect 5089 10761 5123 10795
rect 5457 10761 5491 10795
rect 5917 10761 5951 10795
rect 8217 10761 8251 10795
rect 8677 10761 8711 10795
rect 9045 10761 9079 10795
rect 9137 10761 9171 10795
rect 9505 10761 9539 10795
rect 10333 10761 10367 10795
rect 13645 10761 13679 10795
rect 19993 10761 20027 10795
rect 6745 10693 6779 10727
rect 7205 10693 7239 10727
rect 8585 10693 8619 10727
rect 10793 10693 10827 10727
rect 15761 10693 15795 10727
rect 15945 10693 15979 10727
rect 21106 10693 21140 10727
rect 1409 10625 1443 10659
rect 1685 10625 1719 10659
rect 4721 10625 4755 10659
rect 5549 10625 5583 10659
rect 6009 10625 6043 10659
rect 7849 10625 7883 10659
rect 9597 10625 9631 10659
rect 10701 10625 10735 10659
rect 11161 10625 11195 10659
rect 12653 10625 12687 10659
rect 12909 10625 12943 10659
rect 13185 10625 13219 10659
rect 15402 10625 15436 10659
rect 15669 10625 15703 10659
rect 16681 10625 16715 10659
rect 16937 10625 16971 10659
rect 18685 10625 18719 10659
rect 4537 10557 4571 10591
rect 4629 10557 4663 10591
rect 5365 10557 5399 10591
rect 6469 10557 6503 10591
rect 6653 10557 6687 10591
rect 7573 10557 7607 10591
rect 7757 10557 7791 10591
rect 8493 10557 8527 10591
rect 9689 10557 9723 10591
rect 9965 10557 9999 10591
rect 10885 10557 10919 10591
rect 13369 10557 13403 10591
rect 18429 10557 18463 10591
rect 21373 10557 21407 10591
rect 21465 10557 21499 10591
rect 13001 10489 13035 10523
rect 18153 10489 18187 10523
rect 1593 10421 1627 10455
rect 7113 10421 7147 10455
rect 11529 10421 11563 10455
rect 14289 10421 14323 10455
rect 18061 10421 18095 10455
rect 19809 10421 19843 10455
rect 2145 10217 2179 10251
rect 3157 10217 3191 10251
rect 3341 10217 3375 10251
rect 4813 10217 4847 10251
rect 5641 10217 5675 10251
rect 7205 10217 7239 10251
rect 7297 10217 7331 10251
rect 8309 10217 8343 10251
rect 8953 10217 8987 10251
rect 11713 10217 11747 10251
rect 1593 10149 1627 10183
rect 2605 10081 2639 10115
rect 3893 10081 3927 10115
rect 4077 10081 4111 10115
rect 5549 10081 5583 10115
rect 6101 10081 6135 10115
rect 6285 10081 6319 10115
rect 6653 10081 6687 10115
rect 7849 10081 7883 10115
rect 9505 10081 9539 10115
rect 13093 10081 13127 10115
rect 13277 10081 13311 10115
rect 1409 10013 1443 10047
rect 1685 10013 1719 10047
rect 1961 10013 1995 10047
rect 2329 10013 2363 10047
rect 4721 10013 4755 10047
rect 4997 10013 5031 10047
rect 6745 10013 6779 10047
rect 7665 10013 7699 10047
rect 8217 10013 8251 10047
rect 9321 10013 9355 10047
rect 10149 10013 10183 10047
rect 14197 10013 14231 10047
rect 14453 10013 14487 10047
rect 17049 10013 17083 10047
rect 17141 10013 17175 10047
rect 19257 10013 19291 10047
rect 19513 10013 19547 10047
rect 3617 9945 3651 9979
rect 4169 9945 4203 9979
rect 6837 9945 6871 9979
rect 10394 9945 10428 9979
rect 12848 9945 12882 9979
rect 16782 9945 16816 9979
rect 17386 9945 17420 9979
rect 18613 9945 18647 9979
rect 18797 9945 18831 9979
rect 1869 9877 1903 9911
rect 2697 9877 2731 9911
rect 2789 9877 2823 9911
rect 4537 9877 4571 9911
rect 6009 9877 6043 9911
rect 7757 9877 7791 9911
rect 8585 9877 8619 9911
rect 9413 9877 9447 9911
rect 9781 9877 9815 9911
rect 11529 9877 11563 9911
rect 15577 9877 15611 9911
rect 15669 9877 15703 9911
rect 18521 9877 18555 9911
rect 20637 9877 20671 9911
rect 20821 9877 20855 9911
rect 21465 9877 21499 9911
rect 1409 9673 1443 9707
rect 2881 9673 2915 9707
rect 21189 9673 21223 9707
rect 21373 9673 21407 9707
rect 4905 9605 4939 9639
rect 5457 9605 5491 9639
rect 6653 9605 6687 9639
rect 7205 9605 7239 9639
rect 9321 9605 9355 9639
rect 10793 9605 10827 9639
rect 13492 9605 13526 9639
rect 18398 9605 18432 9639
rect 1777 9537 1811 9571
rect 2053 9537 2087 9571
rect 2329 9537 2363 9571
rect 2605 9537 2639 9571
rect 6745 9537 6779 9571
rect 10333 9537 10367 9571
rect 10425 9537 10459 9571
rect 11161 9537 11195 9571
rect 14942 9537 14976 9571
rect 15209 9537 15243 9571
rect 16037 9537 16071 9571
rect 17805 9537 17839 9571
rect 20841 9537 20875 9571
rect 21097 9537 21131 9571
rect 4629 9469 4663 9503
rect 4813 9469 4847 9503
rect 5549 9469 5583 9503
rect 6469 9469 6503 9503
rect 9137 9469 9171 9503
rect 9229 9469 9263 9503
rect 10609 9469 10643 9503
rect 11897 9469 11931 9503
rect 13737 9469 13771 9503
rect 15853 9469 15887 9503
rect 18061 9469 18095 9503
rect 18153 9469 18187 9503
rect 1593 9401 1627 9435
rect 1869 9401 1903 9435
rect 2145 9401 2179 9435
rect 2421 9401 2455 9435
rect 5273 9401 5307 9435
rect 7113 9401 7147 9435
rect 9689 9401 9723 9435
rect 16681 9401 16715 9435
rect 19533 9401 19567 9435
rect 2789 9333 2823 9367
rect 8769 9333 8803 9367
rect 9781 9333 9815 9367
rect 9965 9333 9999 9367
rect 11069 9333 11103 9367
rect 11713 9333 11747 9367
rect 12357 9333 12391 9367
rect 13829 9333 13863 9367
rect 15301 9333 15335 9367
rect 19717 9333 19751 9367
rect 2145 9129 2179 9163
rect 3065 9129 3099 9163
rect 3341 9129 3375 9163
rect 3893 9129 3927 9163
rect 6101 9129 6135 9163
rect 9689 9129 9723 9163
rect 1593 9061 1627 9095
rect 2973 9061 3007 9095
rect 7021 9061 7055 9095
rect 13461 9061 13495 9095
rect 2421 8993 2455 9027
rect 4629 8993 4663 9027
rect 4813 8993 4847 9027
rect 5549 8993 5583 9027
rect 6837 8993 6871 9027
rect 7665 8993 7699 9027
rect 8493 8993 8527 9027
rect 10149 8993 10183 9027
rect 10333 8993 10367 9027
rect 11069 8993 11103 9027
rect 12081 8993 12115 9027
rect 1409 8925 1443 8959
rect 1685 8925 1719 8959
rect 1961 8925 1995 8959
rect 2605 8925 2639 8959
rect 3249 8925 3283 8959
rect 4077 8925 4111 8959
rect 4905 8925 4939 8959
rect 10977 8925 11011 8959
rect 13829 8925 13863 8959
rect 14105 8925 14139 8959
rect 15577 8925 15611 8959
rect 16313 8925 16347 8959
rect 17785 8925 17819 8959
rect 18153 8925 18187 8959
rect 20646 8925 20680 8959
rect 20913 8925 20947 8959
rect 21005 8925 21039 8959
rect 7389 8857 7423 8891
rect 10885 8857 10919 8891
rect 11345 8857 11379 8891
rect 12348 8857 12382 8891
rect 14372 8857 14406 8891
rect 16580 8857 16614 8891
rect 1869 8789 1903 8823
rect 2513 8789 2547 8823
rect 5273 8789 5307 8823
rect 5641 8789 5675 8823
rect 5733 8789 5767 8823
rect 6193 8789 6227 8823
rect 6561 8789 6595 8823
rect 6653 8789 6687 8823
rect 7481 8789 7515 8823
rect 7849 8789 7883 8823
rect 8217 8789 8251 8823
rect 8309 8789 8343 8823
rect 8769 8789 8803 8823
rect 10057 8789 10091 8823
rect 10517 8789 10551 8823
rect 13645 8789 13679 8823
rect 15485 8789 15519 8823
rect 17693 8789 17727 8823
rect 19533 8789 19567 8823
rect 1685 8585 1719 8619
rect 2697 8585 2731 8619
rect 4353 8585 4387 8619
rect 6193 8585 6227 8619
rect 8033 8585 8067 8619
rect 8585 8585 8619 8619
rect 9965 8585 9999 8619
rect 10517 8585 10551 8619
rect 13829 8585 13863 8619
rect 13921 8585 13955 8619
rect 15577 8585 15611 8619
rect 15761 8585 15795 8619
rect 7297 8517 7331 8551
rect 8125 8517 8159 8551
rect 9413 8517 9447 8551
rect 20729 8517 20763 8551
rect 1409 8449 1443 8483
rect 2237 8449 2271 8483
rect 2881 8449 2915 8483
rect 3065 8449 3099 8483
rect 4445 8449 4479 8483
rect 5825 8449 5859 8483
rect 8953 8449 8987 8483
rect 10057 8449 10091 8483
rect 10885 8449 10919 8483
rect 11529 8449 11563 8483
rect 13378 8449 13412 8483
rect 13645 8449 13679 8483
rect 14197 8449 14231 8483
rect 14453 8449 14487 8483
rect 19165 8449 19199 8483
rect 19432 8449 19466 8483
rect 1961 8381 1995 8415
rect 2145 8381 2179 8415
rect 4261 8381 4295 8415
rect 4905 8381 4939 8415
rect 5549 8381 5583 8415
rect 5733 8381 5767 8415
rect 6377 8381 6411 8415
rect 7389 8381 7423 8415
rect 7573 8381 7607 8415
rect 7941 8381 7975 8415
rect 9045 8381 9079 8415
rect 9229 8381 9263 8415
rect 9873 8381 9907 8415
rect 10977 8381 11011 8415
rect 11069 8381 11103 8415
rect 2605 8313 2639 8347
rect 6929 8313 6963 8347
rect 8493 8313 8527 8347
rect 10425 8313 10459 8347
rect 12265 8313 12299 8347
rect 1593 8245 1627 8279
rect 4813 8245 4847 8279
rect 5273 8245 5307 8279
rect 20545 8245 20579 8279
rect 2605 8041 2639 8075
rect 5457 8041 5491 8075
rect 6469 8041 6503 8075
rect 7573 8041 7607 8075
rect 7849 8041 7883 8075
rect 8677 8041 8711 8075
rect 14841 8041 14875 8075
rect 19441 8041 19475 8075
rect 20913 8041 20947 8075
rect 1593 7973 1627 8007
rect 2513 7973 2547 8007
rect 6101 7973 6135 8007
rect 11897 7973 11931 8007
rect 14381 7973 14415 8007
rect 1961 7905 1995 7939
rect 2881 7905 2915 7939
rect 5733 7905 5767 7939
rect 7113 7905 7147 7939
rect 8493 7905 8527 7939
rect 10425 7905 10459 7939
rect 11253 7905 11287 7939
rect 12449 7905 12483 7939
rect 12817 7905 12851 7939
rect 16681 7905 16715 7939
rect 18521 7905 18555 7939
rect 20821 7905 20855 7939
rect 1409 7837 1443 7871
rect 2789 7837 2823 7871
rect 5641 7837 5675 7871
rect 6285 7837 6319 7871
rect 10149 7837 10183 7871
rect 11345 7837 11379 7871
rect 15761 7837 15795 7871
rect 18337 7837 18371 7871
rect 2053 7769 2087 7803
rect 2145 7769 2179 7803
rect 6837 7769 6871 7803
rect 8217 7769 8251 7803
rect 11437 7769 11471 7803
rect 16405 7769 16439 7803
rect 18245 7769 18279 7803
rect 20554 7769 20588 7803
rect 21097 7769 21131 7803
rect 5917 7701 5951 7735
rect 6929 7701 6963 7735
rect 7297 7701 7331 7735
rect 8309 7701 8343 7735
rect 9781 7701 9815 7735
rect 10241 7701 10275 7735
rect 11805 7701 11839 7735
rect 12265 7701 12299 7735
rect 12357 7701 12391 7735
rect 14289 7701 14323 7735
rect 15853 7701 15887 7735
rect 16037 7701 16071 7735
rect 16497 7701 16531 7735
rect 17509 7701 17543 7735
rect 17693 7701 17727 7735
rect 17877 7701 17911 7735
rect 2145 7497 2179 7531
rect 4905 7497 4939 7531
rect 6193 7497 6227 7531
rect 6837 7497 6871 7531
rect 7481 7497 7515 7531
rect 9045 7497 9079 7531
rect 9597 7497 9631 7531
rect 10517 7497 10551 7531
rect 12081 7497 12115 7531
rect 13461 7497 13495 7531
rect 14657 7497 14691 7531
rect 14749 7497 14783 7531
rect 15577 7497 15611 7531
rect 19349 7497 19383 7531
rect 20821 7497 20855 7531
rect 1961 7429 1995 7463
rect 4997 7429 5031 7463
rect 9505 7429 9539 7463
rect 10977 7429 11011 7463
rect 1409 7361 1443 7395
rect 1685 7361 1719 7395
rect 2329 7361 2363 7395
rect 5825 7361 5859 7395
rect 7297 7361 7331 7395
rect 7849 7361 7883 7395
rect 7941 7361 7975 7395
rect 8677 7361 8711 7395
rect 10885 7361 10919 7395
rect 11529 7361 11563 7395
rect 12449 7361 12483 7395
rect 12909 7361 12943 7395
rect 13829 7361 13863 7395
rect 15485 7361 15519 7395
rect 20462 7361 20496 7395
rect 20729 7361 20763 7395
rect 4813 7293 4847 7327
rect 5549 7293 5583 7327
rect 5733 7293 5767 7327
rect 6929 7293 6963 7327
rect 7113 7293 7147 7327
rect 8125 7293 8159 7327
rect 8493 7293 8527 7327
rect 8585 7293 8619 7327
rect 9689 7293 9723 7327
rect 11069 7293 11103 7327
rect 12541 7293 12575 7327
rect 12725 7293 12759 7327
rect 13921 7293 13955 7327
rect 14105 7293 14139 7327
rect 14933 7293 14967 7327
rect 15761 7293 15795 7327
rect 1593 7225 1627 7259
rect 1869 7225 1903 7259
rect 6469 7225 6503 7259
rect 14289 7225 14323 7259
rect 5365 7157 5399 7191
rect 9137 7157 9171 7191
rect 10057 7157 10091 7191
rect 11897 7157 11931 7191
rect 15117 7157 15151 7191
rect 1961 6953 1995 6987
rect 6469 6953 6503 6987
rect 7297 6953 7331 6987
rect 8401 6953 8435 6987
rect 9321 6953 9355 6987
rect 10149 6953 10183 6987
rect 14105 6953 14139 6987
rect 1593 6885 1627 6919
rect 4077 6817 4111 6851
rect 4169 6817 4203 6851
rect 7113 6817 7147 6851
rect 7849 6817 7883 6851
rect 8953 6817 8987 6851
rect 9229 6817 9263 6851
rect 9781 6817 9815 6851
rect 9873 6817 9907 6851
rect 10793 6817 10827 6851
rect 11989 6817 12023 6851
rect 14749 6817 14783 6851
rect 1409 6749 1443 6783
rect 1685 6749 1719 6783
rect 2145 6749 2179 6783
rect 4261 6749 4295 6783
rect 6101 6749 6135 6783
rect 6837 6749 6871 6783
rect 8033 6749 8067 6783
rect 9689 6749 9723 6783
rect 14565 6749 14599 6783
rect 2329 6681 2363 6715
rect 10517 6681 10551 6715
rect 12081 6681 12115 6715
rect 1869 6613 1903 6647
rect 4629 6613 4663 6647
rect 4721 6613 4755 6647
rect 5457 6613 5491 6647
rect 6285 6613 6319 6647
rect 6929 6613 6963 6647
rect 7573 6613 7607 6647
rect 7941 6613 7975 6647
rect 8585 6613 8619 6647
rect 10609 6613 10643 6647
rect 12173 6613 12207 6647
rect 12541 6613 12575 6647
rect 14473 6613 14507 6647
rect 14933 6613 14967 6647
rect 1593 6409 1627 6443
rect 2053 6409 2087 6443
rect 4353 6409 4387 6443
rect 4813 6409 4847 6443
rect 7113 6409 7147 6443
rect 7481 6409 7515 6443
rect 7941 6409 7975 6443
rect 8769 6409 8803 6443
rect 9229 6409 9263 6443
rect 9965 6409 9999 6443
rect 12265 6409 12299 6443
rect 21373 6409 21407 6443
rect 1961 6341 1995 6375
rect 4445 6341 4479 6375
rect 5733 6341 5767 6375
rect 10057 6341 10091 6375
rect 1409 6273 1443 6307
rect 5273 6273 5307 6307
rect 7021 6273 7055 6307
rect 8309 6273 8343 6307
rect 9137 6273 9171 6307
rect 10977 6273 11011 6307
rect 12633 6273 12667 6307
rect 14289 6273 14323 6307
rect 21281 6273 21315 6307
rect 21557 6273 21591 6307
rect 1869 6205 1903 6239
rect 4261 6205 4295 6239
rect 5089 6205 5123 6239
rect 5181 6205 5215 6239
rect 7573 6205 7607 6239
rect 7757 6205 7791 6239
rect 8401 6205 8435 6239
rect 8585 6205 8619 6239
rect 9321 6205 9355 6239
rect 9873 6205 9907 6239
rect 10701 6205 10735 6239
rect 10885 6205 10919 6239
rect 11897 6205 11931 6239
rect 12725 6205 12759 6239
rect 12909 6205 12943 6239
rect 14013 6205 14047 6239
rect 14197 6205 14231 6239
rect 5641 6137 5675 6171
rect 2421 6069 2455 6103
rect 10425 6069 10459 6103
rect 11345 6069 11379 6103
rect 11713 6069 11747 6103
rect 14657 6069 14691 6103
rect 1961 5865 1995 5899
rect 7205 5865 7239 5899
rect 8769 5865 8803 5899
rect 13277 5865 13311 5899
rect 1593 5797 1627 5831
rect 1869 5797 1903 5831
rect 11161 5797 11195 5831
rect 17325 5797 17359 5831
rect 5825 5729 5859 5763
rect 5917 5729 5951 5763
rect 6653 5729 6687 5763
rect 8125 5729 8159 5763
rect 9689 5729 9723 5763
rect 10609 5729 10643 5763
rect 11529 5729 11563 5763
rect 12725 5729 12759 5763
rect 16681 5729 16715 5763
rect 17601 5729 17635 5763
rect 20085 5729 20119 5763
rect 1409 5661 1443 5695
rect 1685 5661 1719 5695
rect 2513 5661 2547 5695
rect 6009 5661 6043 5695
rect 8401 5661 8435 5695
rect 10793 5661 10827 5695
rect 11805 5661 11839 5695
rect 13369 5661 13403 5695
rect 17693 5661 17727 5695
rect 2697 5593 2731 5627
rect 6837 5593 6871 5627
rect 8309 5593 8343 5627
rect 9505 5593 9539 5627
rect 16957 5593 16991 5627
rect 20361 5593 20395 5627
rect 2237 5525 2271 5559
rect 4905 5525 4939 5559
rect 5273 5525 5307 5559
rect 6377 5525 6411 5559
rect 6745 5525 6779 5559
rect 7297 5525 7331 5559
rect 7941 5525 7975 5559
rect 8953 5525 8987 5559
rect 9137 5525 9171 5559
rect 9597 5525 9631 5559
rect 10701 5525 10735 5559
rect 11713 5525 11747 5559
rect 12173 5525 12207 5559
rect 12817 5525 12851 5559
rect 12909 5525 12943 5559
rect 13553 5525 13587 5559
rect 16865 5525 16899 5559
rect 17785 5525 17819 5559
rect 18153 5525 18187 5559
rect 20269 5525 20303 5559
rect 20729 5525 20763 5559
rect 2237 5321 2271 5355
rect 2605 5321 2639 5355
rect 6653 5321 6687 5355
rect 7113 5321 7147 5355
rect 8309 5321 8343 5355
rect 9321 5321 9355 5355
rect 9689 5321 9723 5355
rect 10149 5321 10183 5355
rect 10977 5321 11011 5355
rect 11897 5321 11931 5355
rect 13185 5321 13219 5355
rect 13553 5321 13587 5355
rect 17233 5321 17267 5355
rect 2145 5253 2179 5287
rect 4629 5253 4663 5287
rect 5549 5253 5583 5287
rect 11989 5253 12023 5287
rect 15393 5253 15427 5287
rect 1501 5185 1535 5219
rect 2697 5185 2731 5219
rect 4721 5185 4755 5219
rect 6745 5185 6779 5219
rect 9781 5185 9815 5219
rect 10609 5185 10643 5219
rect 12817 5185 12851 5219
rect 13277 5185 13311 5219
rect 15853 5185 15887 5219
rect 20821 5185 20855 5219
rect 2053 5117 2087 5151
rect 4537 5117 4571 5151
rect 5273 5117 5307 5151
rect 5457 5117 5491 5151
rect 6009 5117 6043 5151
rect 6561 5117 6595 5151
rect 8401 5117 8435 5151
rect 8493 5117 8527 5151
rect 9505 5117 9539 5151
rect 10333 5117 10367 5151
rect 10517 5117 10551 5151
rect 11805 5117 11839 5151
rect 12541 5117 12575 5151
rect 12725 5117 12759 5151
rect 15485 5117 15519 5151
rect 15577 5117 15611 5151
rect 1685 5049 1719 5083
rect 5089 5049 5123 5083
rect 5917 5049 5951 5083
rect 7941 5049 7975 5083
rect 12357 5049 12391 5083
rect 7757 4981 7791 5015
rect 11161 4981 11195 5015
rect 13461 4981 13495 5015
rect 15025 4981 15059 5015
rect 16037 4981 16071 5015
rect 20637 4981 20671 5015
rect 5825 4777 5859 4811
rect 6285 4777 6319 4811
rect 7113 4777 7147 4811
rect 8493 4777 8527 4811
rect 9045 4777 9079 4811
rect 9781 4777 9815 4811
rect 11437 4777 11471 4811
rect 12357 4777 12391 4811
rect 15485 4777 15519 4811
rect 18061 4777 18095 4811
rect 10977 4709 11011 4743
rect 11253 4709 11287 4743
rect 11621 4709 11655 4743
rect 16773 4709 16807 4743
rect 1961 4641 1995 4675
rect 5181 4641 5215 4675
rect 6929 4641 6963 4675
rect 7849 4641 7883 4675
rect 8677 4641 8711 4675
rect 9689 4641 9723 4675
rect 10425 4641 10459 4675
rect 14841 4641 14875 4675
rect 15025 4641 15059 4675
rect 16037 4641 16071 4675
rect 16405 4641 16439 4675
rect 17509 4641 17543 4675
rect 2237 4573 2271 4607
rect 2329 4573 2363 4607
rect 5457 4573 5491 4607
rect 8033 4573 8067 4607
rect 10241 4573 10275 4607
rect 10609 4573 10643 4607
rect 11897 4573 11931 4607
rect 14749 4573 14783 4607
rect 16589 4573 16623 4607
rect 16865 4573 16899 4607
rect 18797 4573 18831 4607
rect 5365 4505 5399 4539
rect 6653 4505 6687 4539
rect 8125 4505 8159 4539
rect 10793 4505 10827 4539
rect 5917 4437 5951 4471
rect 6745 4437 6779 4471
rect 7297 4437 7331 4471
rect 9413 4437 9447 4471
rect 10149 4437 10183 4471
rect 11713 4437 11747 4471
rect 12081 4437 12115 4471
rect 14381 4437 14415 4471
rect 15853 4437 15887 4471
rect 15945 4437 15979 4471
rect 17601 4437 17635 4471
rect 17693 4437 17727 4471
rect 18981 4437 19015 4471
rect 5825 4233 5859 4267
rect 8953 4233 8987 4267
rect 10057 4233 10091 4267
rect 10517 4233 10551 4267
rect 11897 4233 11931 4267
rect 11989 4233 12023 4267
rect 12449 4233 12483 4267
rect 16681 4233 16715 4267
rect 17601 4233 17635 4267
rect 18521 4233 18555 4267
rect 6745 4165 6779 4199
rect 7757 4165 7791 4199
rect 8493 4165 8527 4199
rect 9321 4165 9355 4199
rect 17049 4165 17083 4199
rect 1961 4097 1995 4131
rect 7665 4097 7699 4131
rect 8585 4097 8619 4131
rect 10149 4097 10183 4131
rect 10885 4097 10919 4131
rect 10977 4097 11011 4131
rect 14381 4097 14415 4131
rect 16313 4097 16347 4131
rect 17969 4097 18003 4131
rect 2237 4029 2271 4063
rect 2513 4029 2547 4063
rect 5641 4029 5675 4063
rect 5733 4029 5767 4063
rect 6837 4029 6871 4063
rect 7021 4029 7055 4063
rect 7573 4029 7607 4063
rect 8401 4029 8435 4063
rect 9229 4029 9263 4063
rect 10241 4029 10275 4063
rect 11161 4029 11195 4063
rect 12173 4029 12207 4063
rect 12725 4029 12759 4063
rect 16129 4029 16163 4063
rect 17141 4029 17175 4063
rect 17325 4029 17359 4063
rect 18061 4029 18095 4063
rect 18245 4029 18279 4063
rect 9689 3961 9723 3995
rect 11529 3961 11563 3995
rect 2329 3893 2363 3927
rect 2789 3893 2823 3927
rect 2973 3893 3007 3927
rect 6193 3893 6227 3927
rect 6377 3893 6411 3927
rect 8125 3893 8159 3927
rect 9505 3893 9539 3927
rect 12633 3893 12667 3927
rect 12909 3893 12943 3927
rect 14565 3893 14599 3927
rect 2697 3689 2731 3723
rect 7113 3689 7147 3723
rect 10517 3689 10551 3723
rect 12449 3689 12483 3723
rect 14105 3689 14139 3723
rect 17233 3689 17267 3723
rect 18429 3689 18463 3723
rect 19993 3689 20027 3723
rect 21373 3689 21407 3723
rect 1685 3621 1719 3655
rect 2053 3621 2087 3655
rect 2605 3621 2639 3655
rect 4813 3621 4847 3655
rect 9689 3621 9723 3655
rect 17417 3621 17451 3655
rect 4261 3553 4295 3587
rect 5549 3553 5583 3587
rect 6561 3553 6595 3587
rect 9137 3553 9171 3587
rect 9229 3553 9263 3587
rect 9873 3553 9907 3587
rect 10057 3553 10091 3587
rect 10701 3553 10735 3587
rect 11529 3553 11563 3587
rect 12541 3553 12575 3587
rect 12817 3553 12851 3587
rect 13185 3553 13219 3587
rect 1501 3485 1535 3519
rect 2145 3485 2179 3519
rect 2421 3485 2455 3519
rect 6745 3485 6779 3519
rect 7389 3485 7423 3519
rect 8309 3485 8343 3519
rect 8585 3485 8619 3519
rect 9321 3485 9355 3519
rect 11805 3485 11839 3519
rect 12265 3485 12299 3519
rect 13369 3485 13403 3519
rect 13829 3485 13863 3519
rect 21281 3485 21315 3519
rect 21557 3485 21591 3519
rect 1869 3417 1903 3451
rect 3065 3417 3099 3451
rect 4445 3417 4479 3451
rect 5273 3417 5307 3451
rect 8217 3417 8251 3451
rect 8769 3417 8803 3451
rect 10885 3417 10919 3451
rect 13277 3417 13311 3451
rect 14289 3417 14323 3451
rect 2329 3349 2363 3383
rect 2881 3349 2915 3383
rect 3249 3349 3283 3383
rect 3433 3349 3467 3383
rect 4353 3349 4387 3383
rect 4905 3349 4939 3383
rect 5365 3349 5399 3383
rect 5733 3349 5767 3383
rect 6653 3349 6687 3383
rect 7297 3349 7331 3383
rect 7573 3349 7607 3383
rect 7757 3349 7791 3383
rect 8033 3349 8067 3383
rect 10149 3349 10183 3383
rect 10977 3349 11011 3383
rect 11345 3349 11379 3383
rect 11713 3349 11747 3383
rect 12173 3349 12207 3383
rect 13737 3349 13771 3383
rect 2881 3145 2915 3179
rect 4261 3145 4295 3179
rect 4629 3145 4663 3179
rect 7389 3145 7423 3179
rect 7757 3145 7791 3179
rect 8493 3145 8527 3179
rect 8953 3145 8987 3179
rect 10057 3145 10091 3179
rect 12449 3145 12483 3179
rect 12909 3145 12943 3179
rect 14841 3145 14875 3179
rect 17693 3145 17727 3179
rect 17969 3145 18003 3179
rect 18245 3145 18279 3179
rect 19073 3145 19107 3179
rect 2421 3077 2455 3111
rect 3801 3077 3835 3111
rect 11253 3077 11287 3111
rect 12817 3077 12851 3111
rect 15209 3077 15243 3111
rect 15945 3077 15979 3111
rect 17233 3077 17267 3111
rect 2697 3009 2731 3043
rect 2973 3009 3007 3043
rect 3249 3009 3283 3043
rect 7849 3009 7883 3043
rect 8217 3009 8251 3043
rect 8861 3009 8895 3043
rect 9689 3009 9723 3043
rect 10149 3009 10183 3043
rect 10425 3009 10459 3043
rect 11529 3009 11563 3043
rect 11805 3009 11839 3043
rect 13461 3009 13495 3043
rect 13553 3009 13587 3043
rect 13829 3009 13863 3043
rect 14105 3009 14139 3043
rect 14381 3009 14415 3043
rect 14657 3009 14691 3043
rect 14933 3009 14967 3043
rect 15485 3009 15519 3043
rect 15669 3009 15703 3043
rect 16129 3009 16163 3043
rect 16681 3009 16715 3043
rect 16957 3009 16991 3043
rect 18061 3009 18095 3043
rect 18521 3009 18555 3043
rect 18613 3009 18647 3043
rect 18889 3009 18923 3043
rect 19349 3009 19383 3043
rect 19625 3009 19659 3043
rect 19901 3009 19935 3043
rect 20361 3009 20395 3043
rect 20729 3009 20763 3043
rect 20913 3009 20947 3043
rect 21281 3009 21315 3043
rect 1961 2941 1995 2975
rect 2237 2941 2271 2975
rect 4721 2941 4755 2975
rect 4905 2941 4939 2975
rect 5089 2941 5123 2975
rect 5365 2941 5399 2975
rect 6193 2941 6227 2975
rect 6469 2941 6503 2975
rect 6745 2941 6779 2975
rect 8033 2941 8067 2975
rect 9137 2941 9171 2975
rect 9413 2941 9447 2975
rect 9597 2941 9631 2975
rect 13001 2941 13035 2975
rect 3433 2873 3467 2907
rect 3709 2873 3743 2907
rect 4169 2873 4203 2907
rect 8401 2873 8435 2907
rect 11069 2873 11103 2907
rect 14013 2873 14047 2907
rect 14289 2873 14323 2907
rect 15117 2873 15151 2907
rect 15853 2873 15887 2907
rect 16865 2873 16899 2907
rect 19165 2873 19199 2907
rect 19441 2873 19475 2907
rect 20177 2873 20211 2907
rect 21097 2873 21131 2907
rect 2513 2805 2547 2839
rect 3157 2805 3191 2839
rect 13277 2805 13311 2839
rect 13737 2805 13771 2839
rect 14565 2805 14599 2839
rect 16313 2805 16347 2839
rect 17141 2805 17175 2839
rect 18337 2805 18371 2839
rect 18797 2805 18831 2839
rect 20085 2805 20119 2839
rect 20545 2805 20579 2839
rect 21465 2805 21499 2839
rect 2973 2601 3007 2635
rect 3985 2601 4019 2635
rect 4813 2601 4847 2635
rect 5273 2601 5307 2635
rect 10149 2601 10183 2635
rect 10425 2601 10459 2635
rect 12127 2601 12161 2635
rect 14289 2601 14323 2635
rect 4353 2533 4387 2567
rect 14657 2533 14691 2567
rect 19717 2533 19751 2567
rect 1961 2465 1995 2499
rect 3065 2465 3099 2499
rect 5917 2465 5951 2499
rect 7205 2465 7239 2499
rect 9505 2465 9539 2499
rect 9689 2465 9723 2499
rect 11345 2465 11379 2499
rect 12449 2465 12483 2499
rect 2237 2397 2271 2431
rect 2329 2397 2363 2431
rect 2789 2397 2823 2431
rect 3249 2397 3283 2431
rect 3801 2397 3835 2431
rect 4169 2397 4203 2431
rect 4629 2397 4663 2431
rect 5089 2397 5123 2431
rect 6193 2397 6227 2431
rect 6929 2397 6963 2431
rect 7849 2397 7883 2431
rect 8125 2397 8159 2431
rect 10241 2397 10275 2431
rect 11069 2397 11103 2431
rect 12357 2397 12391 2431
rect 12725 2397 12759 2431
rect 13369 2397 13403 2431
rect 13737 2397 13771 2431
rect 14105 2397 14139 2431
rect 14473 2397 14507 2431
rect 14841 2397 14875 2431
rect 15209 2397 15243 2431
rect 15669 2397 15703 2431
rect 16129 2397 16163 2431
rect 16681 2397 16715 2431
rect 17325 2397 17359 2431
rect 17509 2397 17543 2431
rect 18245 2397 18279 2431
rect 18705 2397 18739 2431
rect 19533 2397 19567 2431
rect 19901 2397 19935 2431
rect 19993 2397 20027 2431
rect 20361 2397 20395 2431
rect 20729 2397 20763 2431
rect 21189 2397 21223 2431
rect 2697 2329 2731 2363
rect 3617 2329 3651 2363
rect 6469 2329 6503 2363
rect 6653 2329 6687 2363
rect 9137 2329 9171 2363
rect 2513 2261 2547 2295
rect 3433 2261 3467 2295
rect 4537 2261 4571 2295
rect 4997 2261 5031 2295
rect 6745 2261 6779 2295
rect 9229 2261 9263 2295
rect 9781 2261 9815 2295
rect 13553 2261 13587 2295
rect 13921 2261 13955 2295
rect 15025 2261 15059 2295
rect 15393 2261 15427 2295
rect 15853 2261 15887 2295
rect 16313 2261 16347 2295
rect 16865 2261 16899 2295
rect 17141 2261 17175 2295
rect 17693 2261 17727 2295
rect 18061 2261 18095 2295
rect 18521 2261 18555 2295
rect 19349 2261 19383 2295
rect 20177 2261 20211 2295
rect 20545 2261 20579 2295
rect 20913 2261 20947 2295
rect 21373 2261 21407 2295
<< metal1 >>
rect 10502 20952 10508 21004
rect 10560 20992 10566 21004
rect 15194 20992 15200 21004
rect 10560 20964 15200 20992
rect 10560 20952 10566 20964
rect 15194 20952 15200 20964
rect 15252 20952 15258 21004
rect 11790 20884 11796 20936
rect 11848 20924 11854 20936
rect 14090 20924 14096 20936
rect 11848 20896 14096 20924
rect 11848 20884 11854 20896
rect 14090 20884 14096 20896
rect 14148 20884 14154 20936
rect 11882 20816 11888 20868
rect 11940 20856 11946 20868
rect 12802 20856 12808 20868
rect 11940 20828 12808 20856
rect 11940 20816 11946 20828
rect 12802 20816 12808 20828
rect 12860 20816 12866 20868
rect 12158 20748 12164 20800
rect 12216 20788 12222 20800
rect 13906 20788 13912 20800
rect 12216 20760 13912 20788
rect 12216 20748 12222 20760
rect 13906 20748 13912 20760
rect 13964 20748 13970 20800
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 1854 20584 1860 20596
rect 1815 20556 1860 20584
rect 1854 20544 1860 20556
rect 1912 20544 1918 20596
rect 2222 20584 2228 20596
rect 2183 20556 2228 20584
rect 2222 20544 2228 20556
rect 2280 20544 2286 20596
rect 2958 20584 2964 20596
rect 2919 20556 2964 20584
rect 2958 20544 2964 20556
rect 3016 20544 3022 20596
rect 3605 20587 3663 20593
rect 3605 20553 3617 20587
rect 3651 20584 3663 20587
rect 4154 20584 4160 20596
rect 3651 20556 4160 20584
rect 3651 20553 3663 20556
rect 3605 20547 3663 20553
rect 4154 20544 4160 20556
rect 4212 20544 4218 20596
rect 6641 20587 6699 20593
rect 6641 20553 6653 20587
rect 6687 20584 6699 20587
rect 6822 20584 6828 20596
rect 6687 20556 6828 20584
rect 6687 20553 6699 20556
rect 6641 20547 6699 20553
rect 6822 20544 6828 20556
rect 6880 20544 6886 20596
rect 9122 20544 9128 20596
rect 9180 20584 9186 20596
rect 9401 20587 9459 20593
rect 9401 20584 9413 20587
rect 9180 20556 9413 20584
rect 9180 20544 9186 20556
rect 9401 20553 9413 20556
rect 9447 20553 9459 20587
rect 9401 20547 9459 20553
rect 9490 20544 9496 20596
rect 9548 20584 9554 20596
rect 9548 20556 14504 20584
rect 9548 20544 9554 20556
rect 1673 20451 1731 20457
rect 1673 20417 1685 20451
rect 1719 20448 1731 20451
rect 1762 20448 1768 20460
rect 1719 20420 1768 20448
rect 1719 20417 1731 20420
rect 1673 20411 1731 20417
rect 1762 20408 1768 20420
rect 1820 20408 1826 20460
rect 2038 20448 2044 20460
rect 1999 20420 2044 20448
rect 2038 20408 2044 20420
rect 2096 20408 2102 20460
rect 2406 20448 2412 20460
rect 2367 20420 2412 20448
rect 2406 20408 2412 20420
rect 2464 20408 2470 20460
rect 2498 20408 2504 20460
rect 2556 20448 2562 20460
rect 2593 20451 2651 20457
rect 2593 20448 2605 20451
rect 2556 20420 2605 20448
rect 2556 20408 2562 20420
rect 2593 20417 2605 20420
rect 2639 20417 2651 20451
rect 2976 20448 3004 20544
rect 8757 20519 8815 20525
rect 8757 20485 8769 20519
rect 8803 20516 8815 20519
rect 8803 20488 11376 20516
rect 8803 20485 8815 20488
rect 8757 20479 8815 20485
rect 3053 20451 3111 20457
rect 3053 20448 3065 20451
rect 2976 20420 3065 20448
rect 2593 20411 2651 20417
rect 3053 20417 3065 20420
rect 3099 20417 3111 20451
rect 3418 20448 3424 20460
rect 3379 20420 3424 20448
rect 3053 20411 3111 20417
rect 3418 20408 3424 20420
rect 3476 20408 3482 20460
rect 3878 20448 3884 20460
rect 3839 20420 3884 20448
rect 3878 20408 3884 20420
rect 3936 20408 3942 20460
rect 4157 20451 4215 20457
rect 4157 20417 4169 20451
rect 4203 20448 4215 20451
rect 4338 20448 4344 20460
rect 4203 20420 4344 20448
rect 4203 20417 4215 20420
rect 4157 20411 4215 20417
rect 4338 20408 4344 20420
rect 4396 20408 4402 20460
rect 4798 20408 4804 20460
rect 4856 20448 4862 20460
rect 5261 20451 5319 20457
rect 5261 20448 5273 20451
rect 4856 20420 5273 20448
rect 4856 20408 4862 20420
rect 5261 20417 5273 20420
rect 5307 20417 5319 20451
rect 5261 20411 5319 20417
rect 5718 20408 5724 20460
rect 5776 20448 5782 20460
rect 6181 20451 6239 20457
rect 6181 20448 6193 20451
rect 5776 20420 6193 20448
rect 5776 20408 5782 20420
rect 6181 20417 6193 20420
rect 6227 20417 6239 20451
rect 6181 20411 6239 20417
rect 6457 20451 6515 20457
rect 6457 20417 6469 20451
rect 6503 20448 6515 20451
rect 7098 20448 7104 20460
rect 6503 20420 7104 20448
rect 6503 20417 6515 20420
rect 6457 20411 6515 20417
rect 7098 20408 7104 20420
rect 7156 20408 7162 20460
rect 7558 20408 7564 20460
rect 7616 20448 7622 20460
rect 7653 20451 7711 20457
rect 7653 20448 7665 20451
rect 7616 20420 7665 20448
rect 7616 20408 7622 20420
rect 7653 20417 7665 20420
rect 7699 20417 7711 20451
rect 7653 20411 7711 20417
rect 8294 20408 8300 20460
rect 8352 20448 8358 20460
rect 8938 20448 8944 20460
rect 8352 20420 8944 20448
rect 8352 20408 8358 20420
rect 8938 20408 8944 20420
rect 8996 20408 9002 20460
rect 9309 20451 9367 20457
rect 9309 20417 9321 20451
rect 9355 20448 9367 20451
rect 9398 20448 9404 20460
rect 9355 20420 9404 20448
rect 9355 20417 9367 20420
rect 9309 20411 9367 20417
rect 9398 20408 9404 20420
rect 9456 20408 9462 20460
rect 9508 20420 10272 20448
rect 2792 20352 4936 20380
rect 2792 20321 2820 20352
rect 2777 20315 2835 20321
rect 2777 20281 2789 20315
rect 2823 20281 2835 20315
rect 2777 20275 2835 20281
rect 3237 20315 3295 20321
rect 3237 20281 3249 20315
rect 3283 20312 3295 20315
rect 4430 20312 4436 20324
rect 3283 20284 4436 20312
rect 3283 20281 3295 20284
rect 3237 20275 3295 20281
rect 4430 20272 4436 20284
rect 4488 20272 4494 20324
rect 4908 20312 4936 20352
rect 4982 20340 4988 20392
rect 5040 20380 5046 20392
rect 5905 20383 5963 20389
rect 5040 20352 5085 20380
rect 5040 20340 5046 20352
rect 5905 20349 5917 20383
rect 5951 20349 5963 20383
rect 5905 20343 5963 20349
rect 5810 20312 5816 20324
rect 4908 20284 5816 20312
rect 5810 20272 5816 20284
rect 5868 20272 5874 20324
rect 5920 20312 5948 20343
rect 6638 20340 6644 20392
rect 6696 20380 6702 20392
rect 6733 20383 6791 20389
rect 6733 20380 6745 20383
rect 6696 20352 6745 20380
rect 6696 20340 6702 20352
rect 6733 20349 6745 20352
rect 6779 20349 6791 20383
rect 7006 20380 7012 20392
rect 6967 20352 7012 20380
rect 6733 20343 6791 20349
rect 7006 20340 7012 20352
rect 7064 20340 7070 20392
rect 7742 20340 7748 20392
rect 7800 20380 7806 20392
rect 7929 20383 7987 20389
rect 7929 20380 7941 20383
rect 7800 20352 7941 20380
rect 7800 20340 7806 20352
rect 7929 20349 7941 20352
rect 7975 20349 7987 20383
rect 9508 20380 9536 20420
rect 10134 20380 10140 20392
rect 7929 20343 7987 20349
rect 8036 20352 9536 20380
rect 10095 20352 10140 20380
rect 5920 20284 6776 20312
rect 6748 20256 6776 20284
rect 7374 20272 7380 20324
rect 7432 20312 7438 20324
rect 8036 20312 8064 20352
rect 10134 20340 10140 20352
rect 10192 20340 10198 20392
rect 7432 20284 8064 20312
rect 9125 20315 9183 20321
rect 7432 20272 7438 20284
rect 9125 20281 9137 20315
rect 9171 20312 9183 20315
rect 9950 20312 9956 20324
rect 9171 20284 9956 20312
rect 9171 20281 9183 20284
rect 9125 20275 9183 20281
rect 9950 20272 9956 20284
rect 10008 20272 10014 20324
rect 10244 20312 10272 20420
rect 10318 20408 10324 20460
rect 10376 20448 10382 20460
rect 11348 20457 11376 20488
rect 12618 20476 12624 20528
rect 12676 20525 12682 20528
rect 12676 20516 12688 20525
rect 12676 20488 12721 20516
rect 12676 20479 12688 20488
rect 12676 20476 12682 20479
rect 12802 20476 12808 20528
rect 12860 20516 12866 20528
rect 12860 20488 14228 20516
rect 12860 20476 12866 20488
rect 10413 20451 10471 20457
rect 10413 20448 10425 20451
rect 10376 20420 10425 20448
rect 10376 20408 10382 20420
rect 10413 20417 10425 20420
rect 10459 20417 10471 20451
rect 10413 20411 10471 20417
rect 11333 20451 11391 20457
rect 11333 20417 11345 20451
rect 11379 20448 11391 20451
rect 11698 20448 11704 20460
rect 11379 20420 11704 20448
rect 11379 20417 11391 20420
rect 11333 20411 11391 20417
rect 11698 20408 11704 20420
rect 11756 20408 11762 20460
rect 12066 20448 12072 20460
rect 11900 20420 12072 20448
rect 11057 20383 11115 20389
rect 11057 20349 11069 20383
rect 11103 20380 11115 20383
rect 11900 20380 11928 20420
rect 12066 20408 12072 20420
rect 12124 20408 12130 20460
rect 14090 20448 14096 20460
rect 14051 20420 14096 20448
rect 14090 20408 14096 20420
rect 14148 20408 14154 20460
rect 12894 20380 12900 20392
rect 11103 20352 11928 20380
rect 12855 20352 12900 20380
rect 11103 20349 11115 20352
rect 11057 20343 11115 20349
rect 12894 20340 12900 20352
rect 12952 20340 12958 20392
rect 13446 20340 13452 20392
rect 13504 20380 13510 20392
rect 13541 20383 13599 20389
rect 13541 20380 13553 20383
rect 13504 20352 13553 20380
rect 13504 20340 13510 20352
rect 13541 20349 13553 20352
rect 13587 20349 13599 20383
rect 13541 20343 13599 20349
rect 13817 20383 13875 20389
rect 13817 20349 13829 20383
rect 13863 20380 13875 20383
rect 13906 20380 13912 20392
rect 13863 20352 13912 20380
rect 13863 20349 13875 20352
rect 13817 20343 13875 20349
rect 11882 20312 11888 20324
rect 10244 20284 11888 20312
rect 11882 20272 11888 20284
rect 11940 20272 11946 20324
rect 13832 20312 13860 20343
rect 13906 20340 13912 20352
rect 13964 20340 13970 20392
rect 14200 20380 14228 20488
rect 14476 20457 14504 20556
rect 14550 20544 14556 20596
rect 14608 20584 14614 20596
rect 15013 20587 15071 20593
rect 15013 20584 15025 20587
rect 14608 20556 15025 20584
rect 14608 20544 14614 20556
rect 15013 20553 15025 20556
rect 15059 20553 15071 20587
rect 15013 20547 15071 20553
rect 15378 20544 15384 20596
rect 15436 20584 15442 20596
rect 15749 20587 15807 20593
rect 15749 20584 15761 20587
rect 15436 20556 15761 20584
rect 15436 20544 15442 20556
rect 15749 20553 15761 20556
rect 15795 20553 15807 20587
rect 15749 20547 15807 20553
rect 15838 20544 15844 20596
rect 15896 20584 15902 20596
rect 16117 20587 16175 20593
rect 16117 20584 16129 20587
rect 15896 20556 16129 20584
rect 15896 20544 15902 20556
rect 16117 20553 16129 20556
rect 16163 20553 16175 20587
rect 16117 20547 16175 20553
rect 16298 20544 16304 20596
rect 16356 20584 16362 20596
rect 16853 20587 16911 20593
rect 16853 20584 16865 20587
rect 16356 20556 16865 20584
rect 16356 20544 16362 20556
rect 16853 20553 16865 20556
rect 16899 20553 16911 20587
rect 16853 20547 16911 20553
rect 17218 20544 17224 20596
rect 17276 20584 17282 20596
rect 17589 20587 17647 20593
rect 17589 20584 17601 20587
rect 17276 20556 17601 20584
rect 17276 20544 17282 20556
rect 17589 20553 17601 20556
rect 17635 20553 17647 20587
rect 17954 20584 17960 20596
rect 17915 20556 17960 20584
rect 17589 20547 17647 20553
rect 17954 20544 17960 20556
rect 18012 20544 18018 20596
rect 18138 20544 18144 20596
rect 18196 20584 18202 20596
rect 18417 20587 18475 20593
rect 18417 20584 18429 20587
rect 18196 20556 18429 20584
rect 18196 20544 18202 20556
rect 18417 20553 18429 20556
rect 18463 20553 18475 20587
rect 18417 20547 18475 20553
rect 18598 20544 18604 20596
rect 18656 20584 18662 20596
rect 18877 20587 18935 20593
rect 18877 20584 18889 20587
rect 18656 20556 18889 20584
rect 18656 20544 18662 20556
rect 18877 20553 18889 20556
rect 18923 20553 18935 20587
rect 18877 20547 18935 20553
rect 14642 20476 14648 20528
rect 14700 20516 14706 20528
rect 19429 20519 19487 20525
rect 14700 20488 15976 20516
rect 14700 20476 14706 20488
rect 14461 20451 14519 20457
rect 14461 20417 14473 20451
rect 14507 20417 14519 20451
rect 14461 20411 14519 20417
rect 14550 20408 14556 20460
rect 14608 20448 14614 20460
rect 14829 20451 14887 20457
rect 14829 20448 14841 20451
rect 14608 20420 14841 20448
rect 14608 20408 14614 20420
rect 14829 20417 14841 20420
rect 14875 20417 14887 20451
rect 15194 20448 15200 20460
rect 15155 20420 15200 20448
rect 14829 20411 14887 20417
rect 15194 20408 15200 20420
rect 15252 20408 15258 20460
rect 15948 20457 15976 20488
rect 19429 20485 19441 20519
rect 19475 20516 19487 20519
rect 22738 20516 22744 20528
rect 19475 20488 22744 20516
rect 19475 20485 19487 20488
rect 19429 20479 19487 20485
rect 15565 20451 15623 20457
rect 15565 20417 15577 20451
rect 15611 20417 15623 20451
rect 15565 20411 15623 20417
rect 15933 20451 15991 20457
rect 15933 20417 15945 20451
rect 15979 20417 15991 20451
rect 15933 20411 15991 20417
rect 15580 20380 15608 20411
rect 16022 20408 16028 20460
rect 16080 20448 16086 20460
rect 16669 20451 16727 20457
rect 16669 20448 16681 20451
rect 16080 20420 16681 20448
rect 16080 20408 16086 20420
rect 16669 20417 16681 20420
rect 16715 20417 16727 20451
rect 17034 20448 17040 20460
rect 16995 20420 17040 20448
rect 16669 20411 16727 20417
rect 17034 20408 17040 20420
rect 17092 20408 17098 20460
rect 17126 20408 17132 20460
rect 17184 20448 17190 20460
rect 17405 20451 17463 20457
rect 17405 20448 17417 20451
rect 17184 20420 17417 20448
rect 17184 20408 17190 20420
rect 17405 20417 17417 20420
rect 17451 20417 17463 20451
rect 17770 20448 17776 20460
rect 17731 20420 17776 20448
rect 17405 20411 17463 20417
rect 17770 20408 17776 20420
rect 17828 20408 17834 20460
rect 18230 20448 18236 20460
rect 18191 20420 18236 20448
rect 18230 20408 18236 20420
rect 18288 20408 18294 20460
rect 18690 20448 18696 20460
rect 18651 20420 18696 20448
rect 18690 20408 18696 20420
rect 18748 20408 18754 20460
rect 19536 20457 19564 20488
rect 22738 20476 22744 20488
rect 22796 20476 22802 20528
rect 19521 20451 19579 20457
rect 19521 20417 19533 20451
rect 19567 20417 19579 20451
rect 19521 20411 19579 20417
rect 19610 20408 19616 20460
rect 19668 20448 19674 20460
rect 20625 20451 20683 20457
rect 20625 20448 20637 20451
rect 19668 20420 20637 20448
rect 19668 20408 19674 20420
rect 20625 20417 20637 20420
rect 20671 20448 20683 20451
rect 22278 20448 22284 20460
rect 20671 20420 22284 20448
rect 20671 20417 20683 20420
rect 20625 20411 20683 20417
rect 22278 20408 22284 20420
rect 22336 20408 22342 20460
rect 14200 20352 15608 20380
rect 18322 20340 18328 20392
rect 18380 20380 18386 20392
rect 19797 20383 19855 20389
rect 19797 20380 19809 20383
rect 18380 20352 19809 20380
rect 18380 20340 18386 20352
rect 19797 20349 19809 20352
rect 19843 20349 19855 20383
rect 20806 20380 20812 20392
rect 20767 20352 20812 20380
rect 19797 20343 19855 20349
rect 20806 20340 20812 20352
rect 20864 20340 20870 20392
rect 13740 20284 13860 20312
rect 13740 20256 13768 20284
rect 13998 20272 14004 20324
rect 14056 20312 14062 20324
rect 14645 20315 14703 20321
rect 14645 20312 14657 20315
rect 14056 20284 14657 20312
rect 14056 20272 14062 20284
rect 14645 20281 14657 20284
rect 14691 20281 14703 20315
rect 14645 20275 14703 20281
rect 14918 20272 14924 20324
rect 14976 20312 14982 20324
rect 15381 20315 15439 20321
rect 15381 20312 15393 20315
rect 14976 20284 15393 20312
rect 14976 20272 14982 20284
rect 15381 20281 15393 20284
rect 15427 20281 15439 20315
rect 15381 20275 15439 20281
rect 16942 20272 16948 20324
rect 17000 20312 17006 20324
rect 17221 20315 17279 20321
rect 17221 20312 17233 20315
rect 17000 20284 17233 20312
rect 17000 20272 17006 20284
rect 17221 20281 17233 20284
rect 17267 20281 17279 20315
rect 17221 20275 17279 20281
rect 1486 20244 1492 20256
rect 1447 20216 1492 20244
rect 1486 20204 1492 20216
rect 1544 20204 1550 20256
rect 3970 20204 3976 20256
rect 4028 20244 4034 20256
rect 4065 20247 4123 20253
rect 4065 20244 4077 20247
rect 4028 20216 4077 20244
rect 4028 20204 4034 20216
rect 4065 20213 4077 20216
rect 4111 20213 4123 20247
rect 4065 20207 4123 20213
rect 4341 20247 4399 20253
rect 4341 20213 4353 20247
rect 4387 20244 4399 20247
rect 5902 20244 5908 20256
rect 4387 20216 5908 20244
rect 4387 20213 4399 20216
rect 4341 20207 4399 20213
rect 5902 20204 5908 20216
rect 5960 20204 5966 20256
rect 6730 20204 6736 20256
rect 6788 20204 6794 20256
rect 11054 20204 11060 20256
rect 11112 20244 11118 20256
rect 11517 20247 11575 20253
rect 11517 20244 11529 20247
rect 11112 20216 11529 20244
rect 11112 20204 11118 20216
rect 11517 20213 11529 20216
rect 11563 20213 11575 20247
rect 11517 20207 11575 20213
rect 13722 20204 13728 20256
rect 13780 20204 13786 20256
rect 13814 20204 13820 20256
rect 13872 20244 13878 20256
rect 14277 20247 14335 20253
rect 14277 20244 14289 20247
rect 13872 20216 14289 20244
rect 13872 20204 13878 20216
rect 14277 20213 14289 20216
rect 14323 20213 14335 20247
rect 14277 20207 14335 20213
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 2406 20000 2412 20052
rect 2464 20040 2470 20052
rect 2685 20043 2743 20049
rect 2685 20040 2697 20043
rect 2464 20012 2697 20040
rect 2464 20000 2470 20012
rect 2685 20009 2697 20012
rect 2731 20009 2743 20043
rect 2685 20003 2743 20009
rect 3418 20000 3424 20052
rect 3476 20040 3482 20052
rect 3789 20043 3847 20049
rect 3789 20040 3801 20043
rect 3476 20012 3801 20040
rect 3476 20000 3482 20012
rect 3789 20009 3801 20012
rect 3835 20009 3847 20043
rect 3789 20003 3847 20009
rect 3878 20000 3884 20052
rect 3936 20040 3942 20052
rect 4157 20043 4215 20049
rect 4157 20040 4169 20043
rect 3936 20012 4169 20040
rect 3936 20000 3942 20012
rect 4157 20009 4169 20012
rect 4203 20009 4215 20043
rect 4157 20003 4215 20009
rect 4338 20000 4344 20052
rect 4396 20040 4402 20052
rect 4433 20043 4491 20049
rect 4433 20040 4445 20043
rect 4396 20012 4445 20040
rect 4396 20000 4402 20012
rect 4433 20009 4445 20012
rect 4479 20009 4491 20043
rect 4433 20003 4491 20009
rect 4798 20000 4804 20052
rect 4856 20040 4862 20052
rect 4985 20043 5043 20049
rect 4985 20040 4997 20043
rect 4856 20012 4997 20040
rect 4856 20000 4862 20012
rect 4985 20009 4997 20012
rect 5031 20009 5043 20043
rect 5258 20040 5264 20052
rect 5219 20012 5264 20040
rect 4985 20003 5043 20009
rect 5258 20000 5264 20012
rect 5316 20000 5322 20052
rect 5994 20040 6000 20052
rect 5955 20012 6000 20040
rect 5994 20000 6000 20012
rect 6052 20000 6058 20052
rect 6181 20043 6239 20049
rect 6181 20009 6193 20043
rect 6227 20040 6239 20043
rect 7098 20040 7104 20052
rect 6227 20012 7104 20040
rect 6227 20009 6239 20012
rect 6181 20003 6239 20009
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 7466 20040 7472 20052
rect 7427 20012 7472 20040
rect 7466 20000 7472 20012
rect 7524 20000 7530 20052
rect 8757 20043 8815 20049
rect 8757 20009 8769 20043
rect 8803 20040 8815 20043
rect 9214 20040 9220 20052
rect 8803 20012 9220 20040
rect 8803 20009 8815 20012
rect 8757 20003 8815 20009
rect 9214 20000 9220 20012
rect 9272 20000 9278 20052
rect 9585 20043 9643 20049
rect 9585 20009 9597 20043
rect 9631 20040 9643 20043
rect 11790 20040 11796 20052
rect 9631 20012 11796 20040
rect 9631 20009 9643 20012
rect 9585 20003 9643 20009
rect 11790 20000 11796 20012
rect 11848 20000 11854 20052
rect 11882 20000 11888 20052
rect 11940 20040 11946 20052
rect 12894 20040 12900 20052
rect 11940 20012 12900 20040
rect 11940 20000 11946 20012
rect 12894 20000 12900 20012
rect 12952 20040 12958 20052
rect 12989 20043 13047 20049
rect 12989 20040 13001 20043
rect 12952 20012 13001 20040
rect 12952 20000 12958 20012
rect 12989 20009 13001 20012
rect 13035 20009 13047 20043
rect 12989 20003 13047 20009
rect 13078 20000 13084 20052
rect 13136 20040 13142 20052
rect 13357 20043 13415 20049
rect 13357 20040 13369 20043
rect 13136 20012 13369 20040
rect 13136 20000 13142 20012
rect 13357 20009 13369 20012
rect 13403 20009 13415 20043
rect 13357 20003 13415 20009
rect 13722 20000 13728 20052
rect 13780 20040 13786 20052
rect 13817 20043 13875 20049
rect 13817 20040 13829 20043
rect 13780 20012 13829 20040
rect 13780 20000 13786 20012
rect 13817 20009 13829 20012
rect 13863 20009 13875 20043
rect 17770 20040 17776 20052
rect 13817 20003 13875 20009
rect 13924 20012 17776 20040
rect 2130 19932 2136 19984
rect 2188 19972 2194 19984
rect 3145 19975 3203 19981
rect 3145 19972 3157 19975
rect 2188 19944 3157 19972
rect 2188 19932 2194 19944
rect 3145 19941 3157 19944
rect 3191 19941 3203 19975
rect 3145 19935 3203 19941
rect 2590 19904 2596 19916
rect 2056 19876 2596 19904
rect 1670 19836 1676 19848
rect 1631 19808 1676 19836
rect 1670 19796 1676 19808
rect 1728 19796 1734 19848
rect 2056 19845 2084 19876
rect 2590 19864 2596 19876
rect 2648 19864 2654 19916
rect 2961 19907 3019 19913
rect 2961 19904 2973 19907
rect 2700 19876 2973 19904
rect 2041 19839 2099 19845
rect 2041 19805 2053 19839
rect 2087 19805 2099 19839
rect 2041 19799 2099 19805
rect 2130 19796 2136 19848
rect 2188 19836 2194 19848
rect 2409 19839 2467 19845
rect 2188 19808 2233 19836
rect 2188 19796 2194 19808
rect 2409 19805 2421 19839
rect 2455 19836 2467 19839
rect 2700 19836 2728 19876
rect 2961 19873 2973 19876
rect 3007 19873 3019 19907
rect 6012 19904 6040 20000
rect 7745 19975 7803 19981
rect 7745 19941 7757 19975
rect 7791 19972 7803 19975
rect 7791 19944 11560 19972
rect 7791 19941 7803 19944
rect 7745 19935 7803 19941
rect 6273 19907 6331 19913
rect 6273 19904 6285 19907
rect 6012 19876 6285 19904
rect 2961 19867 3019 19873
rect 6273 19873 6285 19876
rect 6319 19873 6331 19907
rect 6273 19867 6331 19873
rect 9858 19864 9864 19916
rect 9916 19904 9922 19916
rect 10505 19907 10563 19913
rect 10505 19904 10517 19907
rect 9916 19876 10517 19904
rect 9916 19864 9922 19876
rect 10505 19873 10517 19876
rect 10551 19904 10563 19907
rect 10686 19904 10692 19916
rect 10551 19876 10692 19904
rect 10551 19873 10563 19876
rect 10505 19867 10563 19873
rect 10686 19864 10692 19876
rect 10744 19864 10750 19916
rect 11238 19864 11244 19916
rect 11296 19904 11302 19916
rect 11425 19907 11483 19913
rect 11425 19904 11437 19907
rect 11296 19876 11437 19904
rect 11296 19864 11302 19876
rect 11425 19873 11437 19876
rect 11471 19873 11483 19907
rect 11425 19867 11483 19873
rect 2455 19808 2728 19836
rect 2869 19839 2927 19845
rect 2455 19805 2467 19808
rect 2409 19799 2467 19805
rect 2869 19805 2881 19839
rect 2915 19805 2927 19839
rect 2869 19799 2927 19805
rect 1578 19728 1584 19780
rect 1636 19768 1642 19780
rect 2424 19768 2452 19799
rect 1636 19740 2452 19768
rect 2884 19768 2912 19799
rect 5258 19796 5264 19848
rect 5316 19836 5322 19848
rect 5353 19839 5411 19845
rect 5353 19836 5365 19839
rect 5316 19808 5365 19836
rect 5316 19796 5322 19808
rect 5353 19805 5365 19808
rect 5399 19805 5411 19839
rect 6546 19836 6552 19848
rect 6507 19808 6552 19836
rect 5353 19799 5411 19805
rect 6546 19796 6552 19808
rect 6604 19796 6610 19848
rect 7098 19796 7104 19848
rect 7156 19836 7162 19848
rect 7285 19839 7343 19845
rect 7285 19836 7297 19839
rect 7156 19808 7297 19836
rect 7156 19796 7162 19808
rect 7285 19805 7297 19808
rect 7331 19805 7343 19839
rect 7285 19799 7343 19805
rect 7561 19839 7619 19845
rect 7561 19805 7573 19839
rect 7607 19836 7619 19839
rect 7650 19836 7656 19848
rect 7607 19808 7656 19836
rect 7607 19805 7619 19808
rect 7561 19799 7619 19805
rect 7650 19796 7656 19808
rect 7708 19796 7714 19848
rect 8018 19836 8024 19848
rect 7979 19808 8024 19836
rect 8018 19796 8024 19808
rect 8076 19796 8082 19848
rect 8110 19796 8116 19848
rect 8168 19836 8174 19848
rect 8205 19839 8263 19845
rect 8205 19836 8217 19839
rect 8168 19808 8217 19836
rect 8168 19796 8174 19808
rect 8205 19805 8217 19808
rect 8251 19805 8263 19839
rect 8205 19799 8263 19805
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19836 8631 19839
rect 8662 19836 8668 19848
rect 8619 19808 8668 19836
rect 8619 19805 8631 19808
rect 8573 19799 8631 19805
rect 8662 19796 8668 19808
rect 8720 19796 8726 19848
rect 9398 19836 9404 19848
rect 9359 19808 9404 19836
rect 9398 19796 9404 19808
rect 9456 19796 9462 19848
rect 10226 19836 10232 19848
rect 10187 19808 10232 19836
rect 10226 19796 10232 19808
rect 10284 19796 10290 19848
rect 11146 19836 11152 19848
rect 11107 19808 11152 19836
rect 11146 19796 11152 19808
rect 11204 19796 11210 19848
rect 11532 19836 11560 19944
rect 13446 19932 13452 19984
rect 13504 19972 13510 19984
rect 13924 19972 13952 20012
rect 17770 20000 17776 20012
rect 17828 20000 17834 20052
rect 18693 20043 18751 20049
rect 18693 20009 18705 20043
rect 18739 20040 18751 20043
rect 19610 20040 19616 20052
rect 18739 20012 19616 20040
rect 18739 20009 18751 20012
rect 18693 20003 18751 20009
rect 19610 20000 19616 20012
rect 19668 20000 19674 20052
rect 21358 20040 21364 20052
rect 20640 20012 21364 20040
rect 13504 19944 13952 19972
rect 14277 19975 14335 19981
rect 13504 19932 13510 19944
rect 14277 19941 14289 19975
rect 14323 19941 14335 19975
rect 14277 19935 14335 19941
rect 14553 19975 14611 19981
rect 14553 19941 14565 19975
rect 14599 19972 14611 19975
rect 18969 19975 19027 19981
rect 14599 19944 18920 19972
rect 14599 19941 14611 19944
rect 14553 19935 14611 19941
rect 12986 19864 12992 19916
rect 13044 19904 13050 19916
rect 13538 19904 13544 19916
rect 13044 19876 13544 19904
rect 13044 19864 13050 19876
rect 13538 19864 13544 19876
rect 13596 19904 13602 19916
rect 14292 19904 14320 19935
rect 13596 19876 13768 19904
rect 14292 19876 18828 19904
rect 13596 19864 13602 19876
rect 11532 19808 12839 19836
rect 5813 19771 5871 19777
rect 2884 19740 5672 19768
rect 1636 19728 1642 19740
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 1854 19700 1860 19712
rect 1815 19672 1860 19700
rect 1854 19660 1860 19672
rect 1912 19660 1918 19712
rect 2314 19700 2320 19712
rect 2275 19672 2320 19700
rect 2314 19660 2320 19672
rect 2372 19660 2378 19712
rect 2593 19703 2651 19709
rect 2593 19669 2605 19703
rect 2639 19700 2651 19703
rect 2682 19700 2688 19712
rect 2639 19672 2688 19700
rect 2639 19669 2651 19672
rect 2593 19663 2651 19669
rect 2682 19660 2688 19672
rect 2740 19660 2746 19712
rect 5534 19700 5540 19712
rect 5495 19672 5540 19700
rect 5534 19660 5540 19672
rect 5592 19660 5598 19712
rect 5644 19700 5672 19740
rect 5813 19737 5825 19771
rect 5859 19768 5871 19771
rect 6638 19768 6644 19780
rect 5859 19740 6644 19768
rect 5859 19737 5871 19740
rect 5813 19731 5871 19737
rect 6638 19728 6644 19740
rect 6696 19728 6702 19780
rect 6748 19740 7880 19768
rect 6748 19700 6776 19740
rect 7852 19709 7880 19740
rect 8478 19728 8484 19780
rect 8536 19768 8542 19780
rect 9033 19771 9091 19777
rect 9033 19768 9045 19771
rect 8536 19740 9045 19768
rect 8536 19728 8542 19740
rect 9033 19737 9045 19740
rect 9079 19737 9091 19771
rect 9214 19768 9220 19780
rect 9175 19740 9220 19768
rect 9033 19731 9091 19737
rect 9214 19728 9220 19740
rect 9272 19728 9278 19780
rect 10042 19728 10048 19780
rect 10100 19768 10106 19780
rect 10100 19740 12434 19768
rect 10100 19728 10106 19740
rect 5644 19672 6776 19700
rect 7837 19703 7895 19709
rect 7837 19669 7849 19703
rect 7883 19669 7895 19703
rect 7837 19663 7895 19669
rect 8297 19703 8355 19709
rect 8297 19669 8309 19703
rect 8343 19700 8355 19703
rect 10594 19700 10600 19712
rect 8343 19672 10600 19700
rect 8343 19669 8355 19672
rect 8297 19663 8355 19669
rect 10594 19660 10600 19672
rect 10652 19660 10658 19712
rect 11517 19703 11575 19709
rect 11517 19669 11529 19703
rect 11563 19700 11575 19703
rect 11790 19700 11796 19712
rect 11563 19672 11796 19700
rect 11563 19669 11575 19672
rect 11517 19663 11575 19669
rect 11790 19660 11796 19672
rect 11848 19660 11854 19712
rect 12406 19700 12434 19740
rect 12618 19728 12624 19780
rect 12676 19777 12682 19780
rect 12676 19768 12688 19777
rect 12811 19768 12839 19808
rect 12894 19796 12900 19848
rect 12952 19836 12958 19848
rect 13170 19836 13176 19848
rect 12952 19808 12997 19836
rect 13131 19808 13176 19836
rect 12952 19796 12958 19808
rect 13170 19796 13176 19808
rect 13228 19796 13234 19848
rect 13740 19845 13768 19876
rect 13725 19839 13783 19845
rect 13725 19805 13737 19839
rect 13771 19805 13783 19839
rect 14090 19836 14096 19848
rect 14051 19808 14096 19836
rect 13725 19799 13783 19805
rect 14090 19796 14096 19808
rect 14148 19796 14154 19848
rect 14369 19839 14427 19845
rect 14369 19805 14381 19839
rect 14415 19836 14427 19839
rect 14458 19836 14464 19848
rect 14415 19808 14464 19836
rect 14415 19805 14427 19808
rect 14369 19799 14427 19805
rect 14458 19796 14464 19808
rect 14516 19836 14522 19848
rect 18800 19845 18828 19876
rect 14829 19839 14887 19845
rect 14829 19836 14841 19839
rect 14516 19808 14841 19836
rect 14516 19796 14522 19808
rect 14829 19805 14841 19808
rect 14875 19805 14887 19839
rect 14829 19799 14887 19805
rect 16301 19839 16359 19845
rect 16301 19805 16313 19839
rect 16347 19805 16359 19839
rect 16301 19799 16359 19805
rect 18785 19839 18843 19845
rect 18785 19805 18797 19839
rect 18831 19805 18843 19839
rect 18892 19836 18920 19944
rect 18969 19941 18981 19975
rect 19015 19941 19027 19975
rect 18969 19935 19027 19941
rect 18984 19904 19012 19935
rect 19058 19932 19064 19984
rect 19116 19972 19122 19984
rect 19429 19975 19487 19981
rect 19429 19972 19441 19975
rect 19116 19944 19441 19972
rect 19116 19932 19122 19944
rect 19429 19941 19441 19944
rect 19475 19941 19487 19975
rect 19429 19935 19487 19941
rect 19518 19932 19524 19984
rect 19576 19972 19582 19984
rect 19797 19975 19855 19981
rect 19797 19972 19809 19975
rect 19576 19944 19809 19972
rect 19576 19932 19582 19944
rect 19797 19941 19809 19944
rect 19843 19941 19855 19975
rect 20640 19972 20668 20012
rect 21358 20000 21364 20012
rect 21416 20000 21422 20052
rect 19797 19935 19855 19941
rect 20180 19944 20668 19972
rect 20180 19904 20208 19944
rect 18984 19876 20208 19904
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 18892 19808 19257 19836
rect 18785 19799 18843 19805
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 14550 19768 14556 19780
rect 12676 19740 12721 19768
rect 12811 19740 14556 19768
rect 12676 19731 12688 19740
rect 12676 19728 12682 19731
rect 14550 19728 14556 19740
rect 14608 19728 14614 19780
rect 16316 19712 16344 19799
rect 19518 19796 19524 19848
rect 19576 19836 19582 19848
rect 19613 19839 19671 19845
rect 19613 19836 19625 19839
rect 19576 19808 19625 19836
rect 19576 19796 19582 19808
rect 19613 19805 19625 19808
rect 19659 19805 19671 19839
rect 21545 19839 21603 19845
rect 21545 19836 21557 19839
rect 19613 19799 19671 19805
rect 20824 19808 21557 19836
rect 20824 19780 20852 19808
rect 21545 19805 21557 19808
rect 21591 19805 21603 19839
rect 21545 19799 21603 19805
rect 20806 19768 20812 19780
rect 19996 19740 20812 19768
rect 19996 19712 20024 19740
rect 20806 19728 20812 19740
rect 20864 19728 20870 19780
rect 21266 19728 21272 19780
rect 21324 19777 21330 19780
rect 21324 19768 21336 19777
rect 21324 19740 21369 19768
rect 21324 19731 21336 19740
rect 21324 19728 21330 19731
rect 13446 19700 13452 19712
rect 12406 19672 13452 19700
rect 13446 19660 13452 19672
rect 13504 19660 13510 19712
rect 13541 19703 13599 19709
rect 13541 19669 13553 19703
rect 13587 19700 13599 19703
rect 13630 19700 13636 19712
rect 13587 19672 13636 19700
rect 13587 19669 13599 19672
rect 13541 19663 13599 19669
rect 13630 19660 13636 19672
rect 13688 19660 13694 19712
rect 14090 19660 14096 19712
rect 14148 19700 14154 19712
rect 14645 19703 14703 19709
rect 14645 19700 14657 19703
rect 14148 19672 14657 19700
rect 14148 19660 14154 19672
rect 14645 19669 14657 19672
rect 14691 19700 14703 19703
rect 14826 19700 14832 19712
rect 14691 19672 14832 19700
rect 14691 19669 14703 19672
rect 14645 19663 14703 19669
rect 14826 19660 14832 19672
rect 14884 19660 14890 19712
rect 16209 19703 16267 19709
rect 16209 19669 16221 19703
rect 16255 19700 16267 19703
rect 16298 19700 16304 19712
rect 16255 19672 16304 19700
rect 16255 19669 16267 19672
rect 16209 19663 16267 19669
rect 16298 19660 16304 19672
rect 16356 19660 16362 19712
rect 16485 19703 16543 19709
rect 16485 19669 16497 19703
rect 16531 19700 16543 19703
rect 19610 19700 19616 19712
rect 16531 19672 19616 19700
rect 16531 19669 16543 19672
rect 16485 19663 16543 19669
rect 19610 19660 19616 19672
rect 19668 19660 19674 19712
rect 19978 19700 19984 19712
rect 19939 19672 19984 19700
rect 19978 19660 19984 19672
rect 20036 19660 20042 19712
rect 20162 19700 20168 19712
rect 20123 19672 20168 19700
rect 20162 19660 20168 19672
rect 20220 19660 20226 19712
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 2498 19456 2504 19508
rect 2556 19496 2562 19508
rect 2685 19499 2743 19505
rect 2685 19496 2697 19499
rect 2556 19468 2697 19496
rect 2556 19456 2562 19468
rect 2685 19465 2697 19468
rect 2731 19465 2743 19499
rect 2685 19459 2743 19465
rect 5718 19456 5724 19508
rect 5776 19496 5782 19508
rect 6365 19499 6423 19505
rect 6365 19496 6377 19499
rect 5776 19468 6377 19496
rect 5776 19456 5782 19468
rect 6365 19465 6377 19468
rect 6411 19465 6423 19499
rect 6365 19459 6423 19465
rect 7101 19499 7159 19505
rect 7101 19465 7113 19499
rect 7147 19496 7159 19499
rect 8110 19496 8116 19508
rect 7147 19468 8116 19496
rect 7147 19465 7159 19468
rect 7101 19459 7159 19465
rect 8110 19456 8116 19468
rect 8168 19456 8174 19508
rect 8297 19499 8355 19505
rect 8297 19465 8309 19499
rect 8343 19496 8355 19499
rect 9582 19496 9588 19508
rect 8343 19468 9588 19496
rect 8343 19465 8355 19468
rect 8297 19459 8355 19465
rect 9582 19456 9588 19468
rect 9640 19456 9646 19508
rect 9766 19496 9772 19508
rect 9727 19468 9772 19496
rect 9766 19456 9772 19468
rect 9824 19456 9830 19508
rect 10042 19496 10048 19508
rect 10003 19468 10048 19496
rect 10042 19456 10048 19468
rect 10100 19456 10106 19508
rect 10689 19499 10747 19505
rect 10689 19465 10701 19499
rect 10735 19465 10747 19499
rect 11238 19496 11244 19508
rect 11199 19468 11244 19496
rect 10689 19459 10747 19465
rect 9674 19428 9680 19440
rect 1688 19400 2728 19428
rect 1688 19369 1716 19400
rect 2700 19372 2728 19400
rect 9324 19400 9680 19428
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19329 1731 19363
rect 1673 19323 1731 19329
rect 1765 19363 1823 19369
rect 1765 19329 1777 19363
rect 1811 19360 1823 19363
rect 1854 19360 1860 19372
rect 1811 19332 1860 19360
rect 1811 19329 1823 19332
rect 1765 19323 1823 19329
rect 1854 19320 1860 19332
rect 1912 19320 1918 19372
rect 2041 19363 2099 19369
rect 2041 19329 2053 19363
rect 2087 19360 2099 19363
rect 2317 19363 2375 19369
rect 2317 19360 2329 19363
rect 2087 19332 2329 19360
rect 2087 19329 2099 19332
rect 2041 19323 2099 19329
rect 2317 19329 2329 19332
rect 2363 19329 2375 19363
rect 2317 19323 2375 19329
rect 198 19252 204 19304
rect 256 19292 262 19304
rect 2056 19292 2084 19323
rect 2682 19320 2688 19372
rect 2740 19320 2746 19372
rect 5994 19360 6000 19372
rect 2792 19332 6000 19360
rect 2792 19292 2820 19332
rect 5994 19320 6000 19332
rect 6052 19320 6058 19372
rect 7193 19363 7251 19369
rect 7193 19360 7205 19363
rect 6932 19332 7205 19360
rect 256 19264 2084 19292
rect 2746 19264 2820 19292
rect 256 19252 262 19264
rect 1118 19184 1124 19236
rect 1176 19224 1182 19236
rect 1854 19224 1860 19236
rect 1176 19196 1860 19224
rect 1176 19184 1182 19196
rect 1854 19184 1860 19196
rect 1912 19224 1918 19236
rect 2501 19227 2559 19233
rect 2501 19224 2513 19227
rect 1912 19196 2513 19224
rect 1912 19184 1918 19196
rect 2501 19193 2513 19196
rect 2547 19193 2559 19227
rect 2501 19187 2559 19193
rect 1486 19156 1492 19168
rect 1447 19128 1492 19156
rect 1486 19116 1492 19128
rect 1544 19116 1550 19168
rect 2225 19159 2283 19165
rect 2225 19125 2237 19159
rect 2271 19156 2283 19159
rect 2746 19156 2774 19264
rect 5534 19184 5540 19236
rect 5592 19224 5598 19236
rect 6932 19233 6960 19332
rect 7193 19329 7205 19332
rect 7239 19329 7251 19363
rect 8113 19363 8171 19369
rect 8113 19360 8125 19363
rect 7193 19323 7251 19329
rect 7576 19332 8125 19360
rect 6917 19227 6975 19233
rect 6917 19224 6929 19227
rect 5592 19196 6929 19224
rect 5592 19184 5598 19196
rect 6917 19193 6929 19196
rect 6963 19193 6975 19227
rect 6917 19187 6975 19193
rect 7190 19184 7196 19236
rect 7248 19224 7254 19236
rect 7576 19224 7604 19332
rect 8113 19329 8125 19332
rect 8159 19329 8171 19363
rect 8386 19360 8392 19372
rect 8347 19332 8392 19360
rect 8113 19323 8171 19329
rect 8386 19320 8392 19332
rect 8444 19320 8450 19372
rect 8938 19320 8944 19372
rect 8996 19360 9002 19372
rect 9324 19369 9352 19400
rect 9674 19388 9680 19400
rect 9732 19388 9738 19440
rect 10410 19428 10416 19440
rect 9876 19400 10416 19428
rect 9033 19363 9091 19369
rect 9033 19360 9045 19363
rect 8996 19332 9045 19360
rect 8996 19320 9002 19332
rect 9033 19329 9045 19332
rect 9079 19329 9091 19363
rect 9033 19323 9091 19329
rect 9309 19363 9367 19369
rect 9309 19329 9321 19363
rect 9355 19329 9367 19363
rect 9582 19360 9588 19372
rect 9543 19332 9588 19360
rect 9309 19323 9367 19329
rect 9582 19320 9588 19332
rect 9640 19320 9646 19372
rect 9876 19369 9904 19400
rect 10410 19388 10416 19400
rect 10468 19388 10474 19440
rect 10704 19428 10732 19459
rect 11238 19456 11244 19468
rect 11296 19456 11302 19508
rect 12434 19496 12440 19508
rect 11348 19468 12440 19496
rect 11348 19428 11376 19468
rect 12434 19456 12440 19468
rect 12492 19456 12498 19508
rect 20070 19456 20076 19508
rect 20128 19496 20134 19508
rect 20993 19499 21051 19505
rect 20993 19496 21005 19499
rect 20128 19468 21005 19496
rect 20128 19456 20134 19468
rect 20993 19465 21005 19468
rect 21039 19465 21051 19499
rect 20993 19459 21051 19465
rect 21361 19499 21419 19505
rect 21361 19465 21373 19499
rect 21407 19465 21419 19499
rect 21361 19459 21419 19465
rect 18230 19428 18236 19440
rect 10704 19400 11376 19428
rect 11624 19400 18236 19428
rect 9861 19363 9919 19369
rect 9861 19360 9873 19363
rect 9784 19332 9873 19360
rect 7653 19295 7711 19301
rect 7653 19261 7665 19295
rect 7699 19292 7711 19295
rect 8294 19292 8300 19304
rect 7699 19264 8300 19292
rect 7699 19261 7711 19264
rect 7653 19255 7711 19261
rect 8294 19252 8300 19264
rect 8352 19252 8358 19304
rect 8849 19295 8907 19301
rect 8849 19261 8861 19295
rect 8895 19292 8907 19295
rect 9784 19292 9812 19332
rect 9861 19329 9873 19332
rect 9907 19329 9919 19363
rect 9861 19323 9919 19329
rect 10134 19320 10140 19372
rect 10192 19360 10198 19372
rect 10229 19363 10287 19369
rect 10229 19360 10241 19363
rect 10192 19332 10241 19360
rect 10192 19320 10198 19332
rect 10229 19329 10241 19332
rect 10275 19329 10287 19363
rect 10229 19323 10287 19329
rect 10505 19363 10563 19369
rect 10505 19329 10517 19363
rect 10551 19329 10563 19363
rect 10505 19323 10563 19329
rect 11057 19363 11115 19369
rect 11057 19329 11069 19363
rect 11103 19329 11115 19363
rect 11624 19360 11652 19400
rect 18230 19388 18236 19400
rect 18288 19388 18294 19440
rect 19978 19428 19984 19440
rect 19352 19400 19984 19428
rect 11057 19323 11115 19329
rect 11164 19332 11652 19360
rect 10520 19292 10548 19323
rect 8895 19264 9812 19292
rect 9876 19264 10548 19292
rect 8895 19261 8907 19264
rect 8849 19255 8907 19261
rect 9876 19236 9904 19264
rect 10778 19252 10784 19304
rect 10836 19292 10842 19304
rect 11072 19292 11100 19323
rect 10836 19264 11100 19292
rect 10836 19252 10842 19264
rect 7745 19227 7803 19233
rect 7745 19224 7757 19227
rect 7248 19196 7757 19224
rect 7248 19184 7254 19196
rect 7745 19193 7757 19196
rect 7791 19193 7803 19227
rect 7745 19187 7803 19193
rect 8021 19227 8079 19233
rect 8021 19193 8033 19227
rect 8067 19224 8079 19227
rect 9306 19224 9312 19236
rect 8067 19196 9312 19224
rect 8067 19193 8079 19196
rect 8021 19187 8079 19193
rect 9306 19184 9312 19196
rect 9364 19184 9370 19236
rect 9490 19224 9496 19236
rect 9451 19196 9496 19224
rect 9490 19184 9496 19196
rect 9548 19184 9554 19236
rect 9858 19184 9864 19236
rect 9916 19184 9922 19236
rect 10413 19227 10471 19233
rect 10413 19193 10425 19227
rect 10459 19224 10471 19227
rect 11164 19224 11192 19332
rect 11698 19320 11704 19372
rect 11756 19360 11762 19372
rect 11756 19332 11801 19360
rect 11756 19320 11762 19332
rect 11882 19320 11888 19372
rect 11940 19360 11946 19372
rect 12158 19369 12164 19372
rect 12152 19360 12164 19369
rect 11940 19332 11985 19360
rect 12119 19332 12164 19360
rect 11940 19320 11946 19332
rect 12152 19323 12164 19332
rect 12158 19320 12164 19323
rect 12216 19320 12222 19372
rect 12434 19320 12440 19372
rect 12492 19360 12498 19372
rect 13170 19360 13176 19372
rect 12492 19332 13176 19360
rect 12492 19320 12498 19332
rect 13170 19320 13176 19332
rect 13228 19320 13234 19372
rect 17034 19360 17040 19372
rect 13280 19332 17040 19360
rect 13280 19236 13308 19332
rect 17034 19320 17040 19332
rect 17092 19320 17098 19372
rect 13538 19292 13544 19304
rect 13499 19264 13544 19292
rect 13538 19252 13544 19264
rect 13596 19252 13602 19304
rect 19352 19301 19380 19400
rect 19978 19388 19984 19400
rect 20036 19388 20042 19440
rect 20438 19388 20444 19440
rect 20496 19428 20502 19440
rect 21376 19428 21404 19459
rect 20496 19400 21404 19428
rect 20496 19388 20502 19400
rect 19604 19363 19662 19369
rect 19604 19329 19616 19363
rect 19650 19360 19662 19363
rect 19886 19360 19892 19372
rect 19650 19332 19892 19360
rect 19650 19329 19662 19332
rect 19604 19323 19662 19329
rect 19886 19320 19892 19332
rect 19944 19320 19950 19372
rect 20714 19320 20720 19372
rect 20772 19360 20778 19372
rect 20809 19363 20867 19369
rect 20809 19360 20821 19363
rect 20772 19332 20821 19360
rect 20772 19320 20778 19332
rect 20809 19329 20821 19332
rect 20855 19329 20867 19363
rect 21174 19360 21180 19372
rect 21135 19332 21180 19360
rect 20809 19323 20867 19329
rect 21174 19320 21180 19332
rect 21232 19320 21238 19372
rect 19337 19295 19395 19301
rect 19337 19292 19349 19295
rect 19168 19264 19349 19292
rect 10459 19196 11192 19224
rect 10459 19193 10471 19196
rect 10413 19187 10471 19193
rect 11238 19184 11244 19236
rect 11296 19224 11302 19236
rect 13262 19224 13268 19236
rect 11296 19196 11744 19224
rect 13175 19196 13268 19224
rect 11296 19184 11302 19196
rect 2271 19128 2774 19156
rect 6733 19159 6791 19165
rect 2271 19125 2283 19128
rect 2225 19119 2283 19125
rect 6733 19125 6745 19159
rect 6779 19156 6791 19159
rect 7098 19156 7104 19168
rect 6779 19128 7104 19156
rect 6779 19125 6791 19128
rect 6733 19119 6791 19125
rect 7098 19116 7104 19128
rect 7156 19116 7162 19168
rect 7374 19156 7380 19168
rect 7335 19128 7380 19156
rect 7374 19116 7380 19128
rect 7432 19116 7438 19168
rect 8570 19156 8576 19168
rect 8531 19128 8576 19156
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 8757 19159 8815 19165
rect 8757 19125 8769 19159
rect 8803 19156 8815 19159
rect 8938 19156 8944 19168
rect 8803 19128 8944 19156
rect 8803 19125 8815 19128
rect 8757 19119 8815 19125
rect 8938 19116 8944 19128
rect 8996 19156 9002 19168
rect 9122 19156 9128 19168
rect 8996 19128 9128 19156
rect 8996 19116 9002 19128
rect 9122 19116 9128 19128
rect 9180 19116 9186 19168
rect 9217 19159 9275 19165
rect 9217 19125 9229 19159
rect 9263 19156 9275 19159
rect 9766 19156 9772 19168
rect 9263 19128 9772 19156
rect 9263 19125 9275 19128
rect 9217 19119 9275 19125
rect 9766 19116 9772 19128
rect 9824 19116 9830 19168
rect 10870 19156 10876 19168
rect 10831 19128 10876 19156
rect 10870 19116 10876 19128
rect 10928 19116 10934 19168
rect 10962 19116 10968 19168
rect 11020 19156 11026 19168
rect 11609 19159 11667 19165
rect 11609 19156 11621 19159
rect 11020 19128 11621 19156
rect 11020 19116 11026 19128
rect 11609 19125 11621 19128
rect 11655 19125 11667 19159
rect 11716 19156 11744 19196
rect 13262 19184 13268 19196
rect 13320 19184 13326 19236
rect 13446 19184 13452 19236
rect 13504 19224 13510 19236
rect 13817 19227 13875 19233
rect 13817 19224 13829 19227
rect 13504 19196 13829 19224
rect 13504 19184 13510 19196
rect 13817 19193 13829 19196
rect 13863 19224 13875 19227
rect 14642 19224 14648 19236
rect 13863 19196 14648 19224
rect 13863 19193 13875 19196
rect 13817 19187 13875 19193
rect 14642 19184 14648 19196
rect 14700 19184 14706 19236
rect 16942 19156 16948 19168
rect 11716 19128 16948 19156
rect 11609 19119 11667 19125
rect 16942 19116 16948 19128
rect 17000 19116 17006 19168
rect 17678 19116 17684 19168
rect 17736 19156 17742 19168
rect 19168 19165 19196 19264
rect 19337 19261 19349 19264
rect 19383 19261 19395 19295
rect 19337 19255 19395 19261
rect 19153 19159 19211 19165
rect 19153 19156 19165 19159
rect 17736 19128 19165 19156
rect 17736 19116 17742 19128
rect 19153 19125 19165 19128
rect 19199 19125 19211 19159
rect 20714 19156 20720 19168
rect 20675 19128 20720 19156
rect 19153 19119 19211 19125
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 7558 18952 7564 18964
rect 7519 18924 7564 18952
rect 7558 18912 7564 18924
rect 7616 18912 7622 18964
rect 8205 18955 8263 18961
rect 8205 18921 8217 18955
rect 8251 18952 8263 18955
rect 8478 18952 8484 18964
rect 8251 18924 8484 18952
rect 8251 18921 8263 18924
rect 8205 18915 8263 18921
rect 8478 18912 8484 18924
rect 8536 18912 8542 18964
rect 9122 18912 9128 18964
rect 9180 18952 9186 18964
rect 9582 18952 9588 18964
rect 9180 18924 9588 18952
rect 9180 18912 9186 18924
rect 9582 18912 9588 18924
rect 9640 18912 9646 18964
rect 9677 18955 9735 18961
rect 9677 18921 9689 18955
rect 9723 18952 9735 18955
rect 17126 18952 17132 18964
rect 9723 18924 12848 18952
rect 9723 18921 9735 18924
rect 9677 18915 9735 18921
rect 6914 18844 6920 18896
rect 6972 18884 6978 18896
rect 9306 18884 9312 18896
rect 6972 18856 9312 18884
rect 6972 18844 6978 18856
rect 9306 18844 9312 18856
rect 9364 18844 9370 18896
rect 9401 18887 9459 18893
rect 9401 18853 9413 18887
rect 9447 18884 9459 18887
rect 10042 18884 10048 18896
rect 9447 18856 10048 18884
rect 9447 18853 9459 18856
rect 9401 18847 9459 18853
rect 658 18776 664 18828
rect 716 18816 722 18828
rect 2041 18819 2099 18825
rect 2041 18816 2053 18819
rect 716 18788 2053 18816
rect 716 18776 722 18788
rect 1670 18748 1676 18760
rect 1631 18720 1676 18748
rect 1670 18708 1676 18720
rect 1728 18708 1734 18760
rect 1780 18757 1808 18788
rect 2041 18785 2053 18788
rect 2087 18785 2099 18819
rect 2041 18779 2099 18785
rect 8021 18819 8079 18825
rect 8021 18785 8033 18819
rect 8067 18816 8079 18819
rect 8570 18816 8576 18828
rect 8067 18788 8576 18816
rect 8067 18785 8079 18788
rect 8021 18779 8079 18785
rect 8570 18776 8576 18788
rect 8628 18776 8634 18828
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18717 1823 18751
rect 8294 18748 8300 18760
rect 8207 18720 8300 18748
rect 1765 18711 1823 18717
rect 8294 18708 8300 18720
rect 8352 18748 8358 18760
rect 8665 18751 8723 18757
rect 8665 18748 8677 18751
rect 8352 18720 8677 18748
rect 8352 18708 8358 18720
rect 8665 18717 8677 18720
rect 8711 18717 8723 18751
rect 8665 18711 8723 18717
rect 8754 18708 8760 18760
rect 8812 18748 8818 18760
rect 9508 18757 9536 18856
rect 10042 18844 10048 18856
rect 10100 18844 10106 18896
rect 12820 18884 12848 18924
rect 13372 18924 17132 18952
rect 13372 18884 13400 18924
rect 17126 18912 17132 18924
rect 17184 18912 17190 18964
rect 20898 18912 20904 18964
rect 20956 18952 20962 18964
rect 21177 18955 21235 18961
rect 21177 18952 21189 18955
rect 20956 18924 21189 18952
rect 20956 18912 20962 18924
rect 21177 18921 21189 18924
rect 21223 18921 21235 18955
rect 21177 18915 21235 18921
rect 12820 18856 13400 18884
rect 13173 18819 13231 18825
rect 13173 18785 13185 18819
rect 13219 18816 13231 18819
rect 13357 18819 13415 18825
rect 13357 18816 13369 18819
rect 13219 18788 13369 18816
rect 13219 18785 13231 18788
rect 13173 18779 13231 18785
rect 13357 18785 13369 18788
rect 13403 18816 13415 18819
rect 13446 18816 13452 18828
rect 13403 18788 13452 18816
rect 13403 18785 13415 18788
rect 13357 18779 13415 18785
rect 13446 18776 13452 18788
rect 13504 18776 13510 18828
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 8812 18720 8953 18748
rect 8812 18708 8818 18720
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 9493 18751 9551 18757
rect 9493 18717 9505 18751
rect 9539 18717 9551 18751
rect 9766 18748 9772 18760
rect 9727 18720 9772 18748
rect 9493 18711 9551 18717
rect 9766 18708 9772 18720
rect 9824 18708 9830 18760
rect 10045 18751 10103 18757
rect 10045 18717 10057 18751
rect 10091 18748 10103 18751
rect 11517 18751 11575 18757
rect 11517 18748 11529 18751
rect 10091 18720 11529 18748
rect 10091 18717 10103 18720
rect 10045 18711 10103 18717
rect 11517 18717 11529 18720
rect 11563 18748 11575 18751
rect 12894 18748 12900 18760
rect 11563 18720 12900 18748
rect 11563 18717 11575 18720
rect 11517 18711 11575 18717
rect 12894 18708 12900 18720
rect 12952 18708 12958 18760
rect 14642 18708 14648 18760
rect 14700 18748 14706 18760
rect 14737 18751 14795 18757
rect 14737 18748 14749 18751
rect 14700 18720 14749 18748
rect 14700 18708 14706 18720
rect 14737 18717 14749 18720
rect 14783 18748 14795 18751
rect 16301 18751 16359 18757
rect 16301 18748 16313 18751
rect 14783 18720 16313 18748
rect 14783 18717 14795 18720
rect 14737 18711 14795 18717
rect 16301 18717 16313 18720
rect 16347 18748 16359 18751
rect 16669 18751 16727 18757
rect 16669 18748 16681 18751
rect 16347 18720 16681 18748
rect 16347 18717 16359 18720
rect 16301 18711 16359 18717
rect 16669 18717 16681 18720
rect 16715 18748 16727 18751
rect 16942 18748 16948 18760
rect 16715 18720 16948 18748
rect 16715 18717 16727 18720
rect 16669 18711 16727 18717
rect 16942 18708 16948 18720
rect 17000 18748 17006 18760
rect 17678 18748 17684 18760
rect 17000 18720 17684 18748
rect 17000 18708 17006 18720
rect 17678 18708 17684 18720
rect 17736 18748 17742 18760
rect 18233 18751 18291 18757
rect 18233 18748 18245 18751
rect 17736 18720 18245 18748
rect 17736 18708 17742 18720
rect 18233 18717 18245 18720
rect 18279 18748 18291 18751
rect 18325 18751 18383 18757
rect 18325 18748 18337 18751
rect 18279 18720 18337 18748
rect 18279 18717 18291 18720
rect 18233 18711 18291 18717
rect 18325 18717 18337 18720
rect 18371 18717 18383 18751
rect 18325 18711 18383 18717
rect 20346 18708 20352 18760
rect 20404 18748 20410 18760
rect 20634 18751 20692 18757
rect 20634 18748 20646 18751
rect 20404 18720 20646 18748
rect 20404 18708 20410 18720
rect 20634 18717 20646 18720
rect 20680 18717 20692 18751
rect 20634 18711 20692 18717
rect 20806 18708 20812 18760
rect 20864 18748 20870 18760
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 20864 18720 20913 18748
rect 20864 18708 20870 18720
rect 20901 18717 20913 18720
rect 20947 18717 20959 18751
rect 20901 18711 20959 18717
rect 7469 18683 7527 18689
rect 7469 18649 7481 18683
rect 7515 18680 7527 18683
rect 7650 18680 7656 18692
rect 7515 18652 7656 18680
rect 7515 18649 7527 18652
rect 7469 18643 7527 18649
rect 7650 18640 7656 18652
rect 7708 18680 7714 18692
rect 8202 18680 8208 18692
rect 7708 18652 8208 18680
rect 7708 18640 7714 18652
rect 8202 18640 8208 18652
rect 8260 18640 8266 18692
rect 10312 18683 10370 18689
rect 9140 18652 10272 18680
rect 1486 18612 1492 18624
rect 1447 18584 1492 18612
rect 1486 18572 1492 18584
rect 1544 18572 1550 18624
rect 1949 18615 2007 18621
rect 1949 18581 1961 18615
rect 1995 18612 2007 18615
rect 5442 18612 5448 18624
rect 1995 18584 5448 18612
rect 1995 18581 2007 18584
rect 1949 18575 2007 18581
rect 5442 18572 5448 18584
rect 5500 18572 5506 18624
rect 8478 18612 8484 18624
rect 8439 18584 8484 18612
rect 8478 18572 8484 18584
rect 8536 18572 8542 18624
rect 9140 18621 9168 18652
rect 9125 18615 9183 18621
rect 9125 18581 9137 18615
rect 9171 18581 9183 18615
rect 9125 18575 9183 18581
rect 9214 18572 9220 18624
rect 9272 18612 9278 18624
rect 9490 18612 9496 18624
rect 9272 18584 9496 18612
rect 9272 18572 9278 18584
rect 9490 18572 9496 18584
rect 9548 18572 9554 18624
rect 9950 18612 9956 18624
rect 9911 18584 9956 18612
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 10244 18612 10272 18652
rect 10312 18649 10324 18683
rect 10358 18680 10370 18683
rect 11054 18680 11060 18692
rect 10358 18652 11060 18680
rect 10358 18649 10370 18652
rect 10312 18643 10370 18649
rect 11054 18640 11060 18652
rect 11112 18640 11118 18692
rect 11784 18683 11842 18689
rect 11784 18649 11796 18683
rect 11830 18649 11842 18683
rect 11784 18643 11842 18649
rect 11238 18612 11244 18624
rect 10244 18584 11244 18612
rect 11238 18572 11244 18584
rect 11296 18572 11302 18624
rect 11425 18615 11483 18621
rect 11425 18581 11437 18615
rect 11471 18612 11483 18615
rect 11808 18612 11836 18643
rect 11882 18640 11888 18692
rect 11940 18680 11946 18692
rect 14982 18683 15040 18689
rect 14982 18680 14994 18683
rect 11940 18652 14994 18680
rect 11940 18640 11946 18652
rect 14982 18649 14994 18652
rect 15028 18649 15040 18683
rect 17988 18683 18046 18689
rect 14982 18643 15040 18649
rect 16132 18652 17908 18680
rect 16132 18624 16160 18652
rect 11974 18612 11980 18624
rect 11471 18584 11980 18612
rect 11471 18581 11483 18584
rect 11425 18575 11483 18581
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 12897 18615 12955 18621
rect 12897 18581 12909 18615
rect 12943 18612 12955 18615
rect 13078 18612 13084 18624
rect 12943 18584 13084 18612
rect 12943 18581 12955 18584
rect 12897 18575 12955 18581
rect 13078 18572 13084 18584
rect 13136 18572 13142 18624
rect 16114 18612 16120 18624
rect 16075 18584 16120 18612
rect 16114 18572 16120 18584
rect 16172 18572 16178 18624
rect 16390 18572 16396 18624
rect 16448 18612 16454 18624
rect 16853 18615 16911 18621
rect 16853 18612 16865 18615
rect 16448 18584 16865 18612
rect 16448 18572 16454 18584
rect 16853 18581 16865 18584
rect 16899 18581 16911 18615
rect 17880 18612 17908 18652
rect 17988 18649 18000 18683
rect 18034 18680 18046 18683
rect 18138 18680 18144 18692
rect 18034 18652 18144 18680
rect 18034 18649 18046 18652
rect 17988 18643 18046 18649
rect 18138 18640 18144 18652
rect 18196 18640 18202 18692
rect 20438 18680 20444 18692
rect 19444 18652 20444 18680
rect 19444 18612 19472 18652
rect 20438 18640 20444 18652
rect 20496 18640 20502 18692
rect 20916 18680 20944 18711
rect 20990 18708 20996 18760
rect 21048 18748 21054 18760
rect 21048 18720 21093 18748
rect 21048 18708 21054 18720
rect 21361 18683 21419 18689
rect 21361 18680 21373 18683
rect 20916 18652 21373 18680
rect 21361 18649 21373 18652
rect 21407 18649 21419 18683
rect 21361 18643 21419 18649
rect 17880 18584 19472 18612
rect 19521 18615 19579 18621
rect 16853 18575 16911 18581
rect 19521 18581 19533 18615
rect 19567 18612 19579 18615
rect 20070 18612 20076 18624
rect 19567 18584 20076 18612
rect 19567 18581 19579 18584
rect 19521 18575 19579 18581
rect 20070 18572 20076 18584
rect 20128 18572 20134 18624
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 2038 18368 2044 18420
rect 2096 18408 2102 18420
rect 2133 18411 2191 18417
rect 2133 18408 2145 18411
rect 2096 18380 2145 18408
rect 2096 18368 2102 18380
rect 2133 18377 2145 18380
rect 2179 18377 2191 18411
rect 2133 18371 2191 18377
rect 5537 18411 5595 18417
rect 5537 18377 5549 18411
rect 5583 18408 5595 18411
rect 5810 18408 5816 18420
rect 5583 18380 5816 18408
rect 5583 18377 5595 18380
rect 5537 18371 5595 18377
rect 5810 18368 5816 18380
rect 5868 18368 5874 18420
rect 5902 18368 5908 18420
rect 5960 18408 5966 18420
rect 8665 18411 8723 18417
rect 8665 18408 8677 18411
rect 5960 18380 8677 18408
rect 5960 18368 5966 18380
rect 8665 18377 8677 18380
rect 8711 18377 8723 18411
rect 8665 18371 8723 18377
rect 9674 18368 9680 18420
rect 9732 18408 9738 18420
rect 9769 18411 9827 18417
rect 9769 18408 9781 18411
rect 9732 18380 9781 18408
rect 9732 18368 9738 18380
rect 9769 18377 9781 18380
rect 9815 18377 9827 18411
rect 9769 18371 9827 18377
rect 10318 18368 10324 18420
rect 10376 18408 10382 18420
rect 10505 18411 10563 18417
rect 10505 18408 10517 18411
rect 10376 18380 10517 18408
rect 10376 18368 10382 18380
rect 10505 18377 10517 18380
rect 10551 18377 10563 18411
rect 19518 18408 19524 18420
rect 10505 18371 10563 18377
rect 10612 18380 19524 18408
rect 5258 18300 5264 18352
rect 5316 18340 5322 18352
rect 5629 18343 5687 18349
rect 5629 18340 5641 18343
rect 5316 18312 5641 18340
rect 5316 18300 5322 18312
rect 5629 18309 5641 18312
rect 5675 18340 5687 18343
rect 5718 18340 5724 18352
rect 5675 18312 5724 18340
rect 5675 18309 5687 18312
rect 5629 18303 5687 18309
rect 5718 18300 5724 18312
rect 5776 18300 5782 18352
rect 6549 18343 6607 18349
rect 6549 18309 6561 18343
rect 6595 18340 6607 18343
rect 6914 18340 6920 18352
rect 6595 18312 6920 18340
rect 6595 18309 6607 18312
rect 6549 18303 6607 18309
rect 6914 18300 6920 18312
rect 6972 18300 6978 18352
rect 10612 18340 10640 18380
rect 19518 18368 19524 18380
rect 19576 18408 19582 18420
rect 19886 18408 19892 18420
rect 19576 18380 19892 18408
rect 19576 18368 19582 18380
rect 19886 18368 19892 18380
rect 19944 18368 19950 18420
rect 20806 18368 20812 18420
rect 20864 18408 20870 18420
rect 21085 18411 21143 18417
rect 21085 18408 21097 18411
rect 20864 18380 21097 18408
rect 20864 18368 20870 18380
rect 10778 18340 10784 18352
rect 8864 18312 10640 18340
rect 10739 18312 10784 18340
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18272 1731 18275
rect 1946 18272 1952 18284
rect 1719 18244 1952 18272
rect 1719 18241 1731 18244
rect 1673 18235 1731 18241
rect 1946 18232 1952 18244
rect 2004 18232 2010 18284
rect 2041 18275 2099 18281
rect 2041 18241 2053 18275
rect 2087 18272 2099 18275
rect 2222 18272 2228 18284
rect 2087 18244 2228 18272
rect 2087 18241 2099 18244
rect 2041 18235 2099 18241
rect 2222 18232 2228 18244
rect 2280 18232 2286 18284
rect 2317 18275 2375 18281
rect 2317 18241 2329 18275
rect 2363 18272 2375 18275
rect 2866 18272 2872 18284
rect 2363 18244 2872 18272
rect 2363 18241 2375 18244
rect 2317 18235 2375 18241
rect 2866 18232 2872 18244
rect 2924 18232 2930 18284
rect 7650 18232 7656 18284
rect 7708 18272 7714 18284
rect 8573 18275 8631 18281
rect 8573 18272 8585 18275
rect 7708 18244 8585 18272
rect 7708 18232 7714 18244
rect 8573 18241 8585 18244
rect 8619 18241 8631 18275
rect 8573 18235 8631 18241
rect 4982 18164 4988 18216
rect 5040 18204 5046 18216
rect 5721 18207 5779 18213
rect 5721 18204 5733 18207
rect 5040 18176 5733 18204
rect 5040 18164 5046 18176
rect 5721 18173 5733 18176
rect 5767 18204 5779 18207
rect 6365 18207 6423 18213
rect 6365 18204 6377 18207
rect 5767 18176 6377 18204
rect 5767 18173 5779 18176
rect 5721 18167 5779 18173
rect 6365 18173 6377 18176
rect 6411 18173 6423 18207
rect 7926 18204 7932 18216
rect 7887 18176 7932 18204
rect 6365 18167 6423 18173
rect 7926 18164 7932 18176
rect 7984 18164 7990 18216
rect 8864 18213 8892 18312
rect 10778 18300 10784 18312
rect 10836 18300 10842 18352
rect 11333 18343 11391 18349
rect 11333 18309 11345 18343
rect 11379 18340 11391 18343
rect 12526 18340 12532 18352
rect 11379 18312 12532 18340
rect 11379 18309 11391 18312
rect 11333 18303 11391 18309
rect 12526 18300 12532 18312
rect 12584 18340 12590 18352
rect 14642 18340 14648 18352
rect 12584 18312 12940 18340
rect 12584 18300 12590 18312
rect 12912 18284 12940 18312
rect 14476 18312 14648 18340
rect 9493 18275 9551 18281
rect 9214 18216 9220 18268
rect 9272 18256 9278 18268
rect 9272 18228 9317 18256
rect 9493 18241 9505 18275
rect 9539 18241 9551 18275
rect 9493 18235 9551 18241
rect 9953 18275 10011 18281
rect 9953 18241 9965 18275
rect 9999 18241 10011 18275
rect 9953 18235 10011 18241
rect 9272 18216 9278 18228
rect 8849 18207 8907 18213
rect 8849 18173 8861 18207
rect 8895 18173 8907 18207
rect 9508 18204 9536 18235
rect 9968 18204 9996 18235
rect 10686 18232 10692 18284
rect 10744 18272 10750 18284
rect 10873 18275 10931 18281
rect 10873 18272 10885 18275
rect 10744 18244 10885 18272
rect 10744 18232 10750 18244
rect 10873 18241 10885 18244
rect 10919 18241 10931 18275
rect 10873 18235 10931 18241
rect 11698 18232 11704 18284
rect 11756 18272 11762 18284
rect 12641 18275 12699 18281
rect 12641 18272 12653 18275
rect 11756 18244 12653 18272
rect 11756 18232 11762 18244
rect 12641 18241 12653 18244
rect 12687 18272 12699 18275
rect 12687 18244 12848 18272
rect 12687 18241 12699 18244
rect 12641 18235 12699 18241
rect 8849 18167 8907 18173
rect 9416 18176 9536 18204
rect 9600 18176 9996 18204
rect 12820 18204 12848 18244
rect 12894 18232 12900 18284
rect 12952 18281 12958 18284
rect 12952 18275 12966 18281
rect 12954 18272 12966 18275
rect 13446 18272 13452 18284
rect 12954 18244 13452 18272
rect 12954 18241 12966 18244
rect 12952 18235 12966 18241
rect 12952 18232 12958 18235
rect 13446 18232 13452 18244
rect 13504 18232 13510 18284
rect 13814 18232 13820 18284
rect 13872 18272 13878 18284
rect 14476 18281 14504 18312
rect 14642 18300 14648 18312
rect 14700 18300 14706 18352
rect 18064 18312 19564 18340
rect 14194 18275 14252 18281
rect 14194 18272 14206 18275
rect 13872 18244 14206 18272
rect 13872 18232 13878 18244
rect 14194 18241 14206 18244
rect 14240 18272 14252 18275
rect 14461 18275 14519 18281
rect 14240 18244 14412 18272
rect 14240 18241 14252 18244
rect 14194 18235 14252 18241
rect 14384 18204 14412 18244
rect 14461 18241 14473 18275
rect 14507 18241 14519 18275
rect 14461 18235 14519 18241
rect 16206 18232 16212 18284
rect 16264 18281 16270 18284
rect 16264 18272 16276 18281
rect 16485 18275 16543 18281
rect 16264 18244 16309 18272
rect 16264 18235 16276 18244
rect 16485 18241 16497 18275
rect 16531 18272 16543 18275
rect 16574 18272 16580 18284
rect 16531 18244 16580 18272
rect 16531 18241 16543 18244
rect 16485 18235 16543 18241
rect 16264 18232 16270 18235
rect 16574 18232 16580 18244
rect 16632 18272 16638 18284
rect 16942 18272 16948 18284
rect 16632 18244 16948 18272
rect 16632 18232 16638 18244
rect 16942 18232 16948 18244
rect 17000 18232 17006 18284
rect 17402 18232 17408 18284
rect 17460 18272 17466 18284
rect 17782 18275 17840 18281
rect 17782 18272 17794 18275
rect 17460 18244 17794 18272
rect 17460 18232 17466 18244
rect 17782 18241 17794 18244
rect 17828 18241 17840 18275
rect 17782 18235 17840 18241
rect 18064 18213 18092 18312
rect 18138 18232 18144 18284
rect 18196 18272 18202 18284
rect 19536 18281 19564 18312
rect 19610 18300 19616 18352
rect 19668 18340 19674 18352
rect 19668 18312 20852 18340
rect 19668 18300 19674 18312
rect 19254 18275 19312 18281
rect 19254 18272 19266 18275
rect 18196 18244 19266 18272
rect 18196 18232 18202 18244
rect 19254 18241 19266 18244
rect 19300 18241 19312 18275
rect 19254 18235 19312 18241
rect 19521 18275 19579 18281
rect 19521 18241 19533 18275
rect 19567 18241 19579 18275
rect 19521 18235 19579 18241
rect 20438 18232 20444 18284
rect 20496 18272 20502 18284
rect 20726 18275 20784 18281
rect 20726 18272 20738 18275
rect 20496 18244 20738 18272
rect 20496 18232 20502 18244
rect 20726 18241 20738 18244
rect 20772 18241 20784 18275
rect 20824 18272 20852 18312
rect 21008 18281 21036 18380
rect 21085 18377 21097 18380
rect 21131 18377 21143 18411
rect 21085 18371 21143 18377
rect 21453 18411 21511 18417
rect 21453 18377 21465 18411
rect 21499 18408 21511 18411
rect 21634 18408 21640 18420
rect 21499 18380 21640 18408
rect 21499 18377 21511 18380
rect 21453 18371 21511 18377
rect 21634 18368 21640 18380
rect 21692 18368 21698 18420
rect 20993 18275 21051 18281
rect 20824 18244 20953 18272
rect 20726 18235 20784 18241
rect 18049 18207 18107 18213
rect 12820 18176 13400 18204
rect 14384 18176 15148 18204
rect 1854 18136 1860 18148
rect 1815 18108 1860 18136
rect 1854 18096 1860 18108
rect 1912 18096 1918 18148
rect 8478 18096 8484 18148
rect 8536 18136 8542 18148
rect 9122 18136 9128 18148
rect 8536 18108 9128 18136
rect 8536 18096 8542 18108
rect 9122 18096 9128 18108
rect 9180 18096 9186 18148
rect 9416 18136 9444 18176
rect 9232 18108 9444 18136
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 5169 18071 5227 18077
rect 5169 18037 5181 18071
rect 5215 18068 5227 18071
rect 5350 18068 5356 18080
rect 5215 18040 5356 18068
rect 5215 18037 5227 18040
rect 5169 18031 5227 18037
rect 5350 18028 5356 18040
rect 5408 18028 5414 18080
rect 7650 18028 7656 18080
rect 7708 18068 7714 18080
rect 7745 18071 7803 18077
rect 7745 18068 7757 18071
rect 7708 18040 7757 18068
rect 7708 18028 7714 18040
rect 7745 18037 7757 18040
rect 7791 18037 7803 18071
rect 7745 18031 7803 18037
rect 7834 18028 7840 18080
rect 7892 18068 7898 18080
rect 8205 18071 8263 18077
rect 8205 18068 8217 18071
rect 7892 18040 8217 18068
rect 7892 18028 7898 18040
rect 8205 18037 8217 18040
rect 8251 18037 8263 18071
rect 8205 18031 8263 18037
rect 8294 18028 8300 18080
rect 8352 18068 8358 18080
rect 9232 18068 9260 18108
rect 9490 18096 9496 18148
rect 9548 18136 9554 18148
rect 9600 18136 9628 18176
rect 9548 18108 9628 18136
rect 9677 18139 9735 18145
rect 9548 18096 9554 18108
rect 9677 18105 9689 18139
rect 9723 18136 9735 18139
rect 9858 18136 9864 18148
rect 9723 18108 9864 18136
rect 9723 18105 9735 18108
rect 9677 18099 9735 18105
rect 9858 18096 9864 18108
rect 9916 18096 9922 18148
rect 8352 18040 9260 18068
rect 8352 18028 8358 18040
rect 9398 18028 9404 18080
rect 9456 18068 9462 18080
rect 10137 18071 10195 18077
rect 9456 18040 9501 18068
rect 9456 18028 9462 18040
rect 10137 18037 10149 18071
rect 10183 18068 10195 18071
rect 10226 18068 10232 18080
rect 10183 18040 10232 18068
rect 10183 18037 10195 18040
rect 10137 18031 10195 18037
rect 10226 18028 10232 18040
rect 10284 18028 10290 18080
rect 10410 18028 10416 18080
rect 10468 18068 10474 18080
rect 10686 18068 10692 18080
rect 10468 18040 10692 18068
rect 10468 18028 10474 18040
rect 10686 18028 10692 18040
rect 10744 18028 10750 18080
rect 11514 18068 11520 18080
rect 11475 18040 11520 18068
rect 11514 18028 11520 18040
rect 11572 18028 11578 18080
rect 12986 18028 12992 18080
rect 13044 18068 13050 18080
rect 13081 18071 13139 18077
rect 13081 18068 13093 18071
rect 13044 18040 13093 18068
rect 13044 18028 13050 18040
rect 13081 18037 13093 18040
rect 13127 18037 13139 18071
rect 13372 18068 13400 18176
rect 15120 18145 15148 18176
rect 18049 18173 18061 18207
rect 18095 18173 18107 18207
rect 20925 18204 20953 18244
rect 20993 18241 21005 18275
rect 21039 18241 21051 18275
rect 20993 18235 21051 18241
rect 21269 18275 21327 18281
rect 21269 18241 21281 18275
rect 21315 18241 21327 18275
rect 21269 18235 21327 18241
rect 21284 18204 21312 18235
rect 20925 18176 21312 18204
rect 18049 18167 18107 18173
rect 15105 18139 15163 18145
rect 15105 18105 15117 18139
rect 15151 18105 15163 18139
rect 15105 18099 15163 18105
rect 14642 18068 14648 18080
rect 13372 18040 14648 18068
rect 13081 18031 13139 18037
rect 14642 18028 14648 18040
rect 14700 18028 14706 18080
rect 16206 18028 16212 18080
rect 16264 18068 16270 18080
rect 16669 18071 16727 18077
rect 16669 18068 16681 18071
rect 16264 18040 16681 18068
rect 16264 18028 16270 18040
rect 16669 18037 16681 18040
rect 16715 18037 16727 18071
rect 16669 18031 16727 18037
rect 17862 18028 17868 18080
rect 17920 18068 17926 18080
rect 18064 18068 18092 18167
rect 19518 18096 19524 18148
rect 19576 18136 19582 18148
rect 19613 18139 19671 18145
rect 19613 18136 19625 18139
rect 19576 18108 19625 18136
rect 19576 18096 19582 18108
rect 19613 18105 19625 18108
rect 19659 18105 19671 18139
rect 19613 18099 19671 18105
rect 17920 18040 18092 18068
rect 17920 18028 17926 18040
rect 18138 18028 18144 18080
rect 18196 18068 18202 18080
rect 18196 18040 18241 18068
rect 18196 18028 18202 18040
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 6914 17824 6920 17876
rect 6972 17824 6978 17876
rect 8573 17867 8631 17873
rect 8573 17833 8585 17867
rect 8619 17864 8631 17867
rect 9490 17864 9496 17876
rect 8619 17836 9496 17864
rect 8619 17833 8631 17836
rect 8573 17827 8631 17833
rect 9490 17824 9496 17836
rect 9548 17824 9554 17876
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 10226 17864 10232 17876
rect 9732 17836 10232 17864
rect 9732 17824 9738 17836
rect 10226 17824 10232 17836
rect 10284 17824 10290 17876
rect 10410 17824 10416 17876
rect 10468 17864 10474 17876
rect 12802 17864 12808 17876
rect 10468 17836 12808 17864
rect 10468 17824 10474 17836
rect 12802 17824 12808 17836
rect 12860 17824 12866 17876
rect 12894 17824 12900 17876
rect 12952 17864 12958 17876
rect 13173 17867 13231 17873
rect 13173 17864 13185 17867
rect 12952 17836 13185 17864
rect 12952 17824 12958 17836
rect 5166 17728 5172 17740
rect 5127 17700 5172 17728
rect 5166 17688 5172 17700
rect 5224 17688 5230 17740
rect 5350 17728 5356 17740
rect 5311 17700 5356 17728
rect 5350 17688 5356 17700
rect 5408 17688 5414 17740
rect 5994 17688 6000 17740
rect 6052 17728 6058 17740
rect 6365 17731 6423 17737
rect 6365 17728 6377 17731
rect 6052 17700 6377 17728
rect 6052 17688 6058 17700
rect 6365 17697 6377 17700
rect 6411 17697 6423 17731
rect 6365 17691 6423 17697
rect 6457 17731 6515 17737
rect 6457 17697 6469 17731
rect 6503 17728 6515 17731
rect 6932 17728 6960 17824
rect 7742 17756 7748 17808
rect 7800 17796 7806 17808
rect 9858 17796 9864 17808
rect 7800 17768 9864 17796
rect 7800 17756 7806 17768
rect 9858 17756 9864 17768
rect 9916 17756 9922 17808
rect 7282 17728 7288 17740
rect 6503 17700 7288 17728
rect 6503 17697 6515 17700
rect 6457 17691 6515 17697
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17660 1731 17663
rect 2498 17660 2504 17672
rect 1719 17632 2504 17660
rect 1719 17629 1731 17632
rect 1673 17623 1731 17629
rect 2498 17620 2504 17632
rect 2556 17620 2562 17672
rect 4798 17620 4804 17672
rect 4856 17660 4862 17672
rect 5442 17660 5448 17672
rect 4856 17632 5448 17660
rect 4856 17620 4862 17632
rect 5442 17620 5448 17632
rect 5500 17660 5506 17672
rect 6273 17663 6331 17669
rect 6273 17660 6285 17663
rect 5500 17632 6285 17660
rect 5500 17620 5506 17632
rect 6273 17629 6285 17632
rect 6319 17629 6331 17663
rect 6380 17660 6408 17691
rect 7282 17688 7288 17700
rect 7340 17688 7346 17740
rect 8021 17731 8079 17737
rect 8021 17697 8033 17731
rect 8067 17728 8079 17731
rect 9674 17728 9680 17740
rect 8067 17700 9680 17728
rect 8067 17697 8079 17700
rect 8021 17691 8079 17697
rect 9674 17688 9680 17700
rect 9732 17688 9738 17740
rect 13096 17737 13124 17836
rect 13173 17833 13185 17836
rect 13219 17864 13231 17867
rect 13541 17867 13599 17873
rect 13541 17864 13553 17867
rect 13219 17836 13553 17864
rect 13219 17833 13231 17836
rect 13173 17827 13231 17833
rect 13541 17833 13553 17836
rect 13587 17833 13599 17867
rect 13541 17827 13599 17833
rect 13722 17824 13728 17876
rect 13780 17864 13786 17876
rect 18322 17864 18328 17876
rect 13780 17836 18328 17864
rect 13780 17824 13786 17836
rect 18322 17824 18328 17836
rect 18380 17824 18386 17876
rect 13449 17799 13507 17805
rect 13449 17765 13461 17799
rect 13495 17796 13507 17799
rect 16390 17796 16396 17808
rect 13495 17768 16396 17796
rect 13495 17765 13507 17768
rect 13449 17759 13507 17765
rect 13081 17731 13139 17737
rect 13081 17697 13093 17731
rect 13127 17697 13139 17731
rect 13081 17691 13139 17697
rect 13170 17688 13176 17740
rect 13228 17728 13234 17740
rect 13464 17728 13492 17759
rect 16390 17756 16396 17768
rect 16448 17756 16454 17808
rect 17770 17756 17776 17808
rect 17828 17796 17834 17808
rect 17865 17799 17923 17805
rect 17865 17796 17877 17799
rect 17828 17768 17877 17796
rect 17828 17756 17834 17768
rect 17865 17765 17877 17768
rect 17911 17765 17923 17799
rect 17865 17759 17923 17765
rect 13228 17700 13492 17728
rect 13228 17688 13234 17700
rect 6546 17660 6552 17672
rect 6380 17632 6552 17660
rect 6273 17623 6331 17629
rect 6546 17620 6552 17632
rect 6604 17620 6610 17672
rect 9398 17620 9404 17672
rect 9456 17660 9462 17672
rect 16206 17660 16212 17672
rect 9456 17632 16212 17660
rect 9456 17620 9462 17632
rect 16206 17620 16212 17632
rect 16264 17620 16270 17672
rect 16485 17663 16543 17669
rect 16485 17629 16497 17663
rect 16531 17660 16543 17663
rect 16574 17660 16580 17672
rect 16531 17632 16580 17660
rect 16531 17629 16543 17632
rect 16485 17623 16543 17629
rect 16574 17620 16580 17632
rect 16632 17660 16638 17672
rect 17862 17660 17868 17672
rect 16632 17632 17868 17660
rect 16632 17620 16638 17632
rect 17862 17620 17868 17632
rect 17920 17660 17926 17672
rect 17957 17663 18015 17669
rect 17957 17660 17969 17663
rect 17920 17632 17969 17660
rect 17920 17620 17926 17632
rect 17957 17629 17969 17632
rect 18003 17660 18015 17663
rect 18141 17663 18199 17669
rect 18141 17660 18153 17663
rect 18003 17632 18153 17660
rect 18003 17629 18015 17632
rect 17957 17623 18015 17629
rect 18141 17629 18153 17632
rect 18187 17660 18199 17663
rect 19613 17663 19671 17669
rect 19613 17660 19625 17663
rect 18187 17632 19625 17660
rect 18187 17629 18199 17632
rect 18141 17623 18199 17629
rect 19613 17629 19625 17632
rect 19659 17660 19671 17663
rect 19797 17663 19855 17669
rect 19797 17660 19809 17663
rect 19659 17632 19809 17660
rect 19659 17629 19671 17632
rect 19613 17623 19671 17629
rect 19797 17629 19809 17632
rect 19843 17629 19855 17663
rect 21266 17660 21272 17672
rect 21227 17632 21272 17660
rect 19797 17623 19855 17629
rect 21266 17620 21272 17632
rect 21324 17620 21330 17672
rect 7466 17552 7472 17604
rect 7524 17592 7530 17604
rect 8205 17595 8263 17601
rect 8205 17592 8217 17595
rect 7524 17564 8217 17592
rect 7524 17552 7530 17564
rect 8205 17561 8217 17564
rect 8251 17561 8263 17595
rect 8205 17555 8263 17561
rect 12158 17552 12164 17604
rect 12216 17592 12222 17604
rect 12814 17595 12872 17601
rect 12814 17592 12826 17595
rect 12216 17564 12826 17592
rect 12216 17552 12222 17564
rect 12814 17561 12826 17564
rect 12860 17561 12872 17595
rect 12814 17555 12872 17561
rect 12986 17552 12992 17604
rect 13044 17592 13050 17604
rect 16390 17592 16396 17604
rect 13044 17564 16396 17592
rect 13044 17552 13050 17564
rect 16390 17552 16396 17564
rect 16448 17552 16454 17604
rect 16752 17595 16810 17601
rect 16752 17561 16764 17595
rect 16798 17592 16810 17595
rect 17034 17592 17040 17604
rect 16798 17564 17040 17592
rect 16798 17561 16810 17564
rect 16752 17555 16810 17561
rect 17034 17552 17040 17564
rect 17092 17552 17098 17604
rect 20070 17601 20076 17604
rect 20064 17592 20076 17601
rect 20031 17564 20076 17592
rect 20064 17555 20076 17564
rect 20070 17552 20076 17555
rect 20128 17552 20134 17604
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 4890 17484 4896 17536
rect 4948 17524 4954 17536
rect 5445 17527 5503 17533
rect 5445 17524 5457 17527
rect 4948 17496 5457 17524
rect 4948 17484 4954 17496
rect 5445 17493 5457 17496
rect 5491 17493 5503 17527
rect 5445 17487 5503 17493
rect 5718 17484 5724 17536
rect 5776 17524 5782 17536
rect 5813 17527 5871 17533
rect 5813 17524 5825 17527
rect 5776 17496 5825 17524
rect 5776 17484 5782 17496
rect 5813 17493 5825 17496
rect 5859 17493 5871 17527
rect 5813 17487 5871 17493
rect 5902 17484 5908 17536
rect 5960 17524 5966 17536
rect 5960 17496 6005 17524
rect 5960 17484 5966 17496
rect 7374 17484 7380 17536
rect 7432 17524 7438 17536
rect 8113 17527 8171 17533
rect 8113 17524 8125 17527
rect 7432 17496 8125 17524
rect 7432 17484 7438 17496
rect 8113 17493 8125 17496
rect 8159 17493 8171 17527
rect 8113 17487 8171 17493
rect 9122 17484 9128 17536
rect 9180 17524 9186 17536
rect 9493 17527 9551 17533
rect 9493 17524 9505 17527
rect 9180 17496 9505 17524
rect 9180 17484 9186 17496
rect 9493 17493 9505 17496
rect 9539 17493 9551 17527
rect 9493 17487 9551 17493
rect 9861 17527 9919 17533
rect 9861 17493 9873 17527
rect 9907 17524 9919 17527
rect 9950 17524 9956 17536
rect 9907 17496 9956 17524
rect 9907 17493 9919 17496
rect 9861 17487 9919 17493
rect 9950 17484 9956 17496
rect 10008 17484 10014 17536
rect 11698 17524 11704 17536
rect 11659 17496 11704 17524
rect 11698 17484 11704 17496
rect 11756 17524 11762 17536
rect 16206 17524 16212 17536
rect 11756 17496 16212 17524
rect 11756 17484 11762 17496
rect 16206 17484 16212 17496
rect 16264 17484 16270 17536
rect 21174 17524 21180 17536
rect 21135 17496 21180 17524
rect 21174 17484 21180 17496
rect 21232 17484 21238 17536
rect 21450 17524 21456 17536
rect 21411 17496 21456 17524
rect 21450 17484 21456 17496
rect 21508 17484 21514 17536
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 1762 17280 1768 17332
rect 1820 17320 1826 17332
rect 2133 17323 2191 17329
rect 2133 17320 2145 17323
rect 1820 17292 2145 17320
rect 1820 17280 1826 17292
rect 2133 17289 2145 17292
rect 2179 17289 2191 17323
rect 2590 17320 2596 17332
rect 2551 17292 2596 17320
rect 2133 17283 2191 17289
rect 2590 17280 2596 17292
rect 2648 17280 2654 17332
rect 2682 17280 2688 17332
rect 2740 17320 2746 17332
rect 2869 17323 2927 17329
rect 2869 17320 2881 17323
rect 2740 17292 2881 17320
rect 2740 17280 2746 17292
rect 2869 17289 2881 17292
rect 2915 17289 2927 17323
rect 2869 17283 2927 17289
rect 3237 17323 3295 17329
rect 3237 17289 3249 17323
rect 3283 17289 3295 17323
rect 4430 17320 4436 17332
rect 4391 17292 4436 17320
rect 3237 17283 3295 17289
rect 3252 17252 3280 17283
rect 4430 17280 4436 17292
rect 4488 17280 4494 17332
rect 4890 17320 4896 17332
rect 4851 17292 4896 17320
rect 4890 17280 4896 17292
rect 4948 17280 4954 17332
rect 5445 17323 5503 17329
rect 5445 17289 5457 17323
rect 5491 17320 5503 17323
rect 5810 17320 5816 17332
rect 5491 17292 5816 17320
rect 5491 17289 5503 17292
rect 5445 17283 5503 17289
rect 5810 17280 5816 17292
rect 5868 17280 5874 17332
rect 5905 17323 5963 17329
rect 5905 17289 5917 17323
rect 5951 17320 5963 17323
rect 6917 17323 6975 17329
rect 6917 17320 6929 17323
rect 5951 17292 6929 17320
rect 5951 17289 5963 17292
rect 5905 17283 5963 17289
rect 6917 17289 6929 17292
rect 6963 17289 6975 17323
rect 7374 17320 7380 17332
rect 7335 17292 7380 17320
rect 6917 17283 6975 17289
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 7926 17320 7932 17332
rect 7887 17292 7932 17320
rect 7926 17280 7932 17292
rect 7984 17280 7990 17332
rect 8018 17280 8024 17332
rect 8076 17320 8082 17332
rect 8297 17323 8355 17329
rect 8297 17320 8309 17323
rect 8076 17292 8309 17320
rect 8076 17280 8082 17292
rect 8297 17289 8309 17292
rect 8343 17289 8355 17323
rect 8297 17283 8355 17289
rect 8478 17280 8484 17332
rect 8536 17320 8542 17332
rect 8665 17323 8723 17329
rect 8665 17320 8677 17323
rect 8536 17292 8677 17320
rect 8536 17280 8542 17292
rect 8665 17289 8677 17292
rect 8711 17289 8723 17323
rect 9122 17320 9128 17332
rect 9083 17292 9128 17320
rect 8665 17283 8723 17289
rect 9122 17280 9128 17292
rect 9180 17280 9186 17332
rect 9217 17323 9275 17329
rect 9217 17289 9229 17323
rect 9263 17320 9275 17323
rect 9585 17323 9643 17329
rect 9585 17320 9597 17323
rect 9263 17292 9597 17320
rect 9263 17289 9275 17292
rect 9217 17283 9275 17289
rect 9585 17289 9597 17292
rect 9631 17289 9643 17323
rect 10042 17320 10048 17332
rect 10003 17292 10048 17320
rect 9585 17283 9643 17289
rect 10042 17280 10048 17292
rect 10100 17280 10106 17332
rect 12802 17320 12808 17332
rect 10152 17292 12808 17320
rect 2792 17224 3280 17252
rect 1670 17184 1676 17196
rect 1631 17156 1676 17184
rect 1670 17144 1676 17156
rect 1728 17144 1734 17196
rect 2792 17193 2820 17224
rect 4154 17212 4160 17264
rect 4212 17252 4218 17264
rect 4525 17255 4583 17261
rect 4525 17252 4537 17255
rect 4212 17224 4537 17252
rect 4212 17212 4218 17224
rect 4525 17221 4537 17224
rect 4571 17252 4583 17255
rect 4614 17252 4620 17264
rect 4571 17224 4620 17252
rect 4571 17221 4583 17224
rect 4525 17215 4583 17221
rect 4614 17212 4620 17224
rect 4672 17212 4678 17264
rect 5718 17212 5724 17264
rect 5776 17252 5782 17264
rect 7009 17255 7067 17261
rect 7009 17252 7021 17255
rect 5776 17224 7021 17252
rect 5776 17212 5782 17224
rect 7009 17221 7021 17224
rect 7055 17221 7067 17255
rect 7834 17252 7840 17264
rect 7795 17224 7840 17252
rect 7009 17215 7067 17221
rect 7834 17212 7840 17224
rect 7892 17212 7898 17264
rect 8110 17212 8116 17264
rect 8168 17252 8174 17264
rect 10152 17252 10180 17292
rect 12802 17280 12808 17292
rect 12860 17280 12866 17332
rect 13170 17280 13176 17332
rect 13228 17280 13234 17332
rect 13464 17292 14596 17320
rect 12434 17252 12440 17264
rect 8168 17224 10180 17252
rect 10244 17224 12440 17252
rect 8168 17212 8174 17224
rect 2317 17187 2375 17193
rect 2317 17153 2329 17187
rect 2363 17153 2375 17187
rect 2317 17147 2375 17153
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17153 2835 17187
rect 3050 17184 3056 17196
rect 3011 17156 3056 17184
rect 2777 17147 2835 17153
rect 2332 17116 2360 17147
rect 3050 17144 3056 17156
rect 3108 17144 3114 17196
rect 3421 17187 3479 17193
rect 3421 17153 3433 17187
rect 3467 17153 3479 17187
rect 3421 17147 3479 17153
rect 2958 17116 2964 17128
rect 2332 17088 2964 17116
rect 2958 17076 2964 17088
rect 3016 17076 3022 17128
rect 3436 17116 3464 17147
rect 3510 17144 3516 17196
rect 3568 17184 3574 17196
rect 3697 17187 3755 17193
rect 3697 17184 3709 17187
rect 3568 17156 3709 17184
rect 3568 17144 3574 17156
rect 3697 17153 3709 17156
rect 3743 17153 3755 17187
rect 3697 17147 3755 17153
rect 4706 17144 4712 17196
rect 4764 17184 4770 17196
rect 5537 17187 5595 17193
rect 5537 17184 5549 17187
rect 4764 17156 5549 17184
rect 4764 17144 4770 17156
rect 5537 17153 5549 17156
rect 5583 17153 5595 17187
rect 8478 17184 8484 17196
rect 8439 17156 8484 17184
rect 5537 17147 5595 17153
rect 8478 17144 8484 17156
rect 8536 17144 8542 17196
rect 9950 17184 9956 17196
rect 9911 17156 9956 17184
rect 9950 17144 9956 17156
rect 10008 17144 10014 17196
rect 4341 17119 4399 17125
rect 3436 17088 3648 17116
rect 3513 17051 3571 17057
rect 3513 17048 3525 17051
rect 2746 17020 3525 17048
rect 1486 16980 1492 16992
rect 1447 16952 1492 16980
rect 1486 16940 1492 16952
rect 1544 16940 1550 16992
rect 1578 16940 1584 16992
rect 1636 16980 1642 16992
rect 2746 16980 2774 17020
rect 3513 17017 3525 17020
rect 3559 17017 3571 17051
rect 3620 17048 3648 17088
rect 4341 17085 4353 17119
rect 4387 17116 4399 17119
rect 4430 17116 4436 17128
rect 4387 17088 4436 17116
rect 4387 17085 4399 17088
rect 4341 17079 4399 17085
rect 4430 17076 4436 17088
rect 4488 17076 4494 17128
rect 5166 17076 5172 17128
rect 5224 17116 5230 17128
rect 5261 17119 5319 17125
rect 5261 17116 5273 17119
rect 5224 17088 5273 17116
rect 5224 17076 5230 17088
rect 5261 17085 5273 17088
rect 5307 17116 5319 17119
rect 5718 17116 5724 17128
rect 5307 17088 5724 17116
rect 5307 17085 5319 17088
rect 5261 17079 5319 17085
rect 5718 17076 5724 17088
rect 5776 17076 5782 17128
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17116 6883 17119
rect 6914 17116 6920 17128
rect 6871 17088 6920 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 6914 17076 6920 17088
rect 6972 17076 6978 17128
rect 7742 17116 7748 17128
rect 7703 17088 7748 17116
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 9398 17116 9404 17128
rect 9359 17088 9404 17116
rect 9398 17076 9404 17088
rect 9456 17076 9462 17128
rect 10244 17125 10272 17224
rect 12434 17212 12440 17224
rect 12492 17212 12498 17264
rect 12652 17255 12710 17261
rect 12652 17252 12664 17255
rect 12544 17224 12664 17252
rect 12544 17184 12572 17224
rect 12652 17221 12664 17224
rect 12698 17252 12710 17255
rect 13188 17252 13216 17280
rect 13262 17261 13268 17264
rect 12698 17224 13216 17252
rect 12698 17221 12710 17224
rect 12652 17215 12710 17221
rect 13256 17215 13268 17261
rect 13320 17252 13326 17264
rect 13320 17224 13356 17252
rect 13262 17212 13268 17215
rect 13320 17212 13326 17224
rect 10428 17156 12572 17184
rect 12897 17187 12955 17193
rect 10229 17119 10287 17125
rect 10229 17085 10241 17119
rect 10275 17085 10287 17119
rect 10229 17079 10287 17085
rect 8757 17051 8815 17057
rect 8757 17048 8769 17051
rect 3620 17020 8769 17048
rect 3513 17011 3571 17017
rect 8757 17017 8769 17020
rect 8803 17017 8815 17051
rect 8757 17011 8815 17017
rect 1636 16952 2774 16980
rect 1636 16940 1642 16952
rect 9674 16940 9680 16992
rect 9732 16980 9738 16992
rect 10428 16989 10456 17156
rect 12897 17153 12909 17187
rect 12943 17184 12955 17187
rect 12986 17184 12992 17196
rect 12943 17156 12992 17184
rect 12943 17153 12955 17156
rect 12897 17147 12955 17153
rect 12986 17144 12992 17156
rect 13044 17144 13050 17196
rect 13464 17184 13492 17292
rect 13722 17212 13728 17264
rect 13780 17252 13786 17264
rect 14461 17255 14519 17261
rect 14461 17252 14473 17255
rect 13780 17224 14473 17252
rect 13780 17212 13786 17224
rect 14461 17221 14473 17224
rect 14507 17221 14519 17255
rect 14568 17252 14596 17292
rect 14642 17280 14648 17332
rect 14700 17320 14706 17332
rect 15105 17323 15163 17329
rect 15105 17320 15117 17323
rect 14700 17292 15117 17320
rect 14700 17280 14706 17292
rect 15105 17289 15117 17292
rect 15151 17289 15163 17323
rect 15105 17283 15163 17289
rect 15212 17292 17071 17320
rect 15212 17252 15240 17292
rect 14568 17224 15240 17252
rect 14461 17215 14519 17221
rect 16206 17212 16212 17264
rect 16264 17261 16270 17264
rect 16264 17252 16276 17261
rect 16264 17224 16309 17252
rect 16264 17215 16276 17224
rect 16264 17212 16270 17215
rect 13096 17156 13492 17184
rect 13096 17116 13124 17156
rect 14366 17144 14372 17196
rect 14424 17184 14430 17196
rect 14642 17184 14648 17196
rect 14424 17156 14648 17184
rect 14424 17144 14430 17156
rect 14642 17144 14648 17156
rect 14700 17184 14706 17196
rect 16942 17184 16948 17196
rect 14700 17156 16948 17184
rect 14700 17144 14706 17156
rect 16942 17144 16948 17156
rect 17000 17144 17006 17196
rect 17043 17184 17071 17292
rect 17862 17280 17868 17332
rect 17920 17320 17926 17332
rect 18141 17323 18199 17329
rect 18141 17320 18153 17323
rect 17920 17292 18153 17320
rect 17920 17280 17926 17292
rect 18064 17193 18092 17292
rect 18141 17289 18153 17292
rect 18187 17289 18199 17323
rect 18141 17283 18199 17289
rect 20441 17255 20499 17261
rect 20441 17252 20453 17255
rect 18984 17224 20453 17252
rect 18984 17193 19012 17224
rect 20441 17221 20453 17224
rect 20487 17252 20499 17255
rect 21269 17255 21327 17261
rect 21269 17252 21281 17255
rect 20487 17224 21281 17252
rect 20487 17221 20499 17224
rect 20441 17215 20499 17221
rect 21269 17221 21281 17224
rect 21315 17221 21327 17255
rect 21269 17215 21327 17221
rect 17793 17187 17851 17193
rect 17793 17184 17805 17187
rect 17043 17156 17805 17184
rect 17793 17153 17805 17156
rect 17839 17184 17851 17187
rect 18049 17187 18107 17193
rect 17839 17156 18000 17184
rect 17839 17153 17851 17156
rect 17793 17147 17851 17153
rect 16482 17116 16488 17128
rect 12912 17088 13124 17116
rect 16443 17088 16488 17116
rect 11517 17051 11575 17057
rect 11517 17017 11529 17051
rect 11563 17048 11575 17051
rect 11790 17048 11796 17060
rect 11563 17020 11796 17048
rect 11563 17017 11575 17020
rect 11517 17011 11575 17017
rect 11790 17008 11796 17020
rect 11848 17008 11854 17060
rect 10413 16983 10471 16989
rect 10413 16980 10425 16983
rect 9732 16952 10425 16980
rect 9732 16940 9738 16952
rect 10413 16949 10425 16952
rect 10459 16949 10471 16983
rect 10413 16943 10471 16949
rect 11606 16940 11612 16992
rect 11664 16980 11670 16992
rect 12912 16980 12940 17088
rect 16482 17076 16488 17088
rect 16540 17076 16546 17128
rect 17972 17116 18000 17156
rect 18049 17153 18061 17187
rect 18095 17184 18107 17187
rect 18969 17187 19027 17193
rect 18969 17184 18981 17187
rect 18095 17156 18981 17184
rect 18095 17153 18107 17156
rect 18049 17147 18107 17153
rect 18969 17153 18981 17156
rect 19015 17153 19027 17187
rect 19225 17187 19283 17193
rect 19225 17184 19237 17187
rect 18969 17147 19027 17153
rect 19076 17156 19237 17184
rect 17972 17088 18092 17116
rect 14292 17020 15608 17048
rect 11664 16952 12940 16980
rect 11664 16940 11670 16952
rect 13170 16940 13176 16992
rect 13228 16980 13234 16992
rect 14292 16980 14320 17020
rect 13228 16952 14320 16980
rect 13228 16940 13234 16952
rect 14366 16940 14372 16992
rect 14424 16980 14430 16992
rect 15580 16980 15608 17020
rect 16669 16983 16727 16989
rect 16669 16980 16681 16983
rect 14424 16952 14469 16980
rect 15580 16952 16681 16980
rect 14424 16940 14430 16952
rect 16669 16949 16681 16952
rect 16715 16980 16727 16983
rect 17402 16980 17408 16992
rect 16715 16952 17408 16980
rect 16715 16949 16727 16952
rect 16669 16943 16727 16949
rect 17402 16940 17408 16952
rect 17460 16940 17466 16992
rect 18064 16980 18092 17088
rect 18138 17076 18144 17128
rect 18196 17116 18202 17128
rect 19076 17116 19104 17156
rect 19225 17153 19237 17156
rect 19271 17153 19283 17187
rect 19225 17147 19283 17153
rect 18196 17088 19104 17116
rect 18196 17076 18202 17088
rect 20162 16980 20168 16992
rect 18064 16952 20168 16980
rect 20162 16940 20168 16952
rect 20220 16940 20226 16992
rect 20346 16980 20352 16992
rect 20307 16952 20352 16980
rect 20346 16940 20352 16952
rect 20404 16940 20410 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 2958 16776 2964 16788
rect 2919 16748 2964 16776
rect 2958 16736 2964 16748
rect 3016 16736 3022 16788
rect 3418 16776 3424 16788
rect 3379 16748 3424 16776
rect 3418 16736 3424 16748
rect 3476 16736 3482 16788
rect 4706 16776 4712 16788
rect 4667 16748 4712 16776
rect 4706 16736 4712 16748
rect 4764 16736 4770 16788
rect 5350 16736 5356 16788
rect 5408 16776 5414 16788
rect 8110 16776 8116 16788
rect 5408 16748 8116 16776
rect 5408 16736 5414 16748
rect 8110 16736 8116 16748
rect 8168 16736 8174 16788
rect 12342 16736 12348 16788
rect 12400 16736 12406 16788
rect 12526 16736 12532 16788
rect 12584 16776 12590 16788
rect 12986 16776 12992 16788
rect 12584 16748 12992 16776
rect 12584 16736 12590 16748
rect 12986 16736 12992 16748
rect 13044 16776 13050 16788
rect 13044 16748 13308 16776
rect 13044 16736 13050 16748
rect 4430 16708 4436 16720
rect 4080 16680 4436 16708
rect 4080 16649 4108 16680
rect 4430 16668 4436 16680
rect 4488 16708 4494 16720
rect 4982 16708 4988 16720
rect 4488 16680 4988 16708
rect 4488 16668 4494 16680
rect 4982 16668 4988 16680
rect 5040 16668 5046 16720
rect 12360 16708 12388 16736
rect 7760 16680 12388 16708
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16609 4123 16643
rect 4246 16640 4252 16652
rect 4207 16612 4252 16640
rect 4065 16603 4123 16609
rect 4246 16600 4252 16612
rect 4304 16640 4310 16652
rect 6178 16640 6184 16652
rect 4304 16612 4660 16640
rect 6139 16612 6184 16640
rect 4304 16600 4310 16612
rect 4632 16584 4660 16612
rect 6178 16600 6184 16612
rect 6236 16600 6242 16652
rect 7558 16640 7564 16652
rect 7519 16612 7564 16640
rect 7558 16600 7564 16612
rect 7616 16600 7622 16652
rect 7760 16649 7788 16680
rect 7745 16643 7803 16649
rect 7745 16609 7757 16643
rect 7791 16609 7803 16643
rect 8110 16640 8116 16652
rect 8071 16612 8116 16640
rect 7745 16603 7803 16609
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 8386 16600 8392 16652
rect 8444 16640 8450 16652
rect 9674 16640 9680 16652
rect 8444 16612 8984 16640
rect 9635 16612 9680 16640
rect 8444 16600 8450 16612
rect 1578 16532 1584 16584
rect 1636 16572 1642 16584
rect 1673 16575 1731 16581
rect 1673 16572 1685 16575
rect 1636 16544 1685 16572
rect 1636 16532 1642 16544
rect 1673 16541 1685 16544
rect 1719 16541 1731 16575
rect 2038 16572 2044 16584
rect 1999 16544 2044 16572
rect 1673 16535 1731 16541
rect 2038 16532 2044 16544
rect 2096 16532 2102 16584
rect 3145 16575 3203 16581
rect 3145 16541 3157 16575
rect 3191 16541 3203 16575
rect 3145 16535 3203 16541
rect 3237 16575 3295 16581
rect 3237 16541 3249 16575
rect 3283 16572 3295 16575
rect 4154 16572 4160 16584
rect 3283 16544 4160 16572
rect 3283 16541 3295 16544
rect 3237 16535 3295 16541
rect 3160 16504 3188 16535
rect 4154 16532 4160 16544
rect 4212 16532 4218 16584
rect 4338 16572 4344 16584
rect 4299 16544 4344 16572
rect 4338 16532 4344 16544
rect 4396 16532 4402 16584
rect 4614 16532 4620 16584
rect 4672 16532 4678 16584
rect 8202 16532 8208 16584
rect 8260 16572 8266 16584
rect 8297 16575 8355 16581
rect 8297 16572 8309 16575
rect 8260 16544 8309 16572
rect 8260 16532 8266 16544
rect 8297 16541 8309 16544
rect 8343 16541 8355 16575
rect 8297 16535 8355 16541
rect 7009 16507 7067 16513
rect 3160 16476 6224 16504
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 1854 16436 1860 16448
rect 1815 16408 1860 16436
rect 1854 16396 1860 16408
rect 1912 16396 1918 16448
rect 3142 16396 3148 16448
rect 3200 16436 3206 16448
rect 5537 16439 5595 16445
rect 5537 16436 5549 16439
rect 3200 16408 5549 16436
rect 3200 16396 3206 16408
rect 5537 16405 5549 16408
rect 5583 16405 5595 16439
rect 5902 16436 5908 16448
rect 5863 16408 5908 16436
rect 5537 16399 5595 16405
rect 5902 16396 5908 16408
rect 5960 16396 5966 16448
rect 5994 16396 6000 16448
rect 6052 16436 6058 16448
rect 6196 16436 6224 16476
rect 7009 16473 7021 16507
rect 7055 16504 7067 16507
rect 7469 16507 7527 16513
rect 7469 16504 7481 16507
rect 7055 16476 7481 16504
rect 7055 16473 7067 16476
rect 7009 16467 7067 16473
rect 7469 16473 7481 16476
rect 7515 16473 7527 16507
rect 7469 16467 7527 16473
rect 7101 16439 7159 16445
rect 7101 16436 7113 16439
rect 6052 16408 6097 16436
rect 6196 16408 7113 16436
rect 6052 16396 6058 16408
rect 7101 16405 7113 16408
rect 7147 16405 7159 16439
rect 7101 16399 7159 16405
rect 8110 16396 8116 16448
rect 8168 16436 8174 16448
rect 8205 16439 8263 16445
rect 8205 16436 8217 16439
rect 8168 16408 8217 16436
rect 8168 16396 8174 16408
rect 8205 16405 8217 16408
rect 8251 16405 8263 16439
rect 8662 16436 8668 16448
rect 8623 16408 8668 16436
rect 8205 16399 8263 16405
rect 8662 16396 8668 16408
rect 8720 16396 8726 16448
rect 8956 16436 8984 16612
rect 9674 16600 9680 16612
rect 9732 16600 9738 16652
rect 10410 16640 10416 16652
rect 9784 16612 10416 16640
rect 9214 16572 9220 16584
rect 9175 16544 9220 16572
rect 9214 16532 9220 16544
rect 9272 16532 9278 16584
rect 9493 16575 9551 16581
rect 9493 16541 9505 16575
rect 9539 16572 9551 16575
rect 9582 16572 9588 16584
rect 9539 16544 9588 16572
rect 9539 16541 9551 16544
rect 9493 16535 9551 16541
rect 9582 16532 9588 16544
rect 9640 16532 9646 16584
rect 9122 16464 9128 16516
rect 9180 16504 9186 16516
rect 9784 16504 9812 16612
rect 10410 16600 10416 16612
rect 10468 16600 10474 16652
rect 10965 16643 11023 16649
rect 10965 16609 10977 16643
rect 11011 16640 11023 16643
rect 11606 16640 11612 16652
rect 11011 16612 11612 16640
rect 11011 16609 11023 16612
rect 10965 16603 11023 16609
rect 11606 16600 11612 16612
rect 11664 16600 11670 16652
rect 13280 16649 13308 16748
rect 15470 16736 15476 16788
rect 15528 16776 15534 16788
rect 16025 16779 16083 16785
rect 16025 16776 16037 16779
rect 15528 16748 16037 16776
rect 15528 16736 15534 16748
rect 16025 16745 16037 16748
rect 16071 16776 16083 16779
rect 16206 16776 16212 16788
rect 16071 16748 16212 16776
rect 16071 16745 16083 16748
rect 16025 16739 16083 16745
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 17954 16736 17960 16788
rect 18012 16776 18018 16788
rect 18417 16779 18475 16785
rect 18417 16776 18429 16779
rect 18012 16748 18429 16776
rect 18012 16736 18018 16748
rect 13265 16643 13323 16649
rect 13265 16609 13277 16643
rect 13311 16640 13323 16643
rect 13630 16640 13636 16652
rect 13311 16612 13636 16640
rect 13311 16609 13323 16612
rect 13265 16603 13323 16609
rect 13630 16600 13636 16612
rect 13688 16600 13694 16652
rect 18340 16649 18368 16748
rect 18417 16745 18429 16748
rect 18463 16745 18475 16779
rect 18417 16739 18475 16745
rect 18325 16643 18383 16649
rect 18325 16609 18337 16643
rect 18371 16640 18383 16643
rect 19334 16640 19340 16652
rect 18371 16612 19340 16640
rect 18371 16609 18383 16612
rect 18325 16603 18383 16609
rect 19334 16600 19340 16612
rect 19392 16600 19398 16652
rect 9953 16575 10011 16581
rect 9953 16541 9965 16575
rect 9999 16572 10011 16575
rect 10226 16572 10232 16584
rect 9999 16544 10232 16572
rect 9999 16541 10011 16544
rect 9953 16535 10011 16541
rect 10226 16532 10232 16544
rect 10284 16572 10290 16584
rect 11241 16575 11299 16581
rect 11241 16572 11253 16575
rect 10284 16544 11253 16572
rect 10284 16532 10290 16544
rect 11241 16541 11253 16544
rect 11287 16541 11299 16575
rect 11241 16535 11299 16541
rect 11882 16532 11888 16584
rect 11940 16572 11946 16584
rect 13009 16575 13067 16581
rect 13009 16572 13021 16575
rect 11940 16544 13021 16572
rect 11940 16532 11946 16544
rect 13009 16541 13021 16544
rect 13055 16572 13067 16575
rect 13541 16575 13599 16581
rect 13541 16572 13553 16575
rect 13055 16544 13553 16572
rect 13055 16541 13067 16544
rect 13009 16535 13067 16541
rect 13541 16541 13553 16544
rect 13587 16572 13599 16575
rect 15746 16572 15752 16584
rect 13587 16544 15608 16572
rect 15707 16544 15752 16572
rect 13587 16541 13599 16544
rect 13541 16535 13599 16541
rect 9180 16476 9812 16504
rect 9180 16464 9186 16476
rect 10042 16464 10048 16516
rect 10100 16504 10106 16516
rect 10100 16476 10456 16504
rect 10100 16464 10106 16476
rect 9033 16439 9091 16445
rect 9033 16436 9045 16439
rect 8956 16408 9045 16436
rect 9033 16405 9045 16408
rect 9079 16405 9091 16439
rect 9306 16436 9312 16448
rect 9267 16408 9312 16436
rect 9033 16399 9091 16405
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 9398 16396 9404 16448
rect 9456 16436 9462 16448
rect 9861 16439 9919 16445
rect 9861 16436 9873 16439
rect 9456 16408 9873 16436
rect 9456 16396 9462 16408
rect 9861 16405 9873 16408
rect 9907 16405 9919 16439
rect 10318 16436 10324 16448
rect 10279 16408 10324 16436
rect 9861 16399 9919 16405
rect 10318 16396 10324 16408
rect 10376 16396 10382 16448
rect 10428 16445 10456 16476
rect 12894 16464 12900 16516
rect 12952 16504 12958 16516
rect 15470 16504 15476 16516
rect 15528 16513 15534 16516
rect 12952 16476 15476 16504
rect 12952 16464 12958 16476
rect 15470 16464 15476 16476
rect 15528 16467 15540 16513
rect 15580 16504 15608 16544
rect 15746 16532 15752 16544
rect 15804 16572 15810 16584
rect 16482 16572 16488 16584
rect 15804 16544 16488 16572
rect 15804 16532 15810 16544
rect 16482 16532 16488 16544
rect 16540 16572 16546 16584
rect 16577 16575 16635 16581
rect 16577 16572 16589 16575
rect 16540 16544 16589 16572
rect 16540 16532 16546 16544
rect 16577 16541 16589 16544
rect 16623 16541 16635 16575
rect 19352 16572 19380 16600
rect 20625 16575 20683 16581
rect 20625 16572 20637 16575
rect 19352 16544 20637 16572
rect 16577 16535 16635 16541
rect 20625 16541 20637 16544
rect 20671 16572 20683 16575
rect 20717 16575 20775 16581
rect 20717 16572 20729 16575
rect 20671 16544 20729 16572
rect 20671 16541 20683 16544
rect 20625 16535 20683 16541
rect 20717 16541 20729 16544
rect 20763 16572 20775 16575
rect 21450 16572 21456 16584
rect 20763 16544 21456 16572
rect 20763 16541 20775 16544
rect 20717 16535 20775 16541
rect 21450 16532 21456 16544
rect 21508 16532 21514 16584
rect 15580 16476 16988 16504
rect 15528 16464 15534 16467
rect 10413 16439 10471 16445
rect 10413 16405 10425 16439
rect 10459 16405 10471 16439
rect 10778 16436 10784 16448
rect 10739 16408 10784 16436
rect 10413 16399 10471 16405
rect 10778 16396 10784 16408
rect 10836 16396 10842 16448
rect 10873 16439 10931 16445
rect 10873 16405 10885 16439
rect 10919 16436 10931 16439
rect 11054 16436 11060 16448
rect 10919 16408 11060 16436
rect 10919 16405 10931 16408
rect 10873 16399 10931 16405
rect 11054 16396 11060 16408
rect 11112 16396 11118 16448
rect 11885 16439 11943 16445
rect 11885 16405 11897 16439
rect 11931 16436 11943 16439
rect 12526 16436 12532 16448
rect 11931 16408 12532 16436
rect 11931 16405 11943 16408
rect 11885 16399 11943 16405
rect 12526 16396 12532 16408
rect 12584 16396 12590 16448
rect 13449 16439 13507 16445
rect 13449 16405 13461 16439
rect 13495 16436 13507 16439
rect 13630 16436 13636 16448
rect 13495 16408 13636 16436
rect 13495 16405 13507 16408
rect 13449 16399 13507 16405
rect 13630 16396 13636 16408
rect 13688 16396 13694 16448
rect 14274 16396 14280 16448
rect 14332 16436 14338 16448
rect 14369 16439 14427 16445
rect 14369 16436 14381 16439
rect 14332 16408 14381 16436
rect 14332 16396 14338 16408
rect 14369 16405 14381 16408
rect 14415 16405 14427 16439
rect 14369 16399 14427 16405
rect 15194 16396 15200 16448
rect 15252 16436 15258 16448
rect 15746 16436 15752 16448
rect 15252 16408 15752 16436
rect 15252 16396 15258 16408
rect 15746 16396 15752 16408
rect 15804 16436 15810 16448
rect 16960 16445 16988 16476
rect 17954 16464 17960 16516
rect 18012 16504 18018 16516
rect 18058 16507 18116 16513
rect 18058 16504 18070 16507
rect 18012 16476 18070 16504
rect 18012 16464 18018 16476
rect 18058 16473 18070 16476
rect 18104 16473 18116 16507
rect 18058 16467 18116 16473
rect 18230 16464 18236 16516
rect 18288 16504 18294 16516
rect 20358 16507 20416 16513
rect 20358 16504 20370 16507
rect 18288 16476 20370 16504
rect 18288 16464 18294 16476
rect 20358 16473 20370 16476
rect 20404 16473 20416 16507
rect 20358 16467 20416 16473
rect 15841 16439 15899 16445
rect 15841 16436 15853 16439
rect 15804 16408 15853 16436
rect 15804 16396 15810 16408
rect 15841 16405 15853 16408
rect 15887 16405 15899 16439
rect 15841 16399 15899 16405
rect 16945 16439 17003 16445
rect 16945 16405 16957 16439
rect 16991 16405 17003 16439
rect 16945 16399 17003 16405
rect 19058 16396 19064 16448
rect 19116 16436 19122 16448
rect 19245 16439 19303 16445
rect 19245 16436 19257 16439
rect 19116 16408 19257 16436
rect 19116 16396 19122 16408
rect 19245 16405 19257 16408
rect 19291 16405 19303 16439
rect 19245 16399 19303 16405
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 2866 16192 2872 16244
rect 2924 16232 2930 16244
rect 2961 16235 3019 16241
rect 2961 16232 2973 16235
rect 2924 16204 2973 16232
rect 2924 16192 2930 16204
rect 2961 16201 2973 16204
rect 3007 16201 3019 16235
rect 2961 16195 3019 16201
rect 3050 16192 3056 16244
rect 3108 16232 3114 16244
rect 3421 16235 3479 16241
rect 3421 16232 3433 16235
rect 3108 16204 3433 16232
rect 3108 16192 3114 16204
rect 3421 16201 3433 16204
rect 3467 16201 3479 16235
rect 3421 16195 3479 16201
rect 5261 16235 5319 16241
rect 5261 16201 5273 16235
rect 5307 16232 5319 16235
rect 5902 16232 5908 16244
rect 5307 16204 5908 16232
rect 5307 16201 5319 16204
rect 5261 16195 5319 16201
rect 5902 16192 5908 16204
rect 5960 16192 5966 16244
rect 6089 16235 6147 16241
rect 6089 16201 6101 16235
rect 6135 16232 6147 16235
rect 7745 16235 7803 16241
rect 7745 16232 7757 16235
rect 6135 16204 7757 16232
rect 6135 16201 6147 16204
rect 6089 16195 6147 16201
rect 7745 16201 7757 16204
rect 7791 16201 7803 16235
rect 8386 16232 8392 16244
rect 8347 16204 8392 16232
rect 7745 16195 7803 16201
rect 8386 16192 8392 16204
rect 8444 16192 8450 16244
rect 8754 16192 8760 16244
rect 8812 16232 8818 16244
rect 9306 16232 9312 16244
rect 8812 16204 9312 16232
rect 8812 16192 8818 16204
rect 9306 16192 9312 16204
rect 9364 16192 9370 16244
rect 9766 16232 9772 16244
rect 9727 16204 9772 16232
rect 9766 16192 9772 16204
rect 9824 16192 9830 16244
rect 10597 16235 10655 16241
rect 9968 16204 10548 16232
rect 6362 16164 6368 16176
rect 5368 16136 6368 16164
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16096 1731 16099
rect 2130 16096 2136 16108
rect 1719 16068 2136 16096
rect 1719 16065 1731 16068
rect 1673 16059 1731 16065
rect 2130 16056 2136 16068
rect 2188 16056 2194 16108
rect 3142 16096 3148 16108
rect 3103 16068 3148 16096
rect 3142 16056 3148 16068
rect 3200 16056 3206 16108
rect 3605 16099 3663 16105
rect 3605 16065 3617 16099
rect 3651 16096 3663 16099
rect 5074 16096 5080 16108
rect 3651 16068 5080 16096
rect 3651 16065 3663 16068
rect 3605 16059 3663 16065
rect 5074 16056 5080 16068
rect 5132 16056 5138 16108
rect 5368 16028 5396 16136
rect 6362 16124 6368 16136
rect 6420 16124 6426 16176
rect 6546 16124 6552 16176
rect 6604 16164 6610 16176
rect 6825 16167 6883 16173
rect 6825 16164 6837 16167
rect 6604 16136 6837 16164
rect 6604 16124 6610 16136
rect 6825 16133 6837 16136
rect 6871 16133 6883 16167
rect 6825 16127 6883 16133
rect 8110 16124 8116 16176
rect 8168 16164 8174 16176
rect 8849 16167 8907 16173
rect 8849 16164 8861 16167
rect 8168 16136 8861 16164
rect 8168 16124 8174 16136
rect 8849 16133 8861 16136
rect 8895 16164 8907 16167
rect 9122 16164 9128 16176
rect 8895 16136 9128 16164
rect 8895 16133 8907 16136
rect 8849 16127 8907 16133
rect 9122 16124 9128 16136
rect 9180 16124 9186 16176
rect 5721 16099 5779 16105
rect 5721 16096 5733 16099
rect 5552 16068 5733 16096
rect 5445 16031 5503 16037
rect 5445 16028 5457 16031
rect 5368 16000 5457 16028
rect 5445 15997 5457 16000
rect 5491 15997 5503 16031
rect 5445 15991 5503 15997
rect 5166 15920 5172 15972
rect 5224 15960 5230 15972
rect 5552 15960 5580 16068
rect 5721 16065 5733 16068
rect 5767 16065 5779 16099
rect 5721 16059 5779 16065
rect 5902 16056 5908 16108
rect 5960 16096 5966 16108
rect 6917 16099 6975 16105
rect 6917 16096 6929 16099
rect 5960 16068 6929 16096
rect 5960 16056 5966 16068
rect 6917 16065 6929 16068
rect 6963 16065 6975 16099
rect 7834 16096 7840 16108
rect 7795 16068 7840 16096
rect 6917 16059 6975 16065
rect 7834 16056 7840 16068
rect 7892 16056 7898 16108
rect 8570 16056 8576 16108
rect 8628 16096 8634 16108
rect 9398 16096 9404 16108
rect 8628 16068 9404 16096
rect 8628 16056 8634 16068
rect 5629 16031 5687 16037
rect 5629 15997 5641 16031
rect 5675 15997 5687 16031
rect 5629 15991 5687 15997
rect 6733 16031 6791 16037
rect 6733 15997 6745 16031
rect 6779 15997 6791 16031
rect 7653 16031 7711 16037
rect 7653 16028 7665 16031
rect 6733 15991 6791 15997
rect 7024 16000 7665 16028
rect 5224 15932 5580 15960
rect 5644 15960 5672 15991
rect 5994 15960 6000 15972
rect 5644 15932 6000 15960
rect 5224 15920 5230 15932
rect 5994 15920 6000 15932
rect 6052 15920 6058 15972
rect 6748 15960 6776 15991
rect 6914 15960 6920 15972
rect 6196 15932 6500 15960
rect 6748 15932 6920 15960
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 4890 15852 4896 15904
rect 4948 15892 4954 15904
rect 5350 15892 5356 15904
rect 4948 15864 5356 15892
rect 4948 15852 4954 15864
rect 5350 15852 5356 15864
rect 5408 15852 5414 15904
rect 5902 15852 5908 15904
rect 5960 15892 5966 15904
rect 6196 15892 6224 15932
rect 6362 15892 6368 15904
rect 5960 15864 6224 15892
rect 6323 15864 6368 15892
rect 5960 15852 5966 15864
rect 6362 15852 6368 15864
rect 6420 15852 6426 15904
rect 6472 15892 6500 15932
rect 6914 15920 6920 15932
rect 6972 15920 6978 15972
rect 7024 15892 7052 16000
rect 7653 15997 7665 16000
rect 7699 16028 7711 16031
rect 7742 16028 7748 16040
rect 7699 16000 7748 16028
rect 7699 15997 7711 16000
rect 7653 15991 7711 15997
rect 7742 15988 7748 16000
rect 7800 15988 7806 16040
rect 7285 15963 7343 15969
rect 7285 15929 7297 15963
rect 7331 15960 7343 15963
rect 8570 15960 8576 15972
rect 7331 15932 8576 15960
rect 7331 15929 7343 15932
rect 7285 15923 7343 15929
rect 8570 15920 8576 15932
rect 8628 15920 8634 15972
rect 6472 15864 7052 15892
rect 7926 15852 7932 15904
rect 7984 15892 7990 15904
rect 8205 15895 8263 15901
rect 8205 15892 8217 15895
rect 7984 15864 8217 15892
rect 7984 15852 7990 15864
rect 8205 15861 8217 15864
rect 8251 15861 8263 15895
rect 8205 15855 8263 15861
rect 8386 15852 8392 15904
rect 8444 15892 8450 15904
rect 9232 15901 9260 16068
rect 9398 16056 9404 16068
rect 9456 16056 9462 16108
rect 9585 16099 9643 16105
rect 9585 16065 9597 16099
rect 9631 16096 9643 16099
rect 9858 16096 9864 16108
rect 9631 16068 9864 16096
rect 9631 16065 9643 16068
rect 9585 16059 9643 16065
rect 9858 16056 9864 16068
rect 9916 16056 9922 16108
rect 9968 16096 9996 16204
rect 10520 16164 10548 16204
rect 10597 16201 10609 16235
rect 10643 16232 10655 16235
rect 10870 16232 10876 16244
rect 10643 16204 10876 16232
rect 10643 16201 10655 16204
rect 10597 16195 10655 16201
rect 10870 16192 10876 16204
rect 10928 16192 10934 16244
rect 11054 16232 11060 16244
rect 11015 16204 11060 16232
rect 11054 16192 11060 16204
rect 11112 16192 11118 16244
rect 11238 16192 11244 16244
rect 11296 16232 11302 16244
rect 11296 16204 13492 16232
rect 11296 16192 11302 16204
rect 10689 16167 10747 16173
rect 10689 16164 10701 16167
rect 10520 16136 10701 16164
rect 10689 16133 10701 16136
rect 10735 16133 10747 16167
rect 10689 16127 10747 16133
rect 10778 16124 10784 16176
rect 10836 16164 10842 16176
rect 11517 16167 11575 16173
rect 11517 16164 11529 16167
rect 10836 16136 11529 16164
rect 10836 16124 10842 16136
rect 11517 16133 11529 16136
rect 11563 16133 11575 16167
rect 11517 16127 11575 16133
rect 13078 16124 13084 16176
rect 13136 16164 13142 16176
rect 13274 16167 13332 16173
rect 13274 16164 13286 16167
rect 13136 16136 13286 16164
rect 13136 16124 13142 16136
rect 13274 16133 13286 16136
rect 13320 16133 13332 16167
rect 13274 16127 13332 16133
rect 12894 16096 12900 16108
rect 9968 16068 10088 16096
rect 9950 16028 9956 16040
rect 9911 16000 9956 16028
rect 9950 15988 9956 16000
rect 10008 15988 10014 16040
rect 10060 15960 10088 16068
rect 9646 15932 10088 15960
rect 10152 16068 12900 16096
rect 9217 15895 9275 15901
rect 9217 15892 9229 15895
rect 8444 15864 9229 15892
rect 8444 15852 8450 15864
rect 9217 15861 9229 15864
rect 9263 15861 9275 15895
rect 9398 15892 9404 15904
rect 9359 15864 9404 15892
rect 9217 15855 9275 15861
rect 9398 15852 9404 15864
rect 9456 15892 9462 15904
rect 9646 15892 9674 15932
rect 9456 15864 9674 15892
rect 9456 15852 9462 15864
rect 9766 15852 9772 15904
rect 9824 15892 9830 15904
rect 10152 15901 10180 16068
rect 12894 16056 12900 16068
rect 12952 16056 12958 16108
rect 10502 16028 10508 16040
rect 10463 16000 10508 16028
rect 10502 15988 10508 16000
rect 10560 15988 10566 16040
rect 11146 16028 11152 16040
rect 11107 16000 11152 16028
rect 11146 15988 11152 16000
rect 11204 15988 11210 16040
rect 13464 16028 13492 16204
rect 14918 16192 14924 16244
rect 14976 16232 14982 16244
rect 17957 16235 18015 16241
rect 17957 16232 17969 16235
rect 14976 16204 17969 16232
rect 14976 16192 14982 16204
rect 17957 16201 17969 16204
rect 18003 16201 18015 16235
rect 17957 16195 18015 16201
rect 15194 16164 15200 16176
rect 13648 16136 15200 16164
rect 13648 16108 13676 16136
rect 15194 16124 15200 16136
rect 15252 16164 15258 16176
rect 15289 16167 15347 16173
rect 15289 16164 15301 16167
rect 15252 16136 15301 16164
rect 15252 16124 15258 16136
rect 15289 16133 15301 16136
rect 15335 16133 15347 16167
rect 20070 16164 20076 16176
rect 15289 16127 15347 16133
rect 18340 16136 20076 16164
rect 13541 16099 13599 16105
rect 13541 16065 13553 16099
rect 13587 16096 13599 16099
rect 13630 16096 13636 16108
rect 13587 16068 13636 16096
rect 13587 16065 13599 16068
rect 13541 16059 13599 16065
rect 13630 16056 13636 16068
rect 13688 16056 13694 16108
rect 14941 16099 14999 16105
rect 14941 16065 14953 16099
rect 14987 16096 14999 16099
rect 15562 16096 15568 16108
rect 14987 16068 15568 16096
rect 14987 16065 14999 16068
rect 14941 16059 14999 16065
rect 15562 16056 15568 16068
rect 15620 16056 15626 16108
rect 15194 16028 15200 16040
rect 13464 16000 14228 16028
rect 15155 16000 15200 16028
rect 12158 15960 12164 15972
rect 12119 15932 12164 15960
rect 12158 15920 12164 15932
rect 12216 15920 12222 15972
rect 13817 15963 13875 15969
rect 13817 15960 13829 15963
rect 13556 15932 13829 15960
rect 10137 15895 10195 15901
rect 10137 15892 10149 15895
rect 9824 15864 10149 15892
rect 9824 15852 9830 15864
rect 10137 15861 10149 15864
rect 10183 15861 10195 15895
rect 10137 15855 10195 15861
rect 12434 15852 12440 15904
rect 12492 15892 12498 15904
rect 13556 15892 13584 15932
rect 13817 15929 13829 15932
rect 13863 15929 13875 15963
rect 13817 15923 13875 15929
rect 12492 15864 13584 15892
rect 14200 15892 14228 16000
rect 15194 15988 15200 16000
rect 15252 15988 15258 16040
rect 18340 15960 18368 16136
rect 20070 16124 20076 16136
rect 20128 16124 20134 16176
rect 19058 16056 19064 16108
rect 19116 16105 19122 16108
rect 19116 16096 19128 16105
rect 19334 16096 19340 16108
rect 19116 16068 19161 16096
rect 19295 16068 19340 16096
rect 19116 16059 19128 16068
rect 19116 16056 19122 16059
rect 19334 16056 19340 16068
rect 19392 16096 19398 16108
rect 19429 16099 19487 16105
rect 19429 16096 19441 16099
rect 19392 16068 19441 16096
rect 19392 16056 19398 16068
rect 19429 16065 19441 16068
rect 19475 16065 19487 16099
rect 21174 16096 21180 16108
rect 21232 16105 21238 16108
rect 21144 16068 21180 16096
rect 19429 16059 19487 16065
rect 21174 16056 21180 16068
rect 21232 16059 21244 16105
rect 21450 16096 21456 16108
rect 21411 16068 21456 16096
rect 21232 16056 21238 16059
rect 21450 16056 21456 16068
rect 21508 16056 21514 16108
rect 15488 15932 18368 15960
rect 15488 15892 15516 15932
rect 14200 15864 15516 15892
rect 12492 15852 12498 15864
rect 15562 15852 15568 15904
rect 15620 15892 15626 15904
rect 16022 15892 16028 15904
rect 15620 15864 16028 15892
rect 15620 15852 15626 15864
rect 16022 15852 16028 15864
rect 16080 15852 16086 15904
rect 16390 15852 16396 15904
rect 16448 15892 16454 15904
rect 20073 15895 20131 15901
rect 20073 15892 20085 15895
rect 16448 15864 20085 15892
rect 16448 15852 16454 15864
rect 20073 15861 20085 15864
rect 20119 15861 20131 15895
rect 20073 15855 20131 15861
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 1670 15648 1676 15700
rect 1728 15688 1734 15700
rect 1857 15691 1915 15697
rect 1857 15688 1869 15691
rect 1728 15660 1869 15688
rect 1728 15648 1734 15660
rect 1857 15657 1869 15660
rect 1903 15657 1915 15691
rect 1857 15651 1915 15657
rect 1946 15648 1952 15700
rect 2004 15688 2010 15700
rect 2225 15691 2283 15697
rect 2225 15688 2237 15691
rect 2004 15660 2237 15688
rect 2004 15648 2010 15660
rect 2225 15657 2237 15660
rect 2271 15657 2283 15691
rect 2498 15688 2504 15700
rect 2459 15660 2504 15688
rect 2225 15651 2283 15657
rect 2498 15648 2504 15660
rect 2556 15648 2562 15700
rect 5166 15688 5172 15700
rect 5127 15660 5172 15688
rect 5166 15648 5172 15660
rect 5224 15648 5230 15700
rect 5994 15688 6000 15700
rect 5955 15660 6000 15688
rect 5994 15648 6000 15660
rect 6052 15648 6058 15700
rect 6086 15648 6092 15700
rect 6144 15688 6150 15700
rect 6144 15660 6189 15688
rect 6144 15648 6150 15660
rect 7834 15648 7840 15700
rect 7892 15688 7898 15700
rect 8941 15691 8999 15697
rect 8941 15688 8953 15691
rect 7892 15660 8953 15688
rect 7892 15648 7898 15660
rect 8941 15657 8953 15660
rect 8987 15657 8999 15691
rect 9766 15688 9772 15700
rect 8941 15651 8999 15657
rect 9324 15660 9772 15688
rect 4890 15620 4896 15632
rect 4540 15592 4896 15620
rect 4062 15552 4068 15564
rect 2424 15524 4068 15552
rect 1394 15444 1400 15496
rect 1452 15484 1458 15496
rect 2424 15493 2452 15524
rect 4062 15512 4068 15524
rect 4120 15512 4126 15564
rect 4540 15561 4568 15592
rect 4890 15580 4896 15592
rect 4948 15580 4954 15632
rect 5442 15580 5448 15632
rect 5500 15620 5506 15632
rect 5718 15620 5724 15632
rect 5500 15592 5724 15620
rect 5500 15580 5506 15592
rect 5718 15580 5724 15592
rect 5776 15580 5782 15632
rect 6362 15580 6368 15632
rect 6420 15620 6426 15632
rect 6420 15592 8064 15620
rect 6420 15580 6426 15592
rect 4525 15555 4583 15561
rect 4525 15521 4537 15555
rect 4571 15521 4583 15555
rect 4525 15515 4583 15521
rect 4709 15555 4767 15561
rect 4709 15521 4721 15555
rect 4755 15552 4767 15555
rect 5258 15552 5264 15564
rect 4755 15524 5264 15552
rect 4755 15521 4767 15524
rect 4709 15515 4767 15521
rect 5258 15512 5264 15524
rect 5316 15512 5322 15564
rect 5350 15512 5356 15564
rect 5408 15552 5414 15564
rect 5408 15524 5453 15552
rect 5408 15512 5414 15524
rect 5626 15512 5632 15564
rect 5684 15552 5690 15564
rect 6549 15555 6607 15561
rect 6549 15552 6561 15555
rect 5684 15524 6561 15552
rect 5684 15512 5690 15524
rect 6549 15521 6561 15524
rect 6595 15521 6607 15555
rect 6730 15552 6736 15564
rect 6691 15524 6736 15552
rect 6549 15515 6607 15521
rect 6730 15512 6736 15524
rect 6788 15512 6794 15564
rect 7742 15552 7748 15564
rect 7703 15524 7748 15552
rect 7742 15512 7748 15524
rect 7800 15512 7806 15564
rect 7926 15552 7932 15564
rect 7887 15524 7932 15552
rect 7926 15512 7932 15524
rect 7984 15512 7990 15564
rect 8036 15552 8064 15592
rect 8294 15580 8300 15632
rect 8352 15620 8358 15632
rect 8389 15623 8447 15629
rect 8389 15620 8401 15623
rect 8352 15592 8401 15620
rect 8352 15580 8358 15592
rect 8389 15589 8401 15592
rect 8435 15589 8447 15623
rect 8389 15583 8447 15589
rect 9324 15552 9352 15660
rect 9508 15561 9536 15660
rect 9766 15648 9772 15660
rect 9824 15648 9830 15700
rect 9861 15691 9919 15697
rect 9861 15657 9873 15691
rect 9907 15688 9919 15691
rect 10410 15688 10416 15700
rect 9907 15660 10416 15688
rect 9907 15657 9919 15660
rect 9861 15651 9919 15657
rect 10410 15648 10416 15660
rect 10468 15648 10474 15700
rect 11330 15648 11336 15700
rect 11388 15688 11394 15700
rect 11790 15688 11796 15700
rect 11388 15660 11796 15688
rect 11388 15648 11394 15660
rect 11790 15648 11796 15660
rect 11848 15688 11854 15700
rect 11848 15660 13492 15688
rect 11848 15648 11854 15660
rect 10229 15623 10287 15629
rect 10229 15620 10241 15623
rect 9692 15592 10241 15620
rect 8036 15524 9352 15552
rect 9493 15555 9551 15561
rect 9493 15521 9505 15555
rect 9539 15521 9551 15555
rect 9493 15515 9551 15521
rect 1673 15487 1731 15493
rect 1673 15484 1685 15487
rect 1452 15456 1685 15484
rect 1452 15444 1458 15456
rect 1673 15453 1685 15456
rect 1719 15453 1731 15487
rect 1673 15447 1731 15453
rect 2041 15487 2099 15493
rect 2041 15453 2053 15487
rect 2087 15453 2099 15487
rect 2041 15447 2099 15453
rect 2409 15487 2467 15493
rect 2409 15453 2421 15487
rect 2455 15453 2467 15487
rect 2409 15447 2467 15453
rect 2685 15487 2743 15493
rect 2685 15453 2697 15487
rect 2731 15484 2743 15487
rect 4430 15484 4436 15496
rect 2731 15456 4436 15484
rect 2731 15453 2743 15456
rect 2685 15447 2743 15453
rect 2056 15416 2084 15447
rect 4430 15444 4436 15456
rect 4488 15444 4494 15496
rect 4614 15444 4620 15496
rect 4672 15484 4678 15496
rect 9306 15484 9312 15496
rect 4672 15456 5672 15484
rect 9267 15456 9312 15484
rect 4672 15444 4678 15456
rect 4246 15416 4252 15428
rect 2056 15388 4252 15416
rect 4246 15376 4252 15388
rect 4304 15376 4310 15428
rect 4522 15376 4528 15428
rect 4580 15416 4586 15428
rect 5644 15425 5672 15456
rect 9306 15444 9312 15456
rect 9364 15444 9370 15496
rect 9398 15444 9404 15496
rect 9456 15484 9462 15496
rect 9692 15484 9720 15592
rect 10229 15589 10241 15592
rect 10275 15589 10287 15623
rect 10229 15583 10287 15589
rect 10594 15580 10600 15632
rect 10652 15620 10658 15632
rect 13464 15620 13492 15660
rect 13740 15660 16160 15688
rect 13740 15620 13768 15660
rect 10652 15592 11376 15620
rect 13464 15592 13768 15620
rect 16132 15620 16160 15660
rect 16206 15648 16212 15700
rect 16264 15688 16270 15700
rect 16301 15691 16359 15697
rect 16301 15688 16313 15691
rect 16264 15660 16313 15688
rect 16264 15648 16270 15660
rect 16301 15657 16313 15660
rect 16347 15657 16359 15691
rect 18230 15688 18236 15700
rect 16301 15651 16359 15657
rect 16408 15660 18236 15688
rect 16408 15620 16436 15660
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 16132 15592 16436 15620
rect 10652 15580 10658 15592
rect 10873 15555 10931 15561
rect 10873 15521 10885 15555
rect 10919 15552 10931 15555
rect 11238 15552 11244 15564
rect 10919 15524 11244 15552
rect 10919 15521 10931 15524
rect 10873 15515 10931 15521
rect 11238 15512 11244 15524
rect 11296 15512 11302 15564
rect 9456 15456 9720 15484
rect 10597 15487 10655 15493
rect 9456 15444 9462 15456
rect 10597 15453 10609 15487
rect 10643 15484 10655 15487
rect 11146 15484 11152 15496
rect 10643 15456 11152 15484
rect 10643 15453 10655 15456
rect 10597 15447 10655 15453
rect 11146 15444 11152 15456
rect 11204 15444 11210 15496
rect 11348 15484 11376 15592
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15552 13415 15555
rect 13630 15552 13636 15564
rect 13403 15524 13636 15552
rect 13403 15521 13415 15524
rect 13357 15515 13415 15521
rect 13630 15512 13636 15524
rect 13688 15512 13694 15564
rect 11348 15456 14596 15484
rect 14568 15428 14596 15456
rect 15378 15444 15384 15496
rect 15436 15484 15442 15496
rect 15473 15487 15531 15493
rect 15473 15484 15485 15487
rect 15436 15456 15485 15484
rect 15436 15444 15442 15456
rect 15473 15453 15485 15456
rect 15519 15484 15531 15487
rect 15565 15487 15623 15493
rect 15565 15484 15577 15487
rect 15519 15456 15577 15484
rect 15519 15453 15531 15456
rect 15473 15447 15531 15453
rect 15565 15453 15577 15456
rect 15611 15453 15623 15487
rect 15565 15447 15623 15453
rect 17586 15444 17592 15496
rect 17644 15484 17650 15496
rect 17681 15487 17739 15493
rect 17681 15484 17693 15487
rect 17644 15456 17693 15484
rect 17644 15444 17650 15456
rect 17681 15453 17693 15456
rect 17727 15484 17739 15487
rect 17773 15487 17831 15493
rect 17773 15484 17785 15487
rect 17727 15456 17785 15484
rect 17727 15453 17739 15456
rect 17681 15447 17739 15453
rect 17773 15453 17785 15456
rect 17819 15453 17831 15487
rect 17773 15447 17831 15453
rect 21450 15444 21456 15496
rect 21508 15484 21514 15496
rect 21545 15487 21603 15493
rect 21545 15484 21557 15487
rect 21508 15456 21557 15484
rect 21508 15444 21514 15456
rect 21545 15453 21557 15456
rect 21591 15453 21603 15487
rect 21545 15447 21603 15453
rect 4801 15419 4859 15425
rect 4801 15416 4813 15419
rect 4580 15388 4813 15416
rect 4580 15376 4586 15388
rect 4801 15385 4813 15388
rect 4847 15385 4859 15419
rect 4801 15379 4859 15385
rect 5629 15419 5687 15425
rect 5629 15385 5641 15419
rect 5675 15385 5687 15419
rect 6546 15416 6552 15428
rect 5629 15379 5687 15385
rect 5736 15388 6552 15416
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 2866 15308 2872 15360
rect 2924 15348 2930 15360
rect 3789 15351 3847 15357
rect 3789 15348 3801 15351
rect 2924 15320 3801 15348
rect 2924 15308 2930 15320
rect 3789 15317 3801 15320
rect 3835 15317 3847 15351
rect 3789 15311 3847 15317
rect 3878 15308 3884 15360
rect 3936 15348 3942 15360
rect 4540 15348 4568 15376
rect 3936 15320 4568 15348
rect 5537 15351 5595 15357
rect 3936 15308 3942 15320
rect 5537 15317 5549 15351
rect 5583 15348 5595 15351
rect 5736 15348 5764 15388
rect 6546 15376 6552 15388
rect 6604 15376 6610 15428
rect 7742 15376 7748 15428
rect 7800 15416 7806 15428
rect 10962 15416 10968 15428
rect 7800 15388 10968 15416
rect 7800 15376 7806 15388
rect 10962 15376 10968 15388
rect 11020 15376 11026 15428
rect 13112 15419 13170 15425
rect 13112 15385 13124 15419
rect 13158 15416 13170 15419
rect 13722 15416 13728 15428
rect 13158 15388 13728 15416
rect 13158 15385 13170 15388
rect 13112 15379 13170 15385
rect 13722 15376 13728 15388
rect 13780 15376 13786 15428
rect 14550 15376 14556 15428
rect 14608 15376 14614 15428
rect 14918 15376 14924 15428
rect 14976 15416 14982 15428
rect 15206 15419 15264 15425
rect 15206 15416 15218 15419
rect 14976 15388 15218 15416
rect 14976 15376 14982 15388
rect 15206 15385 15218 15388
rect 15252 15416 15264 15419
rect 15749 15419 15807 15425
rect 15749 15416 15761 15419
rect 15252 15388 15761 15416
rect 15252 15385 15264 15388
rect 15206 15379 15264 15385
rect 15749 15385 15761 15388
rect 15795 15385 15807 15419
rect 15749 15379 15807 15385
rect 16390 15376 16396 15428
rect 16448 15416 16454 15428
rect 17414 15419 17472 15425
rect 17414 15416 17426 15419
rect 16448 15388 17426 15416
rect 16448 15376 16454 15388
rect 17414 15385 17426 15388
rect 17460 15385 17472 15419
rect 21266 15416 21272 15428
rect 21324 15425 21330 15428
rect 21236 15388 21272 15416
rect 17414 15379 17472 15385
rect 21266 15376 21272 15388
rect 21324 15379 21336 15425
rect 21324 15376 21330 15379
rect 5583 15320 5764 15348
rect 5583 15317 5595 15320
rect 5537 15311 5595 15317
rect 5994 15308 6000 15360
rect 6052 15348 6058 15360
rect 6457 15351 6515 15357
rect 6457 15348 6469 15351
rect 6052 15320 6469 15348
rect 6052 15308 6058 15320
rect 6457 15317 6469 15320
rect 6503 15317 6515 15351
rect 6457 15311 6515 15317
rect 7006 15308 7012 15360
rect 7064 15348 7070 15360
rect 8021 15351 8079 15357
rect 8021 15348 8033 15351
rect 7064 15320 8033 15348
rect 7064 15308 7070 15320
rect 8021 15317 8033 15320
rect 8067 15317 8079 15351
rect 8021 15311 8079 15317
rect 8662 15308 8668 15360
rect 8720 15348 8726 15360
rect 9401 15351 9459 15357
rect 9401 15348 9413 15351
rect 8720 15320 9413 15348
rect 8720 15308 8726 15320
rect 9401 15317 9413 15320
rect 9447 15317 9459 15351
rect 9401 15311 9459 15317
rect 9674 15308 9680 15360
rect 9732 15348 9738 15360
rect 9953 15351 10011 15357
rect 9953 15348 9965 15351
rect 9732 15320 9965 15348
rect 9732 15308 9738 15320
rect 9953 15317 9965 15320
rect 9999 15317 10011 15351
rect 9953 15311 10011 15317
rect 10686 15308 10692 15360
rect 10744 15348 10750 15360
rect 11977 15351 12035 15357
rect 10744 15320 10789 15348
rect 10744 15308 10750 15320
rect 11977 15317 11989 15351
rect 12023 15348 12035 15351
rect 12802 15348 12808 15360
rect 12023 15320 12808 15348
rect 12023 15317 12035 15320
rect 11977 15311 12035 15317
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 13541 15351 13599 15357
rect 13541 15317 13553 15351
rect 13587 15348 13599 15351
rect 13630 15348 13636 15360
rect 13587 15320 13636 15348
rect 13587 15317 13599 15320
rect 13541 15311 13599 15317
rect 13630 15308 13636 15320
rect 13688 15308 13694 15360
rect 13814 15308 13820 15360
rect 13872 15348 13878 15360
rect 14093 15351 14151 15357
rect 14093 15348 14105 15351
rect 13872 15320 14105 15348
rect 13872 15308 13878 15320
rect 14093 15317 14105 15320
rect 14139 15317 14151 15351
rect 19794 15348 19800 15360
rect 19755 15320 19800 15348
rect 14093 15311 14151 15317
rect 19794 15308 19800 15320
rect 19852 15348 19858 15360
rect 19981 15351 20039 15357
rect 19981 15348 19993 15351
rect 19852 15320 19993 15348
rect 19852 15308 19858 15320
rect 19981 15317 19993 15320
rect 20027 15317 20039 15351
rect 19981 15311 20039 15317
rect 20165 15351 20223 15357
rect 20165 15317 20177 15351
rect 20211 15348 20223 15351
rect 20622 15348 20628 15360
rect 20211 15320 20628 15348
rect 20211 15317 20223 15320
rect 20165 15311 20223 15317
rect 20622 15308 20628 15320
rect 20680 15308 20686 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 2038 15104 2044 15156
rect 2096 15144 2102 15156
rect 2133 15147 2191 15153
rect 2133 15144 2145 15147
rect 2096 15116 2145 15144
rect 2096 15104 2102 15116
rect 2133 15113 2145 15116
rect 2179 15113 2191 15147
rect 2133 15107 2191 15113
rect 2222 15104 2228 15156
rect 2280 15144 2286 15156
rect 2593 15147 2651 15153
rect 2593 15144 2605 15147
rect 2280 15116 2605 15144
rect 2280 15104 2286 15116
rect 2593 15113 2605 15116
rect 2639 15113 2651 15147
rect 2593 15107 2651 15113
rect 3329 15147 3387 15153
rect 3329 15113 3341 15147
rect 3375 15144 3387 15147
rect 3878 15144 3884 15156
rect 3375 15116 3884 15144
rect 3375 15113 3387 15116
rect 3329 15107 3387 15113
rect 3878 15104 3884 15116
rect 3936 15104 3942 15156
rect 4985 15147 5043 15153
rect 4985 15144 4997 15147
rect 4448 15116 4997 15144
rect 4338 15076 4344 15088
rect 2792 15048 4344 15076
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 1762 15008 1768 15020
rect 1719 14980 1768 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 1762 14968 1768 14980
rect 1820 14968 1826 15020
rect 2038 15008 2044 15020
rect 1999 14980 2044 15008
rect 2038 14968 2044 14980
rect 2096 14968 2102 15020
rect 2792 15017 2820 15048
rect 4338 15036 4344 15048
rect 4396 15036 4402 15088
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 14977 2375 15011
rect 2317 14971 2375 14977
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 14977 2835 15011
rect 2777 14971 2835 14977
rect 4157 15011 4215 15017
rect 4157 14977 4169 15011
rect 4203 15008 4215 15011
rect 4448 15008 4476 15116
rect 4985 15113 4997 15116
rect 5031 15144 5043 15147
rect 5810 15144 5816 15156
rect 5031 15116 5816 15144
rect 5031 15113 5043 15116
rect 4985 15107 5043 15113
rect 5810 15104 5816 15116
rect 5868 15104 5874 15156
rect 7466 15144 7472 15156
rect 7427 15116 7472 15144
rect 7466 15104 7472 15116
rect 7524 15104 7530 15156
rect 7558 15104 7564 15156
rect 7616 15144 7622 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7616 15116 7849 15144
rect 7616 15104 7622 15116
rect 7837 15113 7849 15116
rect 7883 15113 7895 15147
rect 7837 15107 7895 15113
rect 7926 15104 7932 15156
rect 7984 15144 7990 15156
rect 7984 15116 8432 15144
rect 7984 15104 7990 15116
rect 4798 15076 4804 15088
rect 4203 14980 4476 15008
rect 4540 15048 4804 15076
rect 4203 14977 4215 14980
rect 4157 14971 4215 14977
rect 2332 14940 2360 14971
rect 4540 14952 4568 15048
rect 4798 15036 4804 15048
rect 4856 15036 4862 15088
rect 6822 15036 6828 15088
rect 6880 15076 6886 15088
rect 8297 15079 8355 15085
rect 8297 15076 8309 15079
rect 6880 15048 8309 15076
rect 6880 15036 6886 15048
rect 8297 15045 8309 15048
rect 8343 15045 8355 15079
rect 8297 15039 8355 15045
rect 4724 14980 5580 15008
rect 2958 14940 2964 14952
rect 2332 14912 2964 14940
rect 2958 14900 2964 14912
rect 3016 14900 3022 14952
rect 3053 14943 3111 14949
rect 3053 14909 3065 14943
rect 3099 14909 3111 14943
rect 3053 14903 3111 14909
rect 3237 14943 3295 14949
rect 3237 14909 3249 14943
rect 3283 14909 3295 14943
rect 3237 14903 3295 14909
rect 1854 14872 1860 14884
rect 1815 14844 1860 14872
rect 1854 14832 1860 14844
rect 1912 14832 1918 14884
rect 2866 14832 2872 14884
rect 2924 14872 2930 14884
rect 3068 14872 3096 14903
rect 2924 14844 3096 14872
rect 3252 14872 3280 14903
rect 3418 14900 3424 14952
rect 3476 14940 3482 14952
rect 3881 14943 3939 14949
rect 3881 14940 3893 14943
rect 3476 14912 3893 14940
rect 3476 14900 3482 14912
rect 3881 14909 3893 14912
rect 3927 14909 3939 14943
rect 3881 14903 3939 14909
rect 4065 14943 4123 14949
rect 4065 14909 4077 14943
rect 4111 14940 4123 14943
rect 4522 14940 4528 14952
rect 4111 14912 4528 14940
rect 4111 14909 4123 14912
rect 4065 14903 4123 14909
rect 4522 14900 4528 14912
rect 4580 14900 4586 14952
rect 4724 14949 4752 14980
rect 4709 14943 4767 14949
rect 4709 14909 4721 14943
rect 4755 14909 4767 14943
rect 4890 14940 4896 14952
rect 4851 14912 4896 14940
rect 4709 14903 4767 14909
rect 4890 14900 4896 14912
rect 4948 14900 4954 14952
rect 5350 14900 5356 14952
rect 5408 14940 5414 14952
rect 5445 14943 5503 14949
rect 5445 14940 5457 14943
rect 5408 14912 5457 14940
rect 5408 14900 5414 14912
rect 5445 14909 5457 14912
rect 5491 14909 5503 14943
rect 5552 14940 5580 14980
rect 5718 14968 5724 15020
rect 5776 15008 5782 15020
rect 7101 15011 7159 15017
rect 7101 15008 7113 15011
rect 5776 14980 7113 15008
rect 5776 14968 5782 14980
rect 7101 14977 7113 14980
rect 7147 14977 7159 15011
rect 7101 14971 7159 14977
rect 7745 15011 7803 15017
rect 7745 14977 7757 15011
rect 7791 15008 7803 15011
rect 8202 15008 8208 15020
rect 7791 14980 8208 15008
rect 7791 14977 7803 14980
rect 7745 14971 7803 14977
rect 8202 14968 8208 14980
rect 8260 14968 8266 15020
rect 8404 15008 8432 15116
rect 8570 15104 8576 15156
rect 8628 15144 8634 15156
rect 8941 15147 8999 15153
rect 8941 15144 8953 15147
rect 8628 15116 8953 15144
rect 8628 15104 8634 15116
rect 8941 15113 8953 15116
rect 8987 15113 8999 15147
rect 8941 15107 8999 15113
rect 9030 15104 9036 15156
rect 9088 15144 9094 15156
rect 9490 15144 9496 15156
rect 9088 15116 9133 15144
rect 9451 15116 9496 15144
rect 9088 15104 9094 15116
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 10597 15147 10655 15153
rect 10597 15113 10609 15147
rect 10643 15144 10655 15147
rect 10686 15144 10692 15156
rect 10643 15116 10692 15144
rect 10643 15113 10655 15116
rect 10597 15107 10655 15113
rect 10686 15104 10692 15116
rect 10744 15104 10750 15156
rect 11057 15147 11115 15153
rect 11057 15113 11069 15147
rect 11103 15144 11115 15147
rect 13446 15144 13452 15156
rect 11103 15116 13452 15144
rect 11103 15113 11115 15116
rect 11057 15107 11115 15113
rect 13446 15104 13452 15116
rect 13504 15104 13510 15156
rect 13078 15076 13084 15088
rect 9140 15048 13084 15076
rect 9140 15008 9168 15048
rect 13078 15036 13084 15048
rect 13136 15036 13142 15088
rect 16942 15085 16948 15088
rect 16936 15076 16948 15085
rect 16903 15048 16948 15076
rect 16936 15039 16948 15048
rect 16942 15036 16948 15039
rect 17000 15036 17006 15088
rect 19794 15076 19800 15088
rect 18156 15048 19800 15076
rect 8404 14980 9168 15008
rect 9766 14968 9772 15020
rect 9824 15008 9830 15020
rect 9861 15011 9919 15017
rect 9861 15008 9873 15011
rect 9824 14980 9873 15008
rect 9824 14968 9830 14980
rect 9861 14977 9873 14980
rect 9907 14977 9919 15011
rect 9861 14971 9919 14977
rect 10410 14968 10416 15020
rect 10468 15008 10474 15020
rect 10965 15011 11023 15017
rect 10965 15008 10977 15011
rect 10468 14980 10977 15008
rect 10468 14968 10474 14980
rect 10965 14977 10977 14980
rect 11011 14977 11023 15011
rect 11698 15008 11704 15020
rect 10965 14971 11023 14977
rect 11072 14980 11704 15008
rect 6730 14940 6736 14952
rect 5552 14912 6736 14940
rect 5445 14903 5503 14909
rect 6730 14900 6736 14912
rect 6788 14900 6794 14952
rect 6914 14940 6920 14952
rect 6875 14912 6920 14940
rect 6914 14900 6920 14912
rect 6972 14900 6978 14952
rect 7009 14943 7067 14949
rect 7009 14909 7021 14943
rect 7055 14940 7067 14943
rect 7282 14940 7288 14952
rect 7055 14912 7288 14940
rect 7055 14909 7067 14912
rect 7009 14903 7067 14909
rect 7282 14900 7288 14912
rect 7340 14900 7346 14952
rect 8110 14900 8116 14952
rect 8168 14940 8174 14952
rect 8389 14943 8447 14949
rect 8389 14940 8401 14943
rect 8168 14912 8401 14940
rect 8168 14900 8174 14912
rect 8389 14909 8401 14912
rect 8435 14909 8447 14943
rect 8389 14903 8447 14909
rect 8849 14943 8907 14949
rect 8849 14909 8861 14943
rect 8895 14909 8907 14943
rect 8849 14903 8907 14909
rect 4614 14872 4620 14884
rect 3252 14844 4620 14872
rect 2924 14832 2930 14844
rect 4614 14832 4620 14844
rect 4672 14832 4678 14884
rect 6822 14872 6828 14884
rect 5276 14844 6828 14872
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 3697 14807 3755 14813
rect 3697 14773 3709 14807
rect 3743 14804 3755 14807
rect 3970 14804 3976 14816
rect 3743 14776 3976 14804
rect 3743 14773 3755 14776
rect 3697 14767 3755 14773
rect 3970 14764 3976 14776
rect 4028 14764 4034 14816
rect 4525 14807 4583 14813
rect 4525 14773 4537 14807
rect 4571 14804 4583 14807
rect 5276 14804 5304 14844
rect 6822 14832 6828 14844
rect 6880 14832 6886 14884
rect 7926 14872 7932 14884
rect 6932 14844 7932 14872
rect 4571 14776 5304 14804
rect 5353 14807 5411 14813
rect 4571 14773 4583 14776
rect 4525 14767 4583 14773
rect 5353 14773 5365 14807
rect 5399 14804 5411 14807
rect 5810 14804 5816 14816
rect 5399 14776 5816 14804
rect 5399 14773 5411 14776
rect 5353 14767 5411 14773
rect 5810 14764 5816 14776
rect 5868 14764 5874 14816
rect 5994 14804 6000 14816
rect 5955 14776 6000 14804
rect 5994 14764 6000 14776
rect 6052 14764 6058 14816
rect 6730 14764 6736 14816
rect 6788 14804 6794 14816
rect 6932 14804 6960 14844
rect 7926 14832 7932 14844
rect 7984 14832 7990 14884
rect 8018 14832 8024 14884
rect 8076 14872 8082 14884
rect 8864 14872 8892 14903
rect 9122 14900 9128 14952
rect 9180 14940 9186 14952
rect 9953 14943 10011 14949
rect 9953 14940 9965 14943
rect 9180 14912 9965 14940
rect 9180 14900 9186 14912
rect 9953 14909 9965 14912
rect 9999 14909 10011 14943
rect 9953 14903 10011 14909
rect 10137 14943 10195 14949
rect 10137 14909 10149 14943
rect 10183 14940 10195 14943
rect 11072 14940 11100 14980
rect 11698 14968 11704 14980
rect 11756 14968 11762 15020
rect 12710 15008 12716 15020
rect 12406 14980 12716 15008
rect 11238 14940 11244 14952
rect 10183 14912 11100 14940
rect 11199 14912 11244 14940
rect 10183 14909 10195 14912
rect 10137 14903 10195 14909
rect 11238 14900 11244 14912
rect 11296 14900 11302 14952
rect 9674 14872 9680 14884
rect 8076 14844 9680 14872
rect 8076 14832 8082 14844
rect 9674 14832 9680 14844
rect 9732 14832 9738 14884
rect 12069 14875 12127 14881
rect 12069 14841 12081 14875
rect 12115 14872 12127 14875
rect 12406 14872 12434 14980
rect 12710 14968 12716 14980
rect 12768 14968 12774 15020
rect 12894 14968 12900 15020
rect 12952 15008 12958 15020
rect 13182 15011 13240 15017
rect 13182 15008 13194 15011
rect 12952 14980 13194 15008
rect 12952 14968 12958 14980
rect 13182 14977 13194 14980
rect 13228 14977 13240 15011
rect 13182 14971 13240 14977
rect 15010 14968 15016 15020
rect 15068 15017 15074 15020
rect 15068 15008 15080 15017
rect 15068 14980 15113 15008
rect 15068 14971 15080 14980
rect 15068 14968 15074 14971
rect 15194 14968 15200 15020
rect 15252 15008 15258 15020
rect 15289 15011 15347 15017
rect 15289 15008 15301 15011
rect 15252 14980 15301 15008
rect 15252 14968 15258 14980
rect 15289 14977 15301 14980
rect 15335 15008 15347 15011
rect 15381 15011 15439 15017
rect 15381 15008 15393 15011
rect 15335 14980 15393 15008
rect 15335 14977 15347 14980
rect 15289 14971 15347 14977
rect 15381 14977 15393 14980
rect 15427 15008 15439 15011
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 15427 14980 16681 15008
rect 15427 14977 15439 14980
rect 15381 14971 15439 14977
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 17678 14968 17684 15020
rect 17736 15008 17742 15020
rect 18156 15017 18184 15048
rect 19720 15017 19748 15048
rect 19794 15036 19800 15048
rect 19852 15036 19858 15088
rect 18141 15011 18199 15017
rect 18141 15008 18153 15011
rect 17736 14980 18153 15008
rect 17736 14968 17742 14980
rect 18141 14977 18153 14980
rect 18187 14977 18199 15011
rect 18141 14971 18199 14977
rect 19449 15011 19507 15017
rect 19449 14977 19461 15011
rect 19495 15008 19507 15011
rect 19705 15011 19763 15017
rect 19495 14980 19656 15008
rect 19495 14977 19507 14980
rect 19449 14971 19507 14977
rect 13449 14943 13507 14949
rect 13449 14909 13461 14943
rect 13495 14909 13507 14943
rect 19628 14940 19656 14980
rect 19705 14977 19717 15011
rect 19751 14977 19763 15011
rect 19705 14971 19763 14977
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 21002 15011 21060 15017
rect 21002 15008 21014 15011
rect 20772 14980 21014 15008
rect 20772 14968 20778 14980
rect 21002 14977 21014 14980
rect 21048 14977 21060 15011
rect 21002 14971 21060 14977
rect 19794 14940 19800 14952
rect 19628 14912 19800 14940
rect 13449 14903 13507 14909
rect 12115 14844 12434 14872
rect 13464 14872 13492 14903
rect 19794 14900 19800 14912
rect 19852 14900 19858 14952
rect 21269 14943 21327 14949
rect 21269 14909 21281 14943
rect 21315 14909 21327 14943
rect 21269 14903 21327 14909
rect 13630 14872 13636 14884
rect 13464 14844 13636 14872
rect 12115 14841 12127 14844
rect 12069 14835 12127 14841
rect 13630 14832 13636 14844
rect 13688 14832 13694 14884
rect 14274 14872 14280 14884
rect 13832 14844 14280 14872
rect 6788 14776 6960 14804
rect 6788 14764 6794 14776
rect 7374 14764 7380 14816
rect 7432 14804 7438 14816
rect 8110 14804 8116 14816
rect 7432 14776 8116 14804
rect 7432 14764 7438 14776
rect 8110 14764 8116 14776
rect 8168 14764 8174 14816
rect 9398 14804 9404 14816
rect 9359 14776 9404 14804
rect 9398 14764 9404 14776
rect 9456 14764 9462 14816
rect 10410 14804 10416 14816
rect 10371 14776 10416 14804
rect 10410 14764 10416 14776
rect 10468 14764 10474 14816
rect 12710 14764 12716 14816
rect 12768 14804 12774 14816
rect 13832 14804 13860 14844
rect 14274 14832 14280 14844
rect 14332 14832 14338 14884
rect 17604 14844 18460 14872
rect 12768 14776 13860 14804
rect 13909 14807 13967 14813
rect 12768 14764 12774 14776
rect 13909 14773 13921 14807
rect 13955 14804 13967 14807
rect 14366 14804 14372 14816
rect 13955 14776 14372 14804
rect 13955 14773 13967 14776
rect 13909 14767 13967 14773
rect 14366 14764 14372 14776
rect 14424 14764 14430 14816
rect 15746 14764 15752 14816
rect 15804 14804 15810 14816
rect 16117 14807 16175 14813
rect 16117 14804 16129 14807
rect 15804 14776 16129 14804
rect 15804 14764 15810 14776
rect 16117 14773 16129 14776
rect 16163 14804 16175 14807
rect 17604 14804 17632 14844
rect 18046 14804 18052 14816
rect 16163 14776 17632 14804
rect 18007 14776 18052 14804
rect 16163 14773 16175 14776
rect 16117 14767 16175 14773
rect 18046 14764 18052 14776
rect 18104 14764 18110 14816
rect 18322 14804 18328 14816
rect 18283 14776 18328 14804
rect 18322 14764 18328 14776
rect 18380 14764 18386 14816
rect 18432 14804 18460 14844
rect 19889 14807 19947 14813
rect 19889 14804 19901 14807
rect 18432 14776 19901 14804
rect 19889 14773 19901 14776
rect 19935 14773 19947 14807
rect 19889 14767 19947 14773
rect 21082 14764 21088 14816
rect 21140 14804 21146 14816
rect 21284 14804 21312 14903
rect 21361 14807 21419 14813
rect 21361 14804 21373 14807
rect 21140 14776 21373 14804
rect 21140 14764 21146 14776
rect 21361 14773 21373 14776
rect 21407 14773 21419 14807
rect 21361 14767 21419 14773
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 4617 14603 4675 14609
rect 4617 14569 4629 14603
rect 4663 14600 4675 14603
rect 4890 14600 4896 14612
rect 4663 14572 4896 14600
rect 4663 14569 4675 14572
rect 4617 14563 4675 14569
rect 4890 14560 4896 14572
rect 4948 14560 4954 14612
rect 6641 14603 6699 14609
rect 6641 14569 6653 14603
rect 6687 14600 6699 14603
rect 9122 14600 9128 14612
rect 6687 14572 9128 14600
rect 6687 14569 6699 14572
rect 6641 14563 6699 14569
rect 9122 14560 9128 14572
rect 9180 14560 9186 14612
rect 9858 14600 9864 14612
rect 9819 14572 9864 14600
rect 9858 14560 9864 14572
rect 9916 14560 9922 14612
rect 11238 14560 11244 14612
rect 11296 14600 11302 14612
rect 11296 14572 14596 14600
rect 11296 14560 11302 14572
rect 4706 14492 4712 14544
rect 4764 14532 4770 14544
rect 4764 14504 5212 14532
rect 4764 14492 4770 14504
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 4614 14464 4620 14476
rect 4111 14436 4620 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 4614 14424 4620 14436
rect 4672 14424 4678 14476
rect 5074 14464 5080 14476
rect 5035 14436 5080 14464
rect 5074 14424 5080 14436
rect 5132 14424 5138 14476
rect 5184 14464 5212 14504
rect 5810 14492 5816 14544
rect 5868 14532 5874 14544
rect 8294 14532 8300 14544
rect 5868 14504 6224 14532
rect 5868 14492 5874 14504
rect 6196 14473 6224 14504
rect 8036 14504 8300 14532
rect 6089 14467 6147 14473
rect 5184 14436 5304 14464
rect 5276 14408 5304 14436
rect 6089 14433 6101 14467
rect 6135 14433 6147 14467
rect 6089 14427 6147 14433
rect 6181 14467 6239 14473
rect 6181 14433 6193 14467
rect 6227 14433 6239 14467
rect 6181 14427 6239 14433
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 1854 14396 1860 14408
rect 1719 14368 1860 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 1854 14356 1860 14368
rect 1912 14356 1918 14408
rect 4154 14356 4160 14408
rect 4212 14396 4218 14408
rect 4249 14399 4307 14405
rect 4249 14396 4261 14399
rect 4212 14368 4261 14396
rect 4212 14356 4218 14368
rect 4249 14365 4261 14368
rect 4295 14396 4307 14399
rect 5169 14399 5227 14405
rect 5169 14396 5181 14399
rect 4295 14368 5181 14396
rect 4295 14365 4307 14368
rect 4249 14359 4307 14365
rect 5169 14365 5181 14368
rect 5215 14365 5227 14399
rect 5169 14359 5227 14365
rect 5258 14356 5264 14408
rect 5316 14396 5322 14408
rect 6104 14396 6132 14427
rect 7098 14424 7104 14476
rect 7156 14464 7162 14476
rect 7466 14464 7472 14476
rect 7156 14436 7472 14464
rect 7156 14424 7162 14436
rect 7466 14424 7472 14436
rect 7524 14464 7530 14476
rect 7926 14464 7932 14476
rect 7524 14436 7932 14464
rect 7524 14424 7530 14436
rect 7926 14424 7932 14436
rect 7984 14424 7990 14476
rect 8036 14473 8064 14504
rect 8294 14492 8300 14504
rect 8352 14532 8358 14544
rect 8389 14535 8447 14541
rect 8389 14532 8401 14535
rect 8352 14504 8401 14532
rect 8352 14492 8358 14504
rect 8389 14501 8401 14504
rect 8435 14501 8447 14535
rect 8389 14495 8447 14501
rect 8754 14492 8760 14544
rect 8812 14532 8818 14544
rect 12158 14532 12164 14544
rect 8812 14504 12164 14532
rect 8812 14492 8818 14504
rect 12158 14492 12164 14504
rect 12216 14492 12222 14544
rect 8021 14467 8079 14473
rect 8021 14433 8033 14467
rect 8067 14433 8079 14467
rect 8021 14427 8079 14433
rect 8110 14424 8116 14476
rect 8168 14464 8174 14476
rect 9306 14464 9312 14476
rect 8168 14436 8213 14464
rect 9267 14436 9312 14464
rect 8168 14424 8174 14436
rect 9306 14424 9312 14436
rect 9364 14424 9370 14476
rect 9398 14424 9404 14476
rect 9456 14464 9462 14476
rect 10413 14467 10471 14473
rect 10413 14464 10425 14467
rect 9456 14436 10425 14464
rect 9456 14424 9462 14436
rect 10413 14433 10425 14436
rect 10459 14433 10471 14467
rect 10413 14427 10471 14433
rect 10502 14424 10508 14476
rect 10560 14464 10566 14476
rect 11146 14464 11152 14476
rect 10560 14436 11152 14464
rect 10560 14424 10566 14436
rect 11146 14424 11152 14436
rect 11204 14424 11210 14476
rect 13541 14467 13599 14473
rect 13541 14433 13553 14467
rect 13587 14464 13599 14467
rect 13630 14464 13636 14476
rect 13587 14436 13636 14464
rect 13587 14433 13599 14436
rect 13541 14427 13599 14433
rect 13630 14424 13636 14436
rect 13688 14464 13694 14476
rect 13725 14467 13783 14473
rect 13725 14464 13737 14467
rect 13688 14436 13737 14464
rect 13688 14424 13694 14436
rect 13725 14433 13737 14436
rect 13771 14464 13783 14467
rect 13906 14464 13912 14476
rect 13771 14436 13912 14464
rect 13771 14433 13783 14436
rect 13725 14427 13783 14433
rect 13906 14424 13912 14436
rect 13964 14424 13970 14476
rect 6270 14396 6276 14408
rect 5316 14368 5409 14396
rect 6104 14368 6276 14396
rect 5316 14356 5322 14368
rect 6270 14356 6276 14368
rect 6328 14356 6334 14408
rect 8846 14356 8852 14408
rect 8904 14396 8910 14408
rect 9493 14399 9551 14405
rect 9493 14396 9505 14399
rect 8904 14368 9505 14396
rect 8904 14356 8910 14368
rect 9493 14365 9505 14368
rect 9539 14365 9551 14399
rect 10318 14396 10324 14408
rect 10279 14368 10324 14396
rect 9493 14359 9551 14365
rect 10318 14356 10324 14368
rect 10376 14356 10382 14408
rect 13814 14396 13820 14408
rect 13289 14368 13820 14396
rect 3418 14288 3424 14340
rect 3476 14328 3482 14340
rect 4801 14331 4859 14337
rect 4801 14328 4813 14331
rect 3476 14300 4813 14328
rect 3476 14288 3482 14300
rect 4801 14297 4813 14300
rect 4847 14328 4859 14331
rect 7926 14328 7932 14340
rect 4847 14300 7696 14328
rect 7887 14300 7932 14328
rect 4847 14297 4859 14300
rect 4801 14291 4859 14297
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 4157 14263 4215 14269
rect 4157 14229 4169 14263
rect 4203 14260 4215 14263
rect 4522 14260 4528 14272
rect 4203 14232 4528 14260
rect 4203 14229 4215 14232
rect 4157 14223 4215 14229
rect 4522 14220 4528 14232
rect 4580 14220 4586 14272
rect 5626 14260 5632 14272
rect 5587 14232 5632 14260
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 6273 14263 6331 14269
rect 6273 14229 6285 14263
rect 6319 14260 6331 14263
rect 6546 14260 6552 14272
rect 6319 14232 6552 14260
rect 6319 14229 6331 14232
rect 6273 14223 6331 14229
rect 6546 14220 6552 14232
rect 6604 14220 6610 14272
rect 7558 14260 7564 14272
rect 7519 14232 7564 14260
rect 7558 14220 7564 14232
rect 7616 14220 7622 14272
rect 7668 14260 7696 14300
rect 7926 14288 7932 14300
rect 7984 14288 7990 14340
rect 9401 14331 9459 14337
rect 9401 14297 9413 14331
rect 9447 14328 9459 14331
rect 9447 14300 9996 14328
rect 9447 14297 9459 14300
rect 9401 14291 9459 14297
rect 9858 14260 9864 14272
rect 7668 14232 9864 14260
rect 9858 14220 9864 14232
rect 9916 14220 9922 14272
rect 9968 14269 9996 14300
rect 10962 14288 10968 14340
rect 11020 14328 11026 14340
rect 13289 14337 13317 14368
rect 13814 14356 13820 14368
rect 13872 14356 13878 14408
rect 13274 14331 13332 14337
rect 13274 14328 13286 14331
rect 11020 14300 13286 14328
rect 11020 14288 11026 14300
rect 13274 14297 13286 14300
rect 13320 14297 13332 14331
rect 13274 14291 13332 14297
rect 9953 14263 10011 14269
rect 9953 14229 9965 14263
rect 9999 14229 10011 14263
rect 12158 14260 12164 14272
rect 12119 14232 12164 14260
rect 9953 14223 10011 14229
rect 12158 14220 12164 14232
rect 12216 14220 12222 14272
rect 13538 14220 13544 14272
rect 13596 14260 13602 14272
rect 14458 14260 14464 14272
rect 13596 14232 14464 14260
rect 13596 14220 13602 14232
rect 14458 14220 14464 14232
rect 14516 14220 14522 14272
rect 14568 14260 14596 14572
rect 15194 14560 15200 14612
rect 15252 14600 15258 14612
rect 15933 14603 15991 14609
rect 15933 14600 15945 14603
rect 15252 14572 15945 14600
rect 15252 14560 15258 14572
rect 15856 14473 15884 14572
rect 15933 14569 15945 14572
rect 15979 14569 15991 14603
rect 16206 14600 16212 14612
rect 16119 14572 16212 14600
rect 15933 14563 15991 14569
rect 16206 14560 16212 14572
rect 16264 14600 16270 14612
rect 18138 14600 18144 14612
rect 16264 14572 18144 14600
rect 16264 14560 16270 14572
rect 18138 14560 18144 14572
rect 18196 14560 18202 14612
rect 15841 14467 15899 14473
rect 15841 14433 15853 14467
rect 15887 14433 15899 14467
rect 15841 14427 15899 14433
rect 14826 14356 14832 14408
rect 14884 14396 14890 14408
rect 15574 14399 15632 14405
rect 15574 14396 15586 14399
rect 14884 14368 15586 14396
rect 14884 14356 14890 14368
rect 15574 14365 15586 14368
rect 15620 14396 15632 14399
rect 15746 14396 15752 14408
rect 15620 14368 15752 14396
rect 15620 14365 15632 14368
rect 15574 14359 15632 14365
rect 15746 14356 15752 14368
rect 15804 14356 15810 14408
rect 17586 14396 17592 14408
rect 17547 14368 17592 14396
rect 17586 14356 17592 14368
rect 17644 14396 17650 14408
rect 17681 14399 17739 14405
rect 17681 14396 17693 14399
rect 17644 14368 17693 14396
rect 17644 14356 17650 14368
rect 17681 14365 17693 14368
rect 17727 14396 17739 14399
rect 18141 14399 18199 14405
rect 18141 14396 18153 14399
rect 17727 14368 18153 14396
rect 17727 14365 17739 14368
rect 17681 14359 17739 14365
rect 18141 14365 18153 14368
rect 18187 14365 18199 14399
rect 21082 14396 21088 14408
rect 21043 14368 21088 14396
rect 18141 14359 18199 14365
rect 21082 14356 21088 14368
rect 21140 14396 21146 14408
rect 21177 14399 21235 14405
rect 21177 14396 21189 14399
rect 21140 14368 21189 14396
rect 21140 14356 21146 14368
rect 21177 14365 21189 14368
rect 21223 14365 21235 14399
rect 21177 14359 21235 14365
rect 17344 14331 17402 14337
rect 17344 14297 17356 14331
rect 17390 14328 17402 14331
rect 17494 14328 17500 14340
rect 17390 14300 17500 14328
rect 17390 14297 17402 14300
rect 17344 14291 17402 14297
rect 17494 14288 17500 14300
rect 17552 14288 17558 14340
rect 20346 14328 20352 14340
rect 19628 14300 20352 14328
rect 19628 14260 19656 14300
rect 20346 14288 20352 14300
rect 20404 14288 20410 14340
rect 20898 14337 20904 14340
rect 20840 14331 20904 14337
rect 20840 14297 20852 14331
rect 20886 14297 20904 14331
rect 20840 14291 20904 14297
rect 20898 14288 20904 14291
rect 20956 14288 20962 14340
rect 14568 14232 19656 14260
rect 19705 14263 19763 14269
rect 19705 14229 19717 14263
rect 19751 14260 19763 14263
rect 19794 14260 19800 14272
rect 19751 14232 19800 14260
rect 19751 14229 19763 14232
rect 19705 14223 19763 14229
rect 19794 14220 19800 14232
rect 19852 14220 19858 14272
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 5350 14056 5356 14068
rect 5311 14028 5356 14056
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 5718 14056 5724 14068
rect 5679 14028 5724 14056
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 6365 14059 6423 14065
rect 6365 14025 6377 14059
rect 6411 14056 6423 14059
rect 6546 14056 6552 14068
rect 6411 14028 6552 14056
rect 6411 14025 6423 14028
rect 6365 14019 6423 14025
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 6730 14016 6736 14068
rect 6788 14056 6794 14068
rect 7282 14056 7288 14068
rect 6788 14028 6960 14056
rect 7243 14028 7288 14056
rect 6788 14016 6794 14028
rect 5258 13948 5264 14000
rect 5316 13988 5322 14000
rect 6825 13991 6883 13997
rect 6825 13988 6837 13991
rect 5316 13960 6837 13988
rect 5316 13948 5322 13960
rect 6825 13957 6837 13960
rect 6871 13957 6883 13991
rect 6825 13951 6883 13957
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 1946 13920 1952 13932
rect 1719 13892 1952 13920
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 1946 13880 1952 13892
rect 2004 13880 2010 13932
rect 5442 13920 5448 13932
rect 5092 13892 5448 13920
rect 5092 13861 5120 13892
rect 5442 13880 5448 13892
rect 5500 13880 5506 13932
rect 6733 13923 6791 13929
rect 6733 13889 6745 13923
rect 6779 13889 6791 13923
rect 6733 13883 6791 13889
rect 5077 13855 5135 13861
rect 5077 13821 5089 13855
rect 5123 13821 5135 13855
rect 5077 13815 5135 13821
rect 5166 13812 5172 13864
rect 5224 13852 5230 13864
rect 5261 13855 5319 13861
rect 5261 13852 5273 13855
rect 5224 13824 5273 13852
rect 5224 13812 5230 13824
rect 5261 13821 5273 13824
rect 5307 13821 5319 13855
rect 5261 13815 5319 13821
rect 5460 13784 5488 13880
rect 5534 13812 5540 13864
rect 5592 13852 5598 13864
rect 6089 13855 6147 13861
rect 6089 13852 6101 13855
rect 5592 13824 6101 13852
rect 5592 13812 5598 13824
rect 6089 13821 6101 13824
rect 6135 13852 6147 13855
rect 6748 13852 6776 13883
rect 6932 13864 6960 14028
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 7392 14028 7972 14056
rect 7098 13948 7104 14000
rect 7156 13988 7162 14000
rect 7392 13988 7420 14028
rect 7156 13960 7420 13988
rect 7156 13948 7162 13960
rect 7558 13948 7564 14000
rect 7616 13948 7622 14000
rect 7653 13991 7711 13997
rect 7653 13957 7665 13991
rect 7699 13988 7711 13991
rect 7834 13988 7840 14000
rect 7699 13960 7840 13988
rect 7699 13957 7711 13960
rect 7653 13951 7711 13957
rect 7834 13948 7840 13960
rect 7892 13948 7898 14000
rect 7944 13988 7972 14028
rect 8478 14016 8484 14068
rect 8536 14056 8542 14068
rect 9309 14059 9367 14065
rect 9309 14056 9321 14059
rect 8536 14028 9321 14056
rect 8536 14016 8542 14028
rect 9309 14025 9321 14028
rect 9355 14025 9367 14059
rect 9309 14019 9367 14025
rect 10318 14016 10324 14068
rect 10376 14056 10382 14068
rect 10505 14059 10563 14065
rect 10505 14056 10517 14059
rect 10376 14028 10517 14056
rect 10376 14016 10382 14028
rect 10505 14025 10517 14028
rect 10551 14056 10563 14059
rect 11238 14056 11244 14068
rect 10551 14028 11244 14056
rect 10551 14025 10563 14028
rect 10505 14019 10563 14025
rect 11238 14016 11244 14028
rect 11296 14016 11302 14068
rect 12084 14028 14412 14056
rect 8846 13988 8852 14000
rect 7944 13960 8852 13988
rect 8846 13948 8852 13960
rect 8904 13948 8910 14000
rect 9217 13991 9275 13997
rect 9217 13957 9229 13991
rect 9263 13988 9275 13991
rect 10134 13988 10140 14000
rect 9263 13960 10140 13988
rect 9263 13957 9275 13960
rect 9217 13951 9275 13957
rect 10134 13948 10140 13960
rect 10192 13988 10198 14000
rect 10686 13988 10692 14000
rect 10192 13960 10692 13988
rect 10192 13948 10198 13960
rect 10686 13948 10692 13960
rect 10744 13948 10750 14000
rect 7576 13920 7604 13948
rect 7745 13923 7803 13929
rect 7745 13920 7757 13923
rect 7576 13892 7757 13920
rect 7745 13889 7757 13892
rect 7791 13889 7803 13923
rect 7745 13883 7803 13889
rect 8386 13880 8392 13932
rect 8444 13920 8450 13932
rect 9490 13920 9496 13932
rect 8444 13892 9496 13920
rect 8444 13880 8450 13892
rect 9490 13880 9496 13892
rect 9548 13880 9554 13932
rect 9674 13920 9680 13932
rect 9635 13892 9680 13920
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 9858 13880 9864 13932
rect 9916 13920 9922 13932
rect 11057 13923 11115 13929
rect 11057 13920 11069 13923
rect 9916 13892 11069 13920
rect 9916 13880 9922 13892
rect 6135 13824 6776 13852
rect 6135 13821 6147 13824
rect 6089 13815 6147 13821
rect 6914 13812 6920 13864
rect 6972 13852 6978 13864
rect 7837 13855 7895 13861
rect 6972 13824 7065 13852
rect 6972 13812 6978 13824
rect 7837 13821 7849 13855
rect 7883 13821 7895 13855
rect 7837 13815 7895 13821
rect 7852 13784 7880 13815
rect 7926 13812 7932 13864
rect 7984 13852 7990 13864
rect 10244 13861 10272 13892
rect 11057 13889 11069 13892
rect 11103 13920 11115 13923
rect 12084 13920 12112 14028
rect 12158 13948 12164 14000
rect 12216 13988 12222 14000
rect 14384 13988 14412 14028
rect 14458 14016 14464 14068
rect 14516 14056 14522 14068
rect 14516 14028 16804 14056
rect 14516 14016 14522 14028
rect 14918 13988 14924 14000
rect 12216 13960 13676 13988
rect 14384 13960 14924 13988
rect 12216 13948 12222 13960
rect 12526 13929 12532 13932
rect 12520 13920 12532 13929
rect 11103 13892 12112 13920
rect 12487 13892 12532 13920
rect 11103 13889 11115 13892
rect 11057 13883 11115 13889
rect 12520 13883 12532 13892
rect 12526 13880 12532 13883
rect 12584 13880 12590 13932
rect 12894 13880 12900 13932
rect 12952 13920 12958 13932
rect 12952 13892 13308 13920
rect 12952 13880 12958 13892
rect 9769 13855 9827 13861
rect 9769 13852 9781 13855
rect 7984 13824 9781 13852
rect 7984 13812 7990 13824
rect 9769 13821 9781 13824
rect 9815 13821 9827 13855
rect 9769 13815 9827 13821
rect 9953 13855 10011 13861
rect 9953 13821 9965 13855
rect 9999 13821 10011 13855
rect 9953 13815 10011 13821
rect 10229 13855 10287 13861
rect 10229 13821 10241 13855
rect 10275 13821 10287 13855
rect 10229 13815 10287 13821
rect 10413 13855 10471 13861
rect 10413 13821 10425 13855
rect 10459 13852 10471 13855
rect 10686 13852 10692 13864
rect 10459 13824 10692 13852
rect 10459 13821 10471 13824
rect 10413 13815 10471 13821
rect 5460 13756 7880 13784
rect 9968 13784 9996 13815
rect 10686 13812 10692 13824
rect 10744 13812 10750 13864
rect 12253 13855 12311 13861
rect 12253 13821 12265 13855
rect 12299 13821 12311 13855
rect 13280 13852 13308 13892
rect 13648 13852 13676 13960
rect 14918 13948 14924 13960
rect 14976 13948 14982 14000
rect 16776 13988 16804 14028
rect 17494 14016 17500 14068
rect 17552 14056 17558 14068
rect 18141 14059 18199 14065
rect 18141 14056 18153 14059
rect 17552 14028 18153 14056
rect 17552 14016 17558 14028
rect 18141 14025 18153 14028
rect 18187 14025 18199 14059
rect 18141 14019 18199 14025
rect 21266 14016 21272 14068
rect 21324 14056 21330 14068
rect 21542 14056 21548 14068
rect 21324 14028 21548 14056
rect 21324 14016 21330 14028
rect 21542 14016 21548 14028
rect 21600 14016 21606 14068
rect 16914 13991 16972 13997
rect 16914 13988 16926 13991
rect 15028 13960 16712 13988
rect 16776 13960 16926 13988
rect 13814 13880 13820 13932
rect 13872 13920 13878 13932
rect 15028 13929 15056 13960
rect 16684 13929 16712 13960
rect 16914 13957 16926 13960
rect 16960 13957 16972 13991
rect 16914 13951 16972 13957
rect 15013 13923 15071 13929
rect 15013 13920 15025 13923
rect 13872 13892 15025 13920
rect 13872 13880 13878 13892
rect 15013 13889 15025 13892
rect 15059 13889 15071 13923
rect 15269 13923 15327 13929
rect 15269 13920 15281 13923
rect 15013 13883 15071 13889
rect 15120 13892 15281 13920
rect 15120 13852 15148 13892
rect 15269 13889 15281 13892
rect 15315 13889 15327 13923
rect 15269 13883 15327 13889
rect 16669 13923 16727 13929
rect 16669 13889 16681 13923
rect 16715 13920 16727 13923
rect 17310 13920 17316 13932
rect 16715 13892 17316 13920
rect 16715 13889 16727 13892
rect 16669 13883 16727 13889
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 18322 13880 18328 13932
rect 18380 13920 18386 13932
rect 19254 13923 19312 13929
rect 19254 13920 19266 13923
rect 18380 13892 19266 13920
rect 18380 13880 18386 13892
rect 19254 13889 19266 13892
rect 19300 13889 19312 13923
rect 19254 13883 19312 13889
rect 20254 13880 20260 13932
rect 20312 13920 20318 13932
rect 20421 13923 20479 13929
rect 20421 13920 20433 13923
rect 20312 13892 20433 13920
rect 20312 13880 20318 13892
rect 20421 13889 20433 13892
rect 20467 13889 20479 13923
rect 20421 13883 20479 13889
rect 13280 13824 13584 13852
rect 13648 13824 15148 13852
rect 12253 13815 12311 13821
rect 10778 13784 10784 13796
rect 9968 13756 10784 13784
rect 10778 13744 10784 13756
rect 10836 13744 10842 13796
rect 1486 13716 1492 13728
rect 1447 13688 1492 13716
rect 1486 13676 1492 13688
rect 1544 13676 1550 13728
rect 7650 13676 7656 13728
rect 7708 13716 7714 13728
rect 10594 13716 10600 13728
rect 7708 13688 10600 13716
rect 7708 13676 7714 13688
rect 10594 13676 10600 13688
rect 10652 13676 10658 13728
rect 10870 13716 10876 13728
rect 10831 13688 10876 13716
rect 10870 13676 10876 13688
rect 10928 13676 10934 13728
rect 12268 13716 12296 13815
rect 13556 13784 13584 13824
rect 17954 13812 17960 13864
rect 18012 13852 18018 13864
rect 19518 13852 19524 13864
rect 18012 13824 18092 13852
rect 19479 13824 19524 13852
rect 18012 13812 18018 13824
rect 13633 13787 13691 13793
rect 13633 13784 13645 13787
rect 13556 13756 13645 13784
rect 13633 13753 13645 13756
rect 13679 13753 13691 13787
rect 13814 13784 13820 13796
rect 13775 13756 13820 13784
rect 13633 13747 13691 13753
rect 13814 13744 13820 13756
rect 13872 13744 13878 13796
rect 16022 13744 16028 13796
rect 16080 13784 16086 13796
rect 18064 13793 18092 13824
rect 19518 13812 19524 13824
rect 19576 13852 19582 13864
rect 19613 13855 19671 13861
rect 19613 13852 19625 13855
rect 19576 13824 19625 13852
rect 19576 13812 19582 13824
rect 19613 13821 19625 13824
rect 19659 13852 19671 13855
rect 20165 13855 20223 13861
rect 20165 13852 20177 13855
rect 19659 13824 20177 13852
rect 19659 13821 19671 13824
rect 19613 13815 19671 13821
rect 20165 13821 20177 13824
rect 20211 13821 20223 13855
rect 20165 13815 20223 13821
rect 16393 13787 16451 13793
rect 16393 13784 16405 13787
rect 16080 13756 16405 13784
rect 16080 13744 16086 13756
rect 16393 13753 16405 13756
rect 16439 13753 16451 13787
rect 16393 13747 16451 13753
rect 18049 13787 18107 13793
rect 18049 13753 18061 13787
rect 18095 13753 18107 13787
rect 18049 13747 18107 13753
rect 12618 13716 12624 13728
rect 12268 13688 12624 13716
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 4430 13472 4436 13524
rect 4488 13512 4494 13524
rect 4525 13515 4583 13521
rect 4525 13512 4537 13515
rect 4488 13484 4537 13512
rect 4488 13472 4494 13484
rect 4525 13481 4537 13484
rect 4571 13481 4583 13515
rect 4525 13475 4583 13481
rect 5626 13472 5632 13524
rect 5684 13512 5690 13524
rect 7926 13512 7932 13524
rect 5684 13484 7512 13512
rect 7887 13484 7932 13512
rect 5684 13472 5690 13484
rect 5350 13404 5356 13456
rect 5408 13444 5414 13456
rect 7098 13444 7104 13456
rect 5408 13416 6684 13444
rect 7059 13416 7104 13444
rect 5408 13404 5414 13416
rect 6178 13376 6184 13388
rect 6139 13348 6184 13376
rect 6178 13336 6184 13348
rect 6236 13336 6242 13388
rect 6454 13376 6460 13388
rect 6415 13348 6460 13376
rect 6454 13336 6460 13348
rect 6512 13336 6518 13388
rect 6656 13385 6684 13416
rect 7098 13404 7104 13416
rect 7156 13404 7162 13456
rect 6641 13379 6699 13385
rect 6641 13345 6653 13379
rect 6687 13345 6699 13379
rect 7374 13376 7380 13388
rect 7335 13348 7380 13376
rect 6641 13339 6699 13345
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 7484 13385 7512 13484
rect 7926 13472 7932 13484
rect 7984 13472 7990 13524
rect 9214 13472 9220 13524
rect 9272 13512 9278 13524
rect 9401 13515 9459 13521
rect 9401 13512 9413 13515
rect 9272 13484 9413 13512
rect 9272 13472 9278 13484
rect 9401 13481 9413 13484
rect 9447 13481 9459 13515
rect 11882 13512 11888 13524
rect 9401 13475 9459 13481
rect 9508 13484 11888 13512
rect 8021 13447 8079 13453
rect 8021 13413 8033 13447
rect 8067 13413 8079 13447
rect 8021 13407 8079 13413
rect 7469 13379 7527 13385
rect 7469 13345 7481 13379
rect 7515 13345 7527 13379
rect 7469 13339 7527 13345
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 2041 13311 2099 13317
rect 1719 13280 1900 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 1486 13172 1492 13184
rect 1447 13144 1492 13172
rect 1486 13132 1492 13144
rect 1544 13132 1550 13184
rect 1872 13181 1900 13280
rect 2041 13277 2053 13311
rect 2087 13308 2099 13311
rect 3142 13308 3148 13320
rect 2087 13280 3148 13308
rect 2087 13277 2099 13280
rect 2041 13271 2099 13277
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13308 4767 13311
rect 8036 13308 8064 13407
rect 8754 13404 8760 13456
rect 8812 13444 8818 13456
rect 9508 13444 9536 13484
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 12406 13484 13584 13512
rect 12406 13444 12434 13484
rect 8812 13416 9536 13444
rect 10060 13416 12434 13444
rect 8812 13404 8818 13416
rect 8662 13376 8668 13388
rect 8623 13348 8668 13376
rect 8662 13336 8668 13348
rect 8720 13336 8726 13388
rect 10060 13385 10088 13416
rect 10045 13379 10103 13385
rect 9324 13348 9904 13376
rect 9324 13308 9352 13348
rect 4755 13280 8064 13308
rect 8128 13280 9352 13308
rect 4755 13277 4767 13280
rect 4709 13271 4767 13277
rect 5718 13200 5724 13252
rect 5776 13240 5782 13252
rect 6733 13243 6791 13249
rect 6733 13240 6745 13243
rect 5776 13212 6745 13240
rect 5776 13200 5782 13212
rect 6733 13209 6745 13212
rect 6779 13209 6791 13243
rect 6733 13203 6791 13209
rect 6822 13200 6828 13252
rect 6880 13240 6886 13252
rect 8128 13240 8156 13280
rect 9398 13268 9404 13320
rect 9456 13308 9462 13320
rect 9769 13311 9827 13317
rect 9769 13308 9781 13311
rect 9456 13280 9781 13308
rect 9456 13268 9462 13280
rect 9769 13277 9781 13280
rect 9815 13277 9827 13311
rect 9876 13308 9904 13348
rect 10045 13345 10057 13379
rect 10091 13345 10103 13379
rect 10781 13379 10839 13385
rect 10045 13339 10103 13345
rect 10520 13348 10732 13376
rect 10520 13308 10548 13348
rect 10704 13317 10732 13348
rect 10781 13345 10793 13379
rect 10827 13376 10839 13379
rect 10962 13376 10968 13388
rect 10827 13348 10968 13376
rect 10827 13345 10839 13348
rect 10781 13339 10839 13345
rect 10962 13336 10968 13348
rect 11020 13336 11026 13388
rect 11701 13379 11759 13385
rect 11701 13345 11713 13379
rect 11747 13376 11759 13379
rect 11974 13376 11980 13388
rect 11747 13348 11980 13376
rect 11747 13345 11759 13348
rect 11701 13339 11759 13345
rect 11974 13336 11980 13348
rect 12032 13376 12038 13388
rect 12434 13376 12440 13388
rect 12032 13348 12440 13376
rect 12032 13336 12038 13348
rect 12434 13336 12440 13348
rect 12492 13336 12498 13388
rect 9876 13280 10548 13308
rect 10689 13311 10747 13317
rect 9769 13271 9827 13277
rect 10689 13277 10701 13311
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 10870 13268 10876 13320
rect 10928 13268 10934 13320
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13308 11575 13311
rect 11606 13308 11612 13320
rect 11563 13280 11612 13308
rect 11563 13277 11575 13280
rect 11517 13271 11575 13277
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 12529 13311 12587 13317
rect 12529 13277 12541 13311
rect 12575 13308 12587 13311
rect 12618 13308 12624 13320
rect 12575 13280 12624 13308
rect 12575 13277 12587 13280
rect 12529 13271 12587 13277
rect 12618 13268 12624 13280
rect 12676 13268 12682 13320
rect 12802 13317 12808 13320
rect 12796 13308 12808 13317
rect 12763 13280 12808 13308
rect 12796 13271 12808 13280
rect 12802 13268 12808 13271
rect 12860 13268 12866 13320
rect 13556 13308 13584 13484
rect 17310 13472 17316 13524
rect 17368 13512 17374 13524
rect 17586 13512 17592 13524
rect 17368 13484 17592 13512
rect 17368 13472 17374 13484
rect 15194 13404 15200 13456
rect 15252 13444 15258 13456
rect 16117 13447 16175 13453
rect 16117 13444 16129 13447
rect 15252 13416 16129 13444
rect 15252 13404 15258 13416
rect 16117 13413 16129 13416
rect 16163 13413 16175 13447
rect 16117 13407 16175 13413
rect 17512 13385 17540 13484
rect 17586 13472 17592 13484
rect 17644 13512 17650 13524
rect 19245 13515 19303 13521
rect 19245 13512 19257 13515
rect 17644 13484 19257 13512
rect 17644 13472 17650 13484
rect 19245 13481 19257 13484
rect 19291 13512 19303 13515
rect 19518 13512 19524 13524
rect 19291 13484 19524 13512
rect 19291 13481 19303 13484
rect 19245 13475 19303 13481
rect 19518 13472 19524 13484
rect 19576 13472 19582 13524
rect 20898 13512 20904 13524
rect 20364 13484 20904 13512
rect 18966 13444 18972 13456
rect 18927 13416 18972 13444
rect 18966 13404 18972 13416
rect 19024 13444 19030 13456
rect 20364 13444 20392 13484
rect 20898 13472 20904 13484
rect 20956 13472 20962 13524
rect 19024 13416 20392 13444
rect 19024 13404 19030 13416
rect 17497 13379 17555 13385
rect 17497 13345 17509 13379
rect 17543 13376 17555 13379
rect 17589 13379 17647 13385
rect 17589 13376 17601 13379
rect 17543 13348 17601 13376
rect 17543 13345 17555 13348
rect 17497 13339 17555 13345
rect 17589 13345 17601 13348
rect 17635 13345 17647 13379
rect 17589 13339 17647 13345
rect 17230 13311 17288 13317
rect 17230 13308 17242 13311
rect 13556 13280 17242 13308
rect 17230 13277 17242 13280
rect 17276 13308 17288 13311
rect 17678 13308 17684 13320
rect 17276 13280 17684 13308
rect 17276 13277 17288 13280
rect 17230 13271 17288 13277
rect 17678 13268 17684 13280
rect 17736 13268 17742 13320
rect 21174 13268 21180 13320
rect 21232 13308 21238 13320
rect 21269 13311 21327 13317
rect 21269 13308 21281 13311
rect 21232 13280 21281 13308
rect 21232 13268 21238 13280
rect 21269 13277 21281 13280
rect 21315 13308 21327 13311
rect 21453 13311 21511 13317
rect 21453 13308 21465 13311
rect 21315 13280 21465 13308
rect 21315 13277 21327 13280
rect 21269 13271 21327 13277
rect 21453 13277 21465 13280
rect 21499 13277 21511 13311
rect 21453 13271 21511 13277
rect 6880 13212 8156 13240
rect 8481 13243 8539 13249
rect 6880 13200 6886 13212
rect 8481 13209 8493 13243
rect 8527 13240 8539 13243
rect 9950 13240 9956 13252
rect 8527 13212 9956 13240
rect 8527 13209 8539 13212
rect 8481 13203 8539 13209
rect 9950 13200 9956 13212
rect 10008 13200 10014 13252
rect 10597 13243 10655 13249
rect 10597 13209 10609 13243
rect 10643 13240 10655 13243
rect 10888 13240 10916 13268
rect 10643 13212 10916 13240
rect 10643 13209 10655 13212
rect 10597 13203 10655 13209
rect 11790 13200 11796 13252
rect 11848 13240 11854 13252
rect 17834 13243 17892 13249
rect 17834 13240 17846 13243
rect 11848 13212 17846 13240
rect 11848 13200 11854 13212
rect 17834 13209 17846 13212
rect 17880 13240 17892 13243
rect 18046 13240 18052 13252
rect 17880 13212 18052 13240
rect 17880 13209 17892 13212
rect 17834 13203 17892 13209
rect 18046 13200 18052 13212
rect 18104 13200 18110 13252
rect 20162 13200 20168 13252
rect 20220 13240 20226 13252
rect 21002 13243 21060 13249
rect 21002 13240 21014 13243
rect 20220 13212 21014 13240
rect 20220 13200 20226 13212
rect 21002 13209 21014 13212
rect 21048 13209 21060 13243
rect 21002 13203 21060 13209
rect 1857 13175 1915 13181
rect 1857 13141 1869 13175
rect 1903 13141 1915 13175
rect 1857 13135 1915 13141
rect 7558 13132 7564 13184
rect 7616 13172 7622 13184
rect 8386 13172 8392 13184
rect 7616 13144 7661 13172
rect 8347 13144 8392 13172
rect 7616 13132 7622 13144
rect 8386 13132 8392 13144
rect 8444 13132 8450 13184
rect 9858 13172 9864 13184
rect 9819 13144 9864 13172
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 10229 13175 10287 13181
rect 10229 13141 10241 13175
rect 10275 13172 10287 13175
rect 10410 13172 10416 13184
rect 10275 13144 10416 13172
rect 10275 13141 10287 13144
rect 10229 13135 10287 13141
rect 10410 13132 10416 13144
rect 10468 13132 10474 13184
rect 10870 13132 10876 13184
rect 10928 13172 10934 13184
rect 11057 13175 11115 13181
rect 11057 13172 11069 13175
rect 10928 13144 11069 13172
rect 10928 13132 10934 13144
rect 11057 13141 11069 13144
rect 11103 13141 11115 13175
rect 11057 13135 11115 13141
rect 11238 13132 11244 13184
rect 11296 13172 11302 13184
rect 11425 13175 11483 13181
rect 11425 13172 11437 13175
rect 11296 13144 11437 13172
rect 11296 13132 11302 13144
rect 11425 13141 11437 13144
rect 11471 13141 11483 13175
rect 11425 13135 11483 13141
rect 13262 13132 13268 13184
rect 13320 13172 13326 13184
rect 13909 13175 13967 13181
rect 13909 13172 13921 13175
rect 13320 13144 13921 13172
rect 13320 13132 13326 13144
rect 13909 13141 13921 13144
rect 13955 13141 13967 13175
rect 14090 13172 14096 13184
rect 14051 13144 14096 13172
rect 13909 13135 13967 13141
rect 14090 13132 14096 13144
rect 14148 13132 14154 13184
rect 15930 13172 15936 13184
rect 15891 13144 15936 13172
rect 15930 13132 15936 13144
rect 15988 13132 15994 13184
rect 19886 13172 19892 13184
rect 19847 13144 19892 13172
rect 19886 13132 19892 13144
rect 19944 13132 19950 13184
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 1857 12971 1915 12977
rect 1857 12937 1869 12971
rect 1903 12937 1915 12971
rect 3142 12968 3148 12980
rect 3103 12940 3148 12968
rect 1857 12931 1915 12937
rect 1872 12900 1900 12931
rect 3142 12928 3148 12940
rect 3200 12928 3206 12980
rect 4246 12968 4252 12980
rect 4207 12940 4252 12968
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 5077 12971 5135 12977
rect 4356 12940 5028 12968
rect 4154 12900 4160 12912
rect 1872 12872 4160 12900
rect 4154 12860 4160 12872
rect 4212 12860 4218 12912
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 1670 12832 1676 12844
rect 1631 12804 1676 12832
rect 1670 12792 1676 12804
rect 1728 12832 1734 12844
rect 1949 12835 2007 12841
rect 1949 12832 1961 12835
rect 1728 12804 1961 12832
rect 1728 12792 1734 12804
rect 1949 12801 1961 12804
rect 1995 12801 2007 12835
rect 1949 12795 2007 12801
rect 3329 12835 3387 12841
rect 3329 12801 3341 12835
rect 3375 12801 3387 12835
rect 3329 12795 3387 12801
rect 1412 12764 1440 12792
rect 2133 12767 2191 12773
rect 2133 12764 2145 12767
rect 1412 12736 2145 12764
rect 2133 12733 2145 12736
rect 2179 12733 2191 12767
rect 3344 12764 3372 12795
rect 3878 12792 3884 12844
rect 3936 12832 3942 12844
rect 4356 12832 4384 12940
rect 5000 12900 5028 12940
rect 5077 12937 5089 12971
rect 5123 12968 5135 12971
rect 5445 12971 5503 12977
rect 5445 12968 5457 12971
rect 5123 12940 5457 12968
rect 5123 12937 5135 12940
rect 5077 12931 5135 12937
rect 5445 12937 5457 12940
rect 5491 12937 5503 12971
rect 5445 12931 5503 12937
rect 5905 12971 5963 12977
rect 5905 12937 5917 12971
rect 5951 12968 5963 12971
rect 6365 12971 6423 12977
rect 6365 12968 6377 12971
rect 5951 12940 6377 12968
rect 5951 12937 5963 12940
rect 5905 12931 5963 12937
rect 6365 12937 6377 12940
rect 6411 12937 6423 12971
rect 6365 12931 6423 12937
rect 6454 12928 6460 12980
rect 6512 12968 6518 12980
rect 6730 12968 6736 12980
rect 6512 12940 6736 12968
rect 6512 12928 6518 12940
rect 6730 12928 6736 12940
rect 6788 12928 6794 12980
rect 7285 12971 7343 12977
rect 7285 12937 7297 12971
rect 7331 12968 7343 12971
rect 7331 12940 8340 12968
rect 7331 12937 7343 12940
rect 7285 12931 7343 12937
rect 6825 12903 6883 12909
rect 6825 12900 6837 12903
rect 5000 12872 6837 12900
rect 6825 12869 6837 12872
rect 6871 12869 6883 12903
rect 6825 12863 6883 12869
rect 3936 12804 4384 12832
rect 4433 12835 4491 12841
rect 3936 12792 3942 12804
rect 4433 12801 4445 12835
rect 4479 12832 4491 12835
rect 4982 12832 4988 12844
rect 4479 12804 4844 12832
rect 4943 12804 4988 12832
rect 4479 12801 4491 12804
rect 4433 12795 4491 12801
rect 3344 12736 4660 12764
rect 2133 12727 2191 12733
rect 1581 12699 1639 12705
rect 1581 12665 1593 12699
rect 1627 12696 1639 12699
rect 4522 12696 4528 12708
rect 1627 12668 4528 12696
rect 1627 12665 1639 12668
rect 1581 12659 1639 12665
rect 4522 12656 4528 12668
rect 4580 12656 4586 12708
rect 4632 12705 4660 12736
rect 4617 12699 4675 12705
rect 4617 12665 4629 12699
rect 4663 12665 4675 12699
rect 4816 12696 4844 12804
rect 4982 12792 4988 12804
rect 5040 12792 5046 12844
rect 5810 12832 5816 12844
rect 5771 12804 5816 12832
rect 5810 12792 5816 12804
rect 5868 12792 5874 12844
rect 7300 12776 7328 12931
rect 7650 12860 7656 12912
rect 7708 12900 7714 12912
rect 7929 12903 7987 12909
rect 7929 12900 7941 12903
rect 7708 12872 7941 12900
rect 7708 12860 7714 12872
rect 7929 12869 7941 12872
rect 7975 12869 7987 12903
rect 8312 12900 8340 12940
rect 8386 12928 8392 12980
rect 8444 12968 8450 12980
rect 8573 12971 8631 12977
rect 8573 12968 8585 12971
rect 8444 12940 8585 12968
rect 8444 12928 8450 12940
rect 8573 12937 8585 12940
rect 8619 12937 8631 12971
rect 8573 12931 8631 12937
rect 9582 12928 9588 12980
rect 9640 12968 9646 12980
rect 9953 12971 10011 12977
rect 9953 12968 9965 12971
rect 9640 12940 9965 12968
rect 9640 12928 9646 12940
rect 9953 12937 9965 12940
rect 9999 12937 10011 12971
rect 10410 12968 10416 12980
rect 10371 12940 10416 12968
rect 9953 12931 10011 12937
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 10870 12928 10876 12980
rect 10928 12968 10934 12980
rect 13262 12968 13268 12980
rect 10928 12940 13268 12968
rect 10928 12928 10934 12940
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 14182 12968 14188 12980
rect 13924 12940 14188 12968
rect 8312 12872 10456 12900
rect 7929 12863 7987 12869
rect 7561 12835 7619 12841
rect 7561 12801 7573 12835
rect 7607 12832 7619 12835
rect 8021 12835 8079 12841
rect 8021 12832 8033 12835
rect 7607 12804 8033 12832
rect 7607 12801 7619 12804
rect 7561 12795 7619 12801
rect 8021 12801 8033 12804
rect 8067 12801 8079 12835
rect 8021 12795 8079 12801
rect 8386 12792 8392 12844
rect 8444 12832 8450 12844
rect 8754 12832 8760 12844
rect 8444 12804 8760 12832
rect 8444 12792 8450 12804
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 8941 12835 8999 12841
rect 8941 12801 8953 12835
rect 8987 12832 8999 12835
rect 9306 12832 9312 12844
rect 8987 12804 9312 12832
rect 8987 12801 8999 12804
rect 8941 12795 8999 12801
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 9858 12792 9864 12844
rect 9916 12832 9922 12844
rect 10321 12835 10379 12841
rect 10321 12832 10333 12835
rect 9916 12804 10333 12832
rect 9916 12792 9922 12804
rect 10321 12801 10333 12804
rect 10367 12801 10379 12835
rect 10428 12832 10456 12872
rect 10594 12860 10600 12912
rect 10652 12900 10658 12912
rect 13538 12900 13544 12912
rect 10652 12872 13544 12900
rect 10652 12860 10658 12872
rect 13538 12860 13544 12872
rect 13596 12860 13602 12912
rect 13837 12903 13895 12909
rect 13837 12869 13849 12903
rect 13883 12900 13895 12903
rect 13924 12900 13952 12940
rect 14182 12928 14188 12940
rect 14240 12928 14246 12980
rect 17586 12928 17592 12980
rect 17644 12968 17650 12980
rect 17862 12968 17868 12980
rect 17644 12940 17868 12968
rect 17644 12928 17650 12940
rect 17862 12928 17868 12940
rect 17920 12968 17926 12980
rect 18141 12971 18199 12977
rect 18141 12968 18153 12971
rect 17920 12940 18153 12968
rect 17920 12928 17926 12940
rect 18141 12937 18153 12940
rect 18187 12968 18199 12971
rect 18325 12971 18383 12977
rect 18325 12968 18337 12971
rect 18187 12940 18337 12968
rect 18187 12937 18199 12940
rect 18141 12931 18199 12937
rect 18325 12937 18337 12940
rect 18371 12968 18383 12971
rect 20809 12971 20867 12977
rect 20809 12968 20821 12971
rect 18371 12940 20821 12968
rect 18371 12937 18383 12940
rect 18325 12931 18383 12937
rect 15657 12903 15715 12909
rect 15657 12900 15669 12903
rect 13883 12872 13952 12900
rect 14292 12872 15669 12900
rect 13883 12869 13895 12872
rect 13837 12863 13895 12869
rect 14292 12844 14320 12872
rect 10428 12804 14044 12832
rect 10321 12795 10379 12801
rect 5258 12764 5264 12776
rect 5219 12736 5264 12764
rect 5258 12724 5264 12736
rect 5316 12724 5322 12776
rect 6089 12767 6147 12773
rect 6089 12733 6101 12767
rect 6135 12764 6147 12767
rect 6270 12764 6276 12776
rect 6135 12736 6276 12764
rect 6135 12733 6147 12736
rect 6089 12727 6147 12733
rect 6270 12724 6276 12736
rect 6328 12764 6334 12776
rect 6546 12764 6552 12776
rect 6328 12736 6552 12764
rect 6328 12724 6334 12736
rect 6546 12724 6552 12736
rect 6604 12724 6610 12776
rect 7009 12767 7067 12773
rect 7009 12733 7021 12767
rect 7055 12764 7067 12767
rect 7282 12764 7288 12776
rect 7055 12736 7288 12764
rect 7055 12733 7067 12736
rect 7009 12727 7067 12733
rect 7282 12724 7288 12736
rect 7340 12724 7346 12776
rect 7374 12724 7380 12776
rect 7432 12764 7438 12776
rect 7745 12767 7803 12773
rect 7745 12764 7757 12767
rect 7432 12736 7757 12764
rect 7432 12724 7438 12736
rect 7745 12733 7757 12736
rect 7791 12733 7803 12767
rect 7745 12727 7803 12733
rect 7944 12736 8340 12764
rect 7944 12696 7972 12736
rect 4816 12668 7972 12696
rect 4617 12659 4675 12665
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4890 12628 4896 12640
rect 4212 12600 4896 12628
rect 4212 12588 4218 12600
rect 4890 12588 4896 12600
rect 4948 12588 4954 12640
rect 6914 12588 6920 12640
rect 6972 12628 6978 12640
rect 8018 12628 8024 12640
rect 6972 12600 8024 12628
rect 6972 12588 6978 12600
rect 8018 12588 8024 12600
rect 8076 12588 8082 12640
rect 8312 12628 8340 12736
rect 8570 12724 8576 12776
rect 8628 12764 8634 12776
rect 9033 12767 9091 12773
rect 9033 12764 9045 12767
rect 8628 12736 9045 12764
rect 8628 12724 8634 12736
rect 9033 12733 9045 12736
rect 9079 12733 9091 12767
rect 9033 12727 9091 12733
rect 9217 12767 9275 12773
rect 9217 12733 9229 12767
rect 9263 12764 9275 12767
rect 10597 12767 10655 12773
rect 9263 12736 10548 12764
rect 9263 12733 9275 12736
rect 9217 12727 9275 12733
rect 8389 12699 8447 12705
rect 8389 12665 8401 12699
rect 8435 12696 8447 12699
rect 9674 12696 9680 12708
rect 8435 12668 9680 12696
rect 8435 12665 8447 12668
rect 8389 12659 8447 12665
rect 9674 12656 9680 12668
rect 9732 12656 9738 12708
rect 10520 12696 10548 12736
rect 10597 12733 10609 12767
rect 10643 12764 10655 12767
rect 12158 12764 12164 12776
rect 10643 12736 12164 12764
rect 10643 12733 10655 12736
rect 10597 12727 10655 12733
rect 12158 12724 12164 12736
rect 12216 12724 12222 12776
rect 14016 12764 14044 12804
rect 14090 12792 14096 12844
rect 14148 12832 14154 12844
rect 14274 12832 14280 12844
rect 14148 12804 14280 12832
rect 14148 12792 14154 12804
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 14826 12832 14832 12844
rect 14568 12804 14832 12832
rect 14568 12764 14596 12804
rect 14826 12792 14832 12804
rect 14884 12792 14890 12844
rect 15286 12832 15292 12844
rect 15344 12841 15350 12844
rect 15580 12841 15608 12872
rect 15657 12869 15669 12872
rect 15703 12900 15715 12903
rect 15930 12900 15936 12912
rect 15703 12872 15936 12900
rect 15703 12869 15715 12872
rect 15657 12863 15715 12869
rect 15930 12860 15936 12872
rect 15988 12860 15994 12912
rect 16390 12860 16396 12912
rect 16448 12900 16454 12912
rect 16914 12903 16972 12909
rect 16914 12900 16926 12903
rect 16448 12872 16926 12900
rect 16448 12860 16454 12872
rect 16914 12869 16926 12872
rect 16960 12869 16972 12903
rect 16914 12863 16972 12869
rect 19886 12860 19892 12912
rect 19944 12900 19950 12912
rect 20070 12900 20076 12912
rect 19944 12872 20076 12900
rect 19944 12860 19950 12872
rect 20070 12860 20076 12872
rect 20128 12900 20134 12912
rect 20450 12903 20508 12909
rect 20450 12900 20462 12903
rect 20128 12872 20462 12900
rect 20128 12860 20134 12872
rect 20450 12869 20462 12872
rect 20496 12869 20508 12903
rect 20450 12863 20508 12869
rect 15256 12804 15292 12832
rect 15286 12792 15292 12804
rect 15344 12795 15356 12841
rect 15565 12835 15623 12841
rect 15565 12801 15577 12835
rect 15611 12801 15623 12835
rect 15948 12832 15976 12860
rect 16666 12832 16672 12844
rect 15948 12804 16672 12832
rect 15565 12795 15623 12801
rect 15344 12792 15350 12795
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 20732 12841 20760 12940
rect 20809 12937 20821 12940
rect 20855 12968 20867 12971
rect 21082 12968 21088 12980
rect 20855 12940 21088 12968
rect 20855 12937 20867 12940
rect 20809 12931 20867 12937
rect 21082 12928 21088 12940
rect 21140 12968 21146 12980
rect 21266 12968 21272 12980
rect 21140 12940 21272 12968
rect 21140 12928 21146 12940
rect 21266 12928 21272 12940
rect 21324 12968 21330 12980
rect 21361 12971 21419 12977
rect 21361 12968 21373 12971
rect 21324 12940 21373 12968
rect 21324 12928 21330 12940
rect 21361 12937 21373 12940
rect 21407 12937 21419 12971
rect 21361 12931 21419 12937
rect 20717 12835 20775 12841
rect 20717 12801 20729 12835
rect 20763 12801 20775 12835
rect 20717 12795 20775 12801
rect 14016 12736 14596 12764
rect 10962 12696 10968 12708
rect 10520 12668 10968 12696
rect 10962 12656 10968 12668
rect 11020 12696 11026 12708
rect 11790 12696 11796 12708
rect 11020 12668 11796 12696
rect 11020 12656 11026 12668
rect 11790 12656 11796 12668
rect 11848 12656 11854 12708
rect 17678 12656 17684 12708
rect 17736 12696 17742 12708
rect 18049 12699 18107 12705
rect 18049 12696 18061 12699
rect 17736 12668 18061 12696
rect 17736 12656 17742 12668
rect 18049 12665 18061 12668
rect 18095 12665 18107 12699
rect 18049 12659 18107 12665
rect 8662 12628 8668 12640
rect 8312 12600 8668 12628
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 10226 12588 10232 12640
rect 10284 12628 10290 12640
rect 10594 12628 10600 12640
rect 10284 12600 10600 12628
rect 10284 12588 10290 12600
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 12618 12628 12624 12640
rect 12579 12600 12624 12628
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 12710 12588 12716 12640
rect 12768 12628 12774 12640
rect 12986 12628 12992 12640
rect 12768 12600 12992 12628
rect 12768 12588 12774 12600
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 13446 12588 13452 12640
rect 13504 12628 13510 12640
rect 14185 12631 14243 12637
rect 14185 12628 14197 12631
rect 13504 12600 14197 12628
rect 13504 12588 13510 12600
rect 14185 12597 14197 12600
rect 14231 12597 14243 12631
rect 14185 12591 14243 12597
rect 19337 12631 19395 12637
rect 19337 12597 19349 12631
rect 19383 12628 19395 12631
rect 19518 12628 19524 12640
rect 19383 12600 19524 12628
rect 19383 12597 19395 12600
rect 19337 12591 19395 12597
rect 19518 12588 19524 12600
rect 19576 12588 19582 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 1578 12384 1584 12436
rect 1636 12424 1642 12436
rect 1857 12427 1915 12433
rect 1857 12424 1869 12427
rect 1636 12396 1869 12424
rect 1636 12384 1642 12396
rect 1857 12393 1869 12396
rect 1903 12393 1915 12427
rect 1857 12387 1915 12393
rect 4062 12384 4068 12436
rect 4120 12424 4126 12436
rect 4893 12427 4951 12433
rect 4893 12424 4905 12427
rect 4120 12396 4905 12424
rect 4120 12384 4126 12396
rect 4893 12393 4905 12396
rect 4939 12393 4951 12427
rect 4893 12387 4951 12393
rect 4982 12384 4988 12436
rect 5040 12424 5046 12436
rect 5629 12427 5687 12433
rect 5629 12424 5641 12427
rect 5040 12396 5641 12424
rect 5040 12384 5046 12396
rect 5629 12393 5641 12396
rect 5675 12393 5687 12427
rect 5629 12387 5687 12393
rect 6822 12384 6828 12436
rect 6880 12424 6886 12436
rect 7098 12424 7104 12436
rect 6880 12396 7104 12424
rect 6880 12384 6886 12396
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 7469 12427 7527 12433
rect 7469 12393 7481 12427
rect 7515 12424 7527 12427
rect 7834 12424 7840 12436
rect 7515 12396 7840 12424
rect 7515 12393 7527 12396
rect 7469 12387 7527 12393
rect 7834 12384 7840 12396
rect 7892 12384 7898 12436
rect 8018 12384 8024 12436
rect 8076 12424 8082 12436
rect 8202 12424 8208 12436
rect 8076 12396 8208 12424
rect 8076 12384 8082 12396
rect 8202 12384 8208 12396
rect 8260 12384 8266 12436
rect 8570 12424 8576 12436
rect 8404 12396 8576 12424
rect 5994 12356 6000 12368
rect 5644 12328 6000 12356
rect 5644 12300 5672 12328
rect 5994 12316 6000 12328
rect 6052 12356 6058 12368
rect 8404 12365 8432 12396
rect 8570 12384 8576 12396
rect 8628 12384 8634 12436
rect 8662 12384 8668 12436
rect 8720 12424 8726 12436
rect 8941 12427 8999 12433
rect 8941 12424 8953 12427
rect 8720 12396 8953 12424
rect 8720 12384 8726 12396
rect 8941 12393 8953 12396
rect 8987 12393 8999 12427
rect 8941 12387 8999 12393
rect 9950 12384 9956 12436
rect 10008 12424 10014 12436
rect 10229 12427 10287 12433
rect 10229 12424 10241 12427
rect 10008 12396 10241 12424
rect 10008 12384 10014 12396
rect 10229 12393 10241 12396
rect 10275 12393 10287 12427
rect 10229 12387 10287 12393
rect 10778 12384 10784 12436
rect 10836 12424 10842 12436
rect 10836 12396 17724 12424
rect 10836 12384 10842 12396
rect 8389 12359 8447 12365
rect 8389 12356 8401 12359
rect 6052 12328 8401 12356
rect 6052 12316 6058 12328
rect 8389 12325 8401 12328
rect 8435 12325 8447 12359
rect 8389 12319 8447 12325
rect 9306 12316 9312 12368
rect 9364 12356 9370 12368
rect 11146 12356 11152 12368
rect 9364 12328 9720 12356
rect 9364 12316 9370 12328
rect 5626 12248 5632 12300
rect 5684 12248 5690 12300
rect 6270 12288 6276 12300
rect 6231 12260 6276 12288
rect 6270 12248 6276 12260
rect 6328 12248 6334 12300
rect 6638 12248 6644 12300
rect 6696 12288 6702 12300
rect 7374 12288 7380 12300
rect 6696 12260 7380 12288
rect 6696 12248 6702 12260
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 8110 12288 8116 12300
rect 8071 12260 8116 12288
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 8202 12248 8208 12300
rect 8260 12288 8266 12300
rect 9582 12288 9588 12300
rect 8260 12260 9444 12288
rect 9543 12260 9588 12288
rect 8260 12248 8266 12260
rect 1394 12220 1400 12232
rect 1355 12192 1400 12220
rect 1394 12180 1400 12192
rect 1452 12220 1458 12232
rect 1673 12223 1731 12229
rect 1673 12220 1685 12223
rect 1452 12192 1685 12220
rect 1452 12180 1458 12192
rect 1673 12189 1685 12192
rect 1719 12189 1731 12223
rect 1673 12183 1731 12189
rect 2041 12223 2099 12229
rect 2041 12189 2053 12223
rect 2087 12220 2099 12223
rect 3234 12220 3240 12232
rect 2087 12192 3240 12220
rect 2087 12189 2099 12192
rect 2041 12183 2099 12189
rect 3234 12180 3240 12192
rect 3292 12180 3298 12232
rect 5077 12223 5135 12229
rect 5077 12189 5089 12223
rect 5123 12220 5135 12223
rect 9306 12220 9312 12232
rect 5123 12192 9312 12220
rect 5123 12189 5135 12192
rect 5077 12183 5135 12189
rect 9306 12180 9312 12192
rect 9364 12180 9370 12232
rect 9416 12220 9444 12260
rect 9582 12248 9588 12260
rect 9640 12248 9646 12300
rect 9692 12288 9720 12328
rect 9876 12328 11152 12356
rect 9769 12291 9827 12297
rect 9769 12288 9781 12291
rect 9692 12260 9781 12288
rect 9769 12257 9781 12260
rect 9815 12257 9827 12291
rect 9769 12251 9827 12257
rect 9876 12220 9904 12328
rect 11146 12316 11152 12328
rect 11204 12316 11210 12368
rect 13722 12316 13728 12368
rect 13780 12356 13786 12368
rect 15289 12359 15347 12365
rect 15289 12356 15301 12359
rect 13780 12328 15301 12356
rect 13780 12316 13786 12328
rect 15289 12325 15301 12328
rect 15335 12325 15347 12359
rect 17696 12356 17724 12396
rect 17862 12384 17868 12436
rect 17920 12424 17926 12436
rect 18233 12427 18291 12433
rect 18233 12424 18245 12427
rect 17920 12396 18245 12424
rect 17920 12384 17926 12396
rect 18233 12393 18245 12396
rect 18279 12393 18291 12427
rect 18233 12387 18291 12393
rect 18141 12359 18199 12365
rect 18141 12356 18153 12359
rect 17696 12328 18153 12356
rect 15289 12319 15347 12325
rect 18141 12325 18153 12328
rect 18187 12325 18199 12359
rect 18141 12319 18199 12325
rect 19797 12359 19855 12365
rect 19797 12325 19809 12359
rect 19843 12325 19855 12359
rect 19797 12319 19855 12325
rect 10873 12291 10931 12297
rect 10873 12257 10885 12291
rect 10919 12288 10931 12291
rect 10962 12288 10968 12300
rect 10919 12260 10968 12288
rect 10919 12257 10931 12260
rect 10873 12251 10931 12257
rect 10962 12248 10968 12260
rect 11020 12248 11026 12300
rect 16666 12288 16672 12300
rect 16627 12260 16672 12288
rect 16666 12248 16672 12260
rect 16724 12288 16730 12300
rect 16761 12291 16819 12297
rect 16761 12288 16773 12291
rect 16724 12260 16773 12288
rect 16724 12248 16730 12260
rect 16761 12257 16773 12260
rect 16807 12257 16819 12291
rect 16761 12251 16819 12257
rect 9416 12192 9904 12220
rect 10689 12223 10747 12229
rect 10689 12189 10701 12223
rect 10735 12220 10747 12223
rect 11054 12220 11060 12232
rect 10735 12192 11060 12220
rect 10735 12189 10747 12192
rect 10689 12183 10747 12189
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 12170 12223 12228 12229
rect 12170 12220 12182 12223
rect 11348 12192 12182 12220
rect 5092 12124 6684 12152
rect 5092 12096 5120 12124
rect 1581 12087 1639 12093
rect 1581 12053 1593 12087
rect 1627 12084 1639 12087
rect 2682 12084 2688 12096
rect 1627 12056 2688 12084
rect 1627 12053 1639 12056
rect 1581 12047 1639 12053
rect 2682 12044 2688 12056
rect 2740 12044 2746 12096
rect 5074 12044 5080 12096
rect 5132 12044 5138 12096
rect 5994 12084 6000 12096
rect 5955 12056 6000 12084
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6089 12087 6147 12093
rect 6089 12053 6101 12087
rect 6135 12084 6147 12087
rect 6546 12084 6552 12096
rect 6135 12056 6552 12084
rect 6135 12053 6147 12056
rect 6089 12047 6147 12053
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 6656 12084 6684 12124
rect 7190 12112 7196 12164
rect 7248 12152 7254 12164
rect 7929 12155 7987 12161
rect 7929 12152 7941 12155
rect 7248 12124 7941 12152
rect 7248 12112 7254 12124
rect 7929 12121 7941 12124
rect 7975 12152 7987 12155
rect 8665 12155 8723 12161
rect 8665 12152 8677 12155
rect 7975 12124 8677 12152
rect 7975 12121 7987 12124
rect 7929 12115 7987 12121
rect 8665 12121 8677 12124
rect 8711 12152 8723 12155
rect 10410 12152 10416 12164
rect 8711 12124 10416 12152
rect 8711 12121 8723 12124
rect 8665 12115 8723 12121
rect 10410 12112 10416 12124
rect 10468 12112 10474 12164
rect 10778 12112 10784 12164
rect 10836 12152 10842 12164
rect 11348 12152 11376 12192
rect 12170 12189 12182 12192
rect 12216 12220 12228 12223
rect 12342 12220 12348 12232
rect 12216 12192 12348 12220
rect 12216 12189 12228 12192
rect 12170 12183 12228 12189
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12220 12495 12223
rect 12526 12220 12532 12232
rect 12483 12192 12532 12220
rect 12483 12189 12495 12192
rect 12437 12183 12495 12189
rect 12526 12180 12532 12192
rect 12584 12180 12590 12232
rect 17034 12229 17040 12232
rect 17028 12183 17040 12229
rect 17092 12220 17098 12232
rect 18156 12220 18184 12319
rect 18230 12248 18236 12300
rect 18288 12288 18294 12300
rect 19812 12288 19840 12319
rect 18288 12260 19840 12288
rect 18288 12248 18294 12260
rect 20910 12223 20968 12229
rect 20910 12220 20922 12223
rect 17092 12192 17128 12220
rect 18156 12192 20922 12220
rect 17034 12180 17040 12183
rect 17092 12180 17098 12192
rect 20910 12189 20922 12192
rect 20956 12189 20968 12223
rect 20910 12183 20968 12189
rect 21177 12223 21235 12229
rect 21177 12189 21189 12223
rect 21223 12220 21235 12223
rect 21266 12220 21272 12232
rect 21223 12192 21272 12220
rect 21223 12189 21235 12192
rect 21177 12183 21235 12189
rect 10836 12124 11376 12152
rect 10836 12112 10842 12124
rect 11698 12112 11704 12164
rect 11756 12152 11762 12164
rect 12066 12152 12072 12164
rect 11756 12124 12072 12152
rect 11756 12112 11762 12124
rect 12066 12112 12072 12124
rect 12124 12112 12130 12164
rect 12796 12155 12854 12161
rect 12796 12121 12808 12155
rect 12842 12152 12854 12155
rect 12986 12152 12992 12164
rect 12842 12124 12992 12152
rect 12842 12121 12854 12124
rect 12796 12115 12854 12121
rect 12986 12112 12992 12124
rect 13044 12112 13050 12164
rect 15286 12152 15292 12164
rect 13924 12124 15292 12152
rect 7837 12087 7895 12093
rect 7837 12084 7849 12087
rect 6656 12056 7849 12084
rect 7837 12053 7849 12056
rect 7883 12053 7895 12087
rect 7837 12047 7895 12053
rect 9122 12044 9128 12096
rect 9180 12084 9186 12096
rect 9309 12087 9367 12093
rect 9309 12084 9321 12087
rect 9180 12056 9321 12084
rect 9180 12044 9186 12056
rect 9309 12053 9321 12056
rect 9355 12053 9367 12087
rect 9309 12047 9367 12053
rect 9401 12087 9459 12093
rect 9401 12053 9413 12087
rect 9447 12084 9459 12087
rect 10042 12084 10048 12096
rect 9447 12056 10048 12084
rect 9447 12053 9459 12056
rect 9401 12047 9459 12053
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 10594 12084 10600 12096
rect 10507 12056 10600 12084
rect 10594 12044 10600 12056
rect 10652 12084 10658 12096
rect 10962 12084 10968 12096
rect 10652 12056 10968 12084
rect 10652 12044 10658 12056
rect 10962 12044 10968 12056
rect 11020 12044 11026 12096
rect 11057 12087 11115 12093
rect 11057 12053 11069 12087
rect 11103 12084 11115 12087
rect 11146 12084 11152 12096
rect 11103 12056 11152 12084
rect 11103 12053 11115 12056
rect 11057 12047 11115 12053
rect 11146 12044 11152 12056
rect 11204 12084 11210 12096
rect 13446 12084 13452 12096
rect 11204 12056 13452 12084
rect 11204 12044 11210 12056
rect 13446 12044 13452 12056
rect 13504 12044 13510 12096
rect 13538 12044 13544 12096
rect 13596 12084 13602 12096
rect 13924 12093 13952 12124
rect 15286 12112 15292 12124
rect 15344 12112 15350 12164
rect 16424 12155 16482 12161
rect 16424 12121 16436 12155
rect 16470 12152 16482 12155
rect 19518 12152 19524 12164
rect 16470 12124 19524 12152
rect 16470 12121 16482 12124
rect 16424 12115 16482 12121
rect 19518 12112 19524 12124
rect 19576 12112 19582 12164
rect 20254 12152 20260 12164
rect 19720 12124 20260 12152
rect 13909 12087 13967 12093
rect 13909 12084 13921 12087
rect 13596 12056 13921 12084
rect 13596 12044 13602 12056
rect 13909 12053 13921 12056
rect 13955 12053 13967 12087
rect 14182 12084 14188 12096
rect 14143 12056 14188 12084
rect 13909 12047 13967 12053
rect 14182 12044 14188 12056
rect 14240 12084 14246 12096
rect 14369 12087 14427 12093
rect 14369 12084 14381 12087
rect 14240 12056 14381 12084
rect 14240 12044 14246 12056
rect 14369 12053 14381 12056
rect 14415 12053 14427 12087
rect 14369 12047 14427 12053
rect 15010 12044 15016 12096
rect 15068 12084 15074 12096
rect 19720 12084 19748 12124
rect 20254 12112 20260 12124
rect 20312 12112 20318 12164
rect 15068 12056 19748 12084
rect 15068 12044 15074 12056
rect 20990 12044 20996 12096
rect 21048 12084 21054 12096
rect 21192 12084 21220 12183
rect 21266 12180 21272 12192
rect 21324 12180 21330 12232
rect 21269 12087 21327 12093
rect 21269 12084 21281 12087
rect 21048 12056 21281 12084
rect 21048 12044 21054 12056
rect 21269 12053 21281 12056
rect 21315 12053 21327 12087
rect 21269 12047 21327 12053
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3973 11883 4031 11889
rect 3973 11880 3985 11883
rect 3016 11852 3985 11880
rect 3016 11840 3022 11852
rect 3973 11849 3985 11852
rect 4019 11849 4031 11883
rect 3973 11843 4031 11849
rect 6365 11883 6423 11889
rect 6365 11849 6377 11883
rect 6411 11880 6423 11883
rect 6546 11880 6552 11892
rect 6411 11852 6552 11880
rect 6411 11849 6423 11852
rect 6365 11843 6423 11849
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 7282 11880 7288 11892
rect 7243 11852 7288 11880
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 8389 11883 8447 11889
rect 8389 11849 8401 11883
rect 8435 11880 8447 11883
rect 9674 11880 9680 11892
rect 8435 11852 9680 11880
rect 8435 11849 8447 11852
rect 8389 11843 8447 11849
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 9769 11883 9827 11889
rect 9769 11849 9781 11883
rect 9815 11880 9827 11883
rect 10137 11883 10195 11889
rect 10137 11880 10149 11883
rect 9815 11852 10149 11880
rect 9815 11849 9827 11852
rect 9769 11843 9827 11849
rect 10137 11849 10149 11852
rect 10183 11849 10195 11883
rect 10137 11843 10195 11849
rect 10318 11840 10324 11892
rect 10376 11880 10382 11892
rect 10505 11883 10563 11889
rect 10505 11880 10517 11883
rect 10376 11852 10517 11880
rect 10376 11840 10382 11852
rect 10505 11849 10517 11852
rect 10551 11849 10563 11883
rect 10505 11843 10563 11849
rect 11238 11840 11244 11892
rect 11296 11880 11302 11892
rect 11517 11883 11575 11889
rect 11517 11880 11529 11883
rect 11296 11852 11529 11880
rect 11296 11840 11302 11852
rect 11517 11849 11529 11852
rect 11563 11849 11575 11883
rect 11517 11843 11575 11849
rect 12342 11840 12348 11892
rect 12400 11880 12406 11892
rect 12529 11883 12587 11889
rect 12529 11880 12541 11883
rect 12400 11852 12541 11880
rect 12400 11840 12406 11852
rect 12529 11849 12541 11852
rect 12575 11849 12587 11883
rect 12529 11843 12587 11849
rect 16298 11840 16304 11892
rect 16356 11840 16362 11892
rect 5442 11772 5448 11824
rect 5500 11812 5506 11824
rect 5537 11815 5595 11821
rect 5537 11812 5549 11815
rect 5500 11784 5549 11812
rect 5500 11772 5506 11784
rect 5537 11781 5549 11784
rect 5583 11812 5595 11815
rect 6914 11812 6920 11824
rect 5583 11784 6920 11812
rect 5583 11781 5595 11784
rect 5537 11775 5595 11781
rect 6914 11772 6920 11784
rect 6972 11772 6978 11824
rect 7926 11772 7932 11824
rect 7984 11772 7990 11824
rect 8110 11772 8116 11824
rect 8168 11812 8174 11824
rect 10778 11812 10784 11824
rect 8168 11784 10784 11812
rect 8168 11772 8174 11784
rect 10778 11772 10784 11784
rect 10836 11772 10842 11824
rect 16316 11812 16344 11840
rect 20809 11815 20867 11821
rect 20809 11812 20821 11815
rect 13556 11784 16344 11812
rect 19352 11784 20821 11812
rect 1394 11744 1400 11756
rect 1355 11716 1400 11744
rect 1394 11704 1400 11716
rect 1452 11704 1458 11756
rect 1670 11744 1676 11756
rect 1631 11716 1676 11744
rect 1670 11704 1676 11716
rect 1728 11744 1734 11756
rect 1949 11747 2007 11753
rect 1949 11744 1961 11747
rect 1728 11716 1961 11744
rect 1728 11704 1734 11716
rect 1949 11713 1961 11716
rect 1995 11713 2007 11747
rect 4154 11744 4160 11756
rect 4115 11716 4160 11744
rect 1949 11707 2007 11713
rect 4154 11704 4160 11716
rect 4212 11704 4218 11756
rect 6086 11704 6092 11756
rect 6144 11744 6150 11756
rect 6733 11747 6791 11753
rect 6733 11744 6745 11747
rect 6144 11716 6745 11744
rect 6144 11704 6150 11716
rect 6733 11713 6745 11716
rect 6779 11713 6791 11747
rect 7944 11744 7972 11772
rect 6733 11707 6791 11713
rect 7760 11716 7972 11744
rect 8021 11747 8079 11753
rect 1412 11676 1440 11704
rect 2133 11679 2191 11685
rect 2133 11676 2145 11679
rect 1412 11648 2145 11676
rect 2133 11645 2145 11648
rect 2179 11645 2191 11679
rect 2133 11639 2191 11645
rect 4982 11636 4988 11688
rect 5040 11676 5046 11688
rect 5077 11679 5135 11685
rect 5077 11676 5089 11679
rect 5040 11648 5089 11676
rect 5040 11636 5046 11648
rect 5077 11645 5089 11648
rect 5123 11645 5135 11679
rect 5077 11639 5135 11645
rect 6825 11679 6883 11685
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 7009 11679 7067 11685
rect 6871 11648 6960 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 1857 11543 1915 11549
rect 1857 11509 1869 11543
rect 1903 11540 1915 11543
rect 4522 11540 4528 11552
rect 1903 11512 4528 11540
rect 1903 11509 1915 11512
rect 1857 11503 1915 11509
rect 4522 11500 4528 11512
rect 4580 11500 4586 11552
rect 5997 11543 6055 11549
rect 5997 11509 6009 11543
rect 6043 11540 6055 11543
rect 6086 11540 6092 11552
rect 6043 11512 6092 11540
rect 6043 11509 6055 11512
rect 5997 11503 6055 11509
rect 6086 11500 6092 11512
rect 6144 11500 6150 11552
rect 6181 11543 6239 11549
rect 6181 11509 6193 11543
rect 6227 11540 6239 11543
rect 6932 11540 6960 11648
rect 7009 11645 7021 11679
rect 7055 11676 7067 11679
rect 7282 11676 7288 11688
rect 7055 11648 7288 11676
rect 7055 11645 7067 11648
rect 7009 11639 7067 11645
rect 7282 11636 7288 11648
rect 7340 11636 7346 11688
rect 7760 11685 7788 11716
rect 8021 11713 8033 11747
rect 8067 11744 8079 11747
rect 8662 11744 8668 11756
rect 8067 11716 8668 11744
rect 8067 11713 8079 11716
rect 8021 11707 8079 11713
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 9214 11704 9220 11756
rect 9272 11744 9278 11756
rect 9490 11744 9496 11756
rect 9272 11716 9496 11744
rect 9272 11704 9278 11716
rect 9490 11704 9496 11716
rect 9548 11704 9554 11756
rect 9674 11744 9680 11756
rect 9635 11716 9680 11744
rect 9674 11704 9680 11716
rect 9732 11704 9738 11756
rect 10597 11747 10655 11753
rect 10597 11713 10609 11747
rect 10643 11744 10655 11747
rect 11698 11744 11704 11756
rect 10643 11716 11704 11744
rect 10643 11713 10655 11716
rect 10597 11707 10655 11713
rect 11698 11704 11704 11716
rect 11756 11704 11762 11756
rect 11882 11744 11888 11756
rect 11843 11716 11888 11744
rect 11882 11704 11888 11716
rect 11940 11744 11946 11756
rect 12437 11747 12495 11753
rect 12437 11744 12449 11747
rect 11940 11716 12449 11744
rect 11940 11704 11946 11716
rect 12437 11713 12449 11716
rect 12483 11744 12495 11747
rect 13556 11744 13584 11784
rect 12483 11716 13584 11744
rect 12483 11713 12495 11716
rect 12437 11707 12495 11713
rect 13630 11704 13636 11756
rect 13688 11753 13694 11756
rect 13688 11744 13700 11753
rect 16229 11747 16287 11753
rect 13688 11716 13733 11744
rect 13688 11707 13700 11716
rect 16229 11713 16241 11747
rect 16275 11744 16287 11747
rect 16390 11744 16396 11756
rect 16275 11716 16396 11744
rect 16275 11713 16287 11716
rect 16229 11707 16287 11713
rect 13688 11704 13694 11707
rect 16390 11704 16396 11716
rect 16448 11704 16454 11756
rect 16482 11704 16488 11756
rect 16540 11744 16546 11756
rect 16761 11747 16819 11753
rect 16761 11744 16773 11747
rect 16540 11716 16773 11744
rect 16540 11704 16546 11716
rect 16761 11713 16773 11716
rect 16807 11744 16819 11747
rect 16945 11747 17003 11753
rect 16945 11744 16957 11747
rect 16807 11716 16957 11744
rect 16807 11713 16819 11716
rect 16761 11707 16819 11713
rect 16945 11713 16957 11716
rect 16991 11744 17003 11747
rect 17129 11747 17187 11753
rect 17129 11744 17141 11747
rect 16991 11716 17141 11744
rect 16991 11713 17003 11716
rect 16945 11707 17003 11713
rect 17129 11713 17141 11716
rect 17175 11744 17187 11747
rect 17497 11747 17555 11753
rect 17497 11744 17509 11747
rect 17175 11716 17509 11744
rect 17175 11713 17187 11716
rect 17129 11707 17187 11713
rect 17497 11713 17509 11716
rect 17543 11713 17555 11747
rect 17753 11747 17811 11753
rect 17753 11744 17765 11747
rect 17497 11707 17555 11713
rect 17604 11716 17765 11744
rect 7745 11679 7803 11685
rect 7745 11645 7757 11679
rect 7791 11645 7803 11679
rect 7926 11676 7932 11688
rect 7887 11648 7932 11676
rect 7745 11639 7803 11645
rect 7926 11636 7932 11648
rect 7984 11636 7990 11688
rect 9950 11676 9956 11688
rect 9911 11648 9956 11676
rect 9950 11636 9956 11648
rect 10008 11636 10014 11688
rect 10778 11676 10784 11688
rect 10739 11648 10784 11676
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 10962 11636 10968 11688
rect 11020 11676 11026 11688
rect 11149 11679 11207 11685
rect 11149 11676 11161 11679
rect 11020 11648 11161 11676
rect 11020 11636 11026 11648
rect 11149 11645 11161 11648
rect 11195 11676 11207 11679
rect 11790 11676 11796 11688
rect 11195 11648 11796 11676
rect 11195 11645 11207 11648
rect 11149 11639 11207 11645
rect 11790 11636 11796 11648
rect 11848 11636 11854 11688
rect 11974 11676 11980 11688
rect 11935 11648 11980 11676
rect 11974 11636 11980 11648
rect 12032 11636 12038 11688
rect 12069 11679 12127 11685
rect 12069 11645 12081 11679
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 13909 11679 13967 11685
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 14182 11676 14188 11688
rect 13955 11648 14188 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 9306 11608 9312 11620
rect 9267 11580 9312 11608
rect 9306 11568 9312 11580
rect 9364 11568 9370 11620
rect 11054 11568 11060 11620
rect 11112 11608 11118 11620
rect 12084 11608 12112 11639
rect 12618 11608 12624 11620
rect 11112 11580 12624 11608
rect 11112 11568 11118 11580
rect 12618 11568 12624 11580
rect 12676 11568 12682 11620
rect 7098 11540 7104 11552
rect 6227 11512 7104 11540
rect 6227 11509 6239 11512
rect 6181 11503 6239 11509
rect 7098 11500 7104 11512
rect 7156 11540 7162 11552
rect 7834 11540 7840 11552
rect 7156 11512 7840 11540
rect 7156 11500 7162 11512
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 11146 11500 11152 11552
rect 11204 11540 11210 11552
rect 11333 11543 11391 11549
rect 11333 11540 11345 11543
rect 11204 11512 11345 11540
rect 11204 11500 11210 11512
rect 11333 11509 11345 11512
rect 11379 11540 11391 11543
rect 11698 11540 11704 11552
rect 11379 11512 11704 11540
rect 11379 11509 11391 11512
rect 11333 11503 11391 11509
rect 11698 11500 11704 11512
rect 11756 11500 11762 11552
rect 12526 11500 12532 11552
rect 12584 11540 12590 11552
rect 13262 11540 13268 11552
rect 12584 11512 13268 11540
rect 12584 11500 12590 11512
rect 13262 11500 13268 11512
rect 13320 11540 13326 11552
rect 13924 11540 13952 11639
rect 14182 11636 14188 11648
rect 14240 11636 14246 11688
rect 17604 11676 17632 11716
rect 17753 11713 17765 11716
rect 17799 11713 17811 11747
rect 17753 11707 17811 11713
rect 19352 11685 19380 11784
rect 20809 11781 20821 11784
rect 20855 11812 20867 11815
rect 20990 11812 20996 11824
rect 20855 11784 20996 11812
rect 20855 11781 20867 11784
rect 20809 11775 20867 11781
rect 20990 11772 20996 11784
rect 21048 11772 21054 11824
rect 19604 11747 19662 11753
rect 19604 11713 19616 11747
rect 19650 11744 19662 11747
rect 19886 11744 19892 11756
rect 19650 11716 19892 11744
rect 19650 11713 19662 11716
rect 19604 11707 19662 11713
rect 19886 11704 19892 11716
rect 19944 11704 19950 11756
rect 19337 11679 19395 11685
rect 19337 11676 19349 11679
rect 16500 11648 17632 11676
rect 18984 11648 19349 11676
rect 16500 11620 16528 11648
rect 16482 11568 16488 11620
rect 16540 11568 16546 11620
rect 18984 11617 19012 11648
rect 19337 11645 19349 11648
rect 19383 11645 19395 11679
rect 19337 11639 19395 11645
rect 18969 11611 19027 11617
rect 18969 11608 18981 11611
rect 18432 11580 18981 11608
rect 18432 11552 18460 11580
rect 18969 11577 18981 11580
rect 19015 11577 19027 11611
rect 18969 11571 19027 11577
rect 14001 11543 14059 11549
rect 14001 11540 14013 11543
rect 13320 11512 14013 11540
rect 13320 11500 13326 11512
rect 14001 11509 14013 11512
rect 14047 11509 14059 11543
rect 14001 11503 14059 11509
rect 15010 11500 15016 11552
rect 15068 11540 15074 11552
rect 15105 11543 15163 11549
rect 15105 11540 15117 11543
rect 15068 11512 15117 11540
rect 15068 11500 15074 11512
rect 15105 11509 15117 11512
rect 15151 11509 15163 11543
rect 15105 11503 15163 11509
rect 15470 11500 15476 11552
rect 15528 11540 15534 11552
rect 18230 11540 18236 11552
rect 15528 11512 18236 11540
rect 15528 11500 15534 11512
rect 18230 11500 18236 11512
rect 18288 11500 18294 11552
rect 18414 11500 18420 11552
rect 18472 11500 18478 11552
rect 18877 11543 18935 11549
rect 18877 11509 18889 11543
rect 18923 11540 18935 11543
rect 19610 11540 19616 11552
rect 18923 11512 19616 11540
rect 18923 11509 18935 11512
rect 18877 11503 18935 11509
rect 19610 11500 19616 11512
rect 19668 11500 19674 11552
rect 20717 11543 20775 11549
rect 20717 11509 20729 11543
rect 20763 11540 20775 11543
rect 20898 11540 20904 11552
rect 20763 11512 20904 11540
rect 20763 11509 20775 11512
rect 20717 11503 20775 11509
rect 20898 11500 20904 11512
rect 20956 11500 20962 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 1762 11296 1768 11348
rect 1820 11336 1826 11348
rect 1857 11339 1915 11345
rect 1857 11336 1869 11339
rect 1820 11308 1869 11336
rect 1820 11296 1826 11308
rect 1857 11305 1869 11308
rect 1903 11305 1915 11339
rect 2130 11336 2136 11348
rect 2091 11308 2136 11336
rect 1857 11299 1915 11305
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 5258 11336 5264 11348
rect 2746 11308 5264 11336
rect 1581 11271 1639 11277
rect 1581 11237 1593 11271
rect 1627 11268 1639 11271
rect 2746 11268 2774 11308
rect 5258 11296 5264 11308
rect 5316 11296 5322 11348
rect 5353 11339 5411 11345
rect 5353 11305 5365 11339
rect 5399 11336 5411 11339
rect 5718 11336 5724 11348
rect 5399 11308 5724 11336
rect 5399 11305 5411 11308
rect 5353 11299 5411 11305
rect 5718 11296 5724 11308
rect 5776 11296 5782 11348
rect 5994 11296 6000 11348
rect 6052 11336 6058 11348
rect 6181 11339 6239 11345
rect 6181 11336 6193 11339
rect 6052 11308 6193 11336
rect 6052 11296 6058 11308
rect 6181 11305 6193 11308
rect 6227 11305 6239 11339
rect 7006 11336 7012 11348
rect 6967 11308 7012 11336
rect 6181 11299 6239 11305
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 7282 11296 7288 11348
rect 7340 11336 7346 11348
rect 7377 11339 7435 11345
rect 7377 11336 7389 11339
rect 7340 11308 7389 11336
rect 7340 11296 7346 11308
rect 7377 11305 7389 11308
rect 7423 11305 7435 11339
rect 12802 11336 12808 11348
rect 7377 11299 7435 11305
rect 9600 11308 12808 11336
rect 1627 11240 2774 11268
rect 1627 11237 1639 11240
rect 1581 11231 1639 11237
rect 4154 11228 4160 11280
rect 4212 11268 4218 11280
rect 8941 11271 8999 11277
rect 8941 11268 8953 11271
rect 4212 11240 8953 11268
rect 4212 11228 4218 11240
rect 8941 11237 8953 11240
rect 8987 11237 8999 11271
rect 8941 11231 8999 11237
rect 4801 11203 4859 11209
rect 4801 11169 4813 11203
rect 4847 11200 4859 11203
rect 5442 11200 5448 11212
rect 4847 11172 5448 11200
rect 4847 11169 4859 11172
rect 4801 11163 4859 11169
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 5629 11203 5687 11209
rect 5629 11169 5641 11203
rect 5675 11169 5687 11203
rect 5629 11163 5687 11169
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11132 1458 11144
rect 1673 11135 1731 11141
rect 1673 11132 1685 11135
rect 1452 11104 1685 11132
rect 1452 11092 1458 11104
rect 1673 11101 1685 11104
rect 1719 11101 1731 11135
rect 1673 11095 1731 11101
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11101 2099 11135
rect 2041 11095 2099 11101
rect 2317 11135 2375 11141
rect 2317 11101 2329 11135
rect 2363 11132 2375 11135
rect 3878 11132 3884 11144
rect 2363 11104 3884 11132
rect 2363 11101 2375 11104
rect 2317 11095 2375 11101
rect 2056 11064 2084 11095
rect 3878 11092 3884 11104
rect 3936 11092 3942 11144
rect 4982 11132 4988 11144
rect 4943 11104 4988 11132
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 5644 11132 5672 11163
rect 5902 11160 5908 11212
rect 5960 11200 5966 11212
rect 6365 11203 6423 11209
rect 6365 11200 6377 11203
rect 5960 11172 6377 11200
rect 5960 11160 5966 11172
rect 6365 11169 6377 11172
rect 6411 11169 6423 11203
rect 6914 11200 6920 11212
rect 6365 11163 6423 11169
rect 6472 11172 6920 11200
rect 6472 11132 6500 11172
rect 6914 11160 6920 11172
rect 6972 11200 6978 11212
rect 7282 11200 7288 11212
rect 6972 11172 7288 11200
rect 6972 11160 6978 11172
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 9600 11209 9628 11308
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 15930 11336 15936 11348
rect 13004 11308 15936 11336
rect 10042 11268 10048 11280
rect 10003 11240 10048 11268
rect 10042 11228 10048 11240
rect 10100 11228 10106 11280
rect 10318 11228 10324 11280
rect 10376 11268 10382 11280
rect 10965 11271 11023 11277
rect 10965 11268 10977 11271
rect 10376 11240 10977 11268
rect 10376 11228 10382 11240
rect 10965 11237 10977 11240
rect 11011 11237 11023 11271
rect 10965 11231 11023 11237
rect 11241 11271 11299 11277
rect 11241 11237 11253 11271
rect 11287 11268 11299 11271
rect 11514 11268 11520 11280
rect 11287 11240 11520 11268
rect 11287 11237 11299 11240
rect 11241 11231 11299 11237
rect 9585 11203 9643 11209
rect 9585 11169 9597 11203
rect 9631 11169 9643 11203
rect 9950 11200 9956 11212
rect 9911 11172 9956 11200
rect 9585 11163 9643 11169
rect 9950 11160 9956 11172
rect 10008 11200 10014 11212
rect 10505 11203 10563 11209
rect 10505 11200 10517 11203
rect 10008 11172 10517 11200
rect 10008 11160 10014 11172
rect 10505 11169 10517 11172
rect 10551 11169 10563 11203
rect 10505 11163 10563 11169
rect 10410 11132 10416 11144
rect 5644 11104 6500 11132
rect 10371 11104 10416 11132
rect 10410 11092 10416 11104
rect 10468 11092 10474 11144
rect 3050 11064 3056 11076
rect 2056 11036 3056 11064
rect 3050 11024 3056 11036
rect 3108 11024 3114 11076
rect 4246 11024 4252 11076
rect 4304 11064 4310 11076
rect 4433 11067 4491 11073
rect 4433 11064 4445 11067
rect 4304 11036 4445 11064
rect 4304 11024 4310 11036
rect 4433 11033 4445 11036
rect 4479 11064 4491 11067
rect 4479 11036 4568 11064
rect 4479 11033 4491 11036
rect 4433 11027 4491 11033
rect 4540 10996 4568 11036
rect 4614 11024 4620 11076
rect 4672 11064 4678 11076
rect 4890 11064 4896 11076
rect 4672 11036 4896 11064
rect 4672 11024 4678 11036
rect 4890 11024 4896 11036
rect 4948 11024 4954 11076
rect 5626 11064 5632 11076
rect 5000 11036 5632 11064
rect 5000 10996 5028 11036
rect 5626 11024 5632 11036
rect 5684 11064 5690 11076
rect 5721 11067 5779 11073
rect 5721 11064 5733 11067
rect 5684 11036 5733 11064
rect 5684 11024 5690 11036
rect 5721 11033 5733 11036
rect 5767 11033 5779 11067
rect 5721 11027 5779 11033
rect 5813 11067 5871 11073
rect 5813 11033 5825 11067
rect 5859 11064 5871 11067
rect 7101 11067 7159 11073
rect 7101 11064 7113 11067
rect 5859 11036 7113 11064
rect 5859 11033 5871 11036
rect 5813 11027 5871 11033
rect 7101 11033 7113 11036
rect 7147 11033 7159 11067
rect 9306 11064 9312 11076
rect 9267 11036 9312 11064
rect 7101 11027 7159 11033
rect 9306 11024 9312 11036
rect 9364 11024 9370 11076
rect 10520 11064 10548 11163
rect 10594 11160 10600 11212
rect 10652 11200 10658 11212
rect 10870 11200 10876 11212
rect 10652 11172 10876 11200
rect 10652 11160 10658 11172
rect 10870 11160 10876 11172
rect 10928 11160 10934 11212
rect 10980 11200 11008 11231
rect 11514 11228 11520 11240
rect 11572 11228 11578 11280
rect 12618 11228 12624 11280
rect 12676 11268 12682 11280
rect 13004 11277 13032 11308
rect 15930 11296 15936 11308
rect 15988 11296 15994 11348
rect 16114 11296 16120 11348
rect 16172 11336 16178 11348
rect 16482 11336 16488 11348
rect 16172 11308 16488 11336
rect 16172 11296 16178 11308
rect 16482 11296 16488 11308
rect 16540 11336 16546 11348
rect 16577 11339 16635 11345
rect 16577 11336 16589 11339
rect 16540 11308 16589 11336
rect 16540 11296 16546 11308
rect 16577 11305 16589 11308
rect 16623 11305 16635 11339
rect 19613 11339 19671 11345
rect 19613 11336 19625 11339
rect 16577 11299 16635 11305
rect 17052 11308 19625 11336
rect 12989 11271 13047 11277
rect 12989 11268 13001 11271
rect 12676 11240 13001 11268
rect 12676 11228 12682 11240
rect 12989 11237 13001 11240
rect 13035 11237 13047 11271
rect 12989 11231 13047 11237
rect 16669 11271 16727 11277
rect 16669 11237 16681 11271
rect 16715 11268 16727 11271
rect 16942 11268 16948 11280
rect 16715 11240 16948 11268
rect 16715 11237 16727 11240
rect 16669 11231 16727 11237
rect 16942 11228 16948 11240
rect 17000 11228 17006 11280
rect 10980 11172 11652 11200
rect 11238 11092 11244 11144
rect 11296 11132 11302 11144
rect 11517 11135 11575 11141
rect 11517 11132 11529 11135
rect 11296 11104 11529 11132
rect 11296 11092 11302 11104
rect 11517 11101 11529 11104
rect 11563 11101 11575 11135
rect 11624 11132 11652 11172
rect 14274 11160 14280 11212
rect 14332 11200 14338 11212
rect 15194 11200 15200 11212
rect 14332 11172 15200 11200
rect 14332 11160 14338 11172
rect 15194 11160 15200 11172
rect 15252 11160 15258 11212
rect 16390 11160 16396 11212
rect 16448 11200 16454 11212
rect 17052 11200 17080 11308
rect 19613 11305 19625 11308
rect 19659 11305 19671 11339
rect 19613 11299 19671 11305
rect 18325 11203 18383 11209
rect 18325 11200 18337 11203
rect 16448 11172 17080 11200
rect 17972 11172 18337 11200
rect 16448 11160 16454 11172
rect 12250 11132 12256 11144
rect 11624 11104 12256 11132
rect 11517 11095 11575 11101
rect 12250 11092 12256 11104
rect 12308 11092 12314 11144
rect 15286 11092 15292 11144
rect 15344 11132 15350 11144
rect 16408 11132 16436 11160
rect 15344 11104 16436 11132
rect 15344 11092 15350 11104
rect 17972 11076 18000 11172
rect 18325 11169 18337 11172
rect 18371 11169 18383 11203
rect 20990 11200 20996 11212
rect 20951 11172 20996 11200
rect 18325 11163 18383 11169
rect 20990 11160 20996 11172
rect 21048 11200 21054 11212
rect 21085 11203 21143 11209
rect 21085 11200 21097 11203
rect 21048 11172 21097 11200
rect 21048 11160 21054 11172
rect 21085 11169 21097 11172
rect 21131 11169 21143 11203
rect 21085 11163 21143 11169
rect 18049 11135 18107 11141
rect 18049 11101 18061 11135
rect 18095 11132 18107 11135
rect 18095 11104 18184 11132
rect 18095 11101 18107 11104
rect 18049 11095 18107 11101
rect 11422 11064 11428 11076
rect 10520 11036 11284 11064
rect 11383 11036 11428 11064
rect 6546 10996 6552 11008
rect 4540 10968 5028 10996
rect 6507 10968 6552 10996
rect 6546 10956 6552 10968
rect 6604 10956 6610 11008
rect 6638 10956 6644 11008
rect 6696 10996 6702 11008
rect 8573 10999 8631 11005
rect 6696 10968 6741 10996
rect 6696 10956 6702 10968
rect 8573 10965 8585 10999
rect 8619 10996 8631 10999
rect 8754 10996 8760 11008
rect 8619 10968 8760 10996
rect 8619 10965 8631 10968
rect 8573 10959 8631 10965
rect 8754 10956 8760 10968
rect 8812 10956 8818 11008
rect 9398 10956 9404 11008
rect 9456 10996 9462 11008
rect 11256 10996 11284 11036
rect 11422 11024 11428 11036
rect 11480 11024 11486 11076
rect 11606 11024 11612 11076
rect 11664 11064 11670 11076
rect 11784 11067 11842 11073
rect 11784 11064 11796 11067
rect 11664 11036 11796 11064
rect 11664 11024 11670 11036
rect 11784 11033 11796 11036
rect 11830 11033 11842 11067
rect 11784 11027 11842 11033
rect 12158 11024 12164 11076
rect 12216 11064 12222 11076
rect 15464 11067 15522 11073
rect 12216 11036 12940 11064
rect 12216 11024 12222 11036
rect 12526 10996 12532 11008
rect 9456 10968 9501 10996
rect 11256 10968 12532 10996
rect 9456 10956 9462 10968
rect 12526 10956 12532 10968
rect 12584 10956 12590 11008
rect 12912 11005 12940 11036
rect 15464 11033 15476 11067
rect 15510 11064 15522 11067
rect 15562 11064 15568 11076
rect 15510 11036 15568 11064
rect 15510 11033 15522 11036
rect 15464 11027 15522 11033
rect 15562 11024 15568 11036
rect 15620 11024 15626 11076
rect 17804 11067 17862 11073
rect 17804 11033 17816 11067
rect 17850 11064 17862 11067
rect 17954 11064 17960 11076
rect 17850 11036 17960 11064
rect 17850 11033 17862 11036
rect 17804 11027 17862 11033
rect 17954 11024 17960 11036
rect 18012 11024 18018 11076
rect 12897 10999 12955 11005
rect 12897 10965 12909 10999
rect 12943 10965 12955 10999
rect 13262 10996 13268 11008
rect 13223 10968 13268 10996
rect 12897 10959 12955 10965
rect 13262 10956 13268 10968
rect 13320 10956 13326 11008
rect 13354 10956 13360 11008
rect 13412 10996 13418 11008
rect 13449 10999 13507 11005
rect 13449 10996 13461 10999
rect 13412 10968 13461 10996
rect 13412 10956 13418 10968
rect 13449 10965 13461 10968
rect 13495 10996 13507 10999
rect 14642 10996 14648 11008
rect 13495 10968 14648 10996
rect 13495 10965 13507 10968
rect 13449 10959 13507 10965
rect 14642 10956 14648 10968
rect 14700 10956 14706 11008
rect 18156 11005 18184 11104
rect 19794 11024 19800 11076
rect 19852 11064 19858 11076
rect 20726 11067 20784 11073
rect 20726 11064 20738 11067
rect 19852 11036 20738 11064
rect 19852 11024 19858 11036
rect 20726 11033 20738 11036
rect 20772 11033 20784 11067
rect 20726 11027 20784 11033
rect 18141 10999 18199 11005
rect 18141 10965 18153 10999
rect 18187 10996 18199 10999
rect 18414 10996 18420 11008
rect 18187 10968 18420 10996
rect 18187 10965 18199 10968
rect 18141 10959 18199 10965
rect 18414 10956 18420 10968
rect 18472 10996 18478 11008
rect 18601 10999 18659 11005
rect 18601 10996 18613 10999
rect 18472 10968 18613 10996
rect 18472 10956 18478 10968
rect 18601 10965 18613 10968
rect 18647 10965 18659 10999
rect 18601 10959 18659 10965
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 5077 10795 5135 10801
rect 5077 10761 5089 10795
rect 5123 10792 5135 10795
rect 5166 10792 5172 10804
rect 5123 10764 5172 10792
rect 5123 10761 5135 10764
rect 5077 10755 5135 10761
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 5258 10752 5264 10804
rect 5316 10792 5322 10804
rect 5445 10795 5503 10801
rect 5445 10792 5457 10795
rect 5316 10764 5457 10792
rect 5316 10752 5322 10764
rect 5445 10761 5457 10764
rect 5491 10761 5503 10795
rect 5445 10755 5503 10761
rect 5905 10795 5963 10801
rect 5905 10761 5917 10795
rect 5951 10792 5963 10795
rect 6638 10792 6644 10804
rect 5951 10764 6644 10792
rect 5951 10761 5963 10764
rect 5905 10755 5963 10761
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 7926 10752 7932 10804
rect 7984 10792 7990 10804
rect 8205 10795 8263 10801
rect 8205 10792 8217 10795
rect 7984 10764 8217 10792
rect 7984 10752 7990 10764
rect 8205 10761 8217 10764
rect 8251 10761 8263 10795
rect 8205 10755 8263 10761
rect 8665 10795 8723 10801
rect 8665 10761 8677 10795
rect 8711 10792 8723 10795
rect 8754 10792 8760 10804
rect 8711 10764 8760 10792
rect 8711 10761 8723 10764
rect 8665 10755 8723 10761
rect 8754 10752 8760 10764
rect 8812 10752 8818 10804
rect 9030 10792 9036 10804
rect 8991 10764 9036 10792
rect 9030 10752 9036 10764
rect 9088 10752 9094 10804
rect 9125 10795 9183 10801
rect 9125 10761 9137 10795
rect 9171 10792 9183 10795
rect 9398 10792 9404 10804
rect 9171 10764 9404 10792
rect 9171 10761 9183 10764
rect 9125 10755 9183 10761
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 9490 10752 9496 10804
rect 9548 10792 9554 10804
rect 9548 10764 9593 10792
rect 9548 10752 9554 10764
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 10321 10795 10379 10801
rect 10321 10792 10333 10795
rect 9732 10764 10333 10792
rect 9732 10752 9738 10764
rect 10321 10761 10333 10764
rect 10367 10761 10379 10795
rect 10321 10755 10379 10761
rect 11698 10752 11704 10804
rect 11756 10792 11762 10804
rect 12434 10792 12440 10804
rect 11756 10764 12440 10792
rect 11756 10752 11762 10764
rect 12434 10752 12440 10764
rect 12492 10752 12498 10804
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 13354 10792 13360 10804
rect 12860 10764 13360 10792
rect 12860 10752 12866 10764
rect 13354 10752 13360 10764
rect 13412 10792 13418 10804
rect 13633 10795 13691 10801
rect 13633 10792 13645 10795
rect 13412 10764 13645 10792
rect 13412 10752 13418 10764
rect 13633 10761 13645 10764
rect 13679 10792 13691 10795
rect 19981 10795 20039 10801
rect 19981 10792 19993 10795
rect 13679 10764 19993 10792
rect 13679 10761 13691 10764
rect 13633 10755 13691 10761
rect 19981 10761 19993 10764
rect 20027 10761 20039 10795
rect 19981 10755 20039 10761
rect 3142 10684 3148 10736
rect 3200 10724 3206 10736
rect 6733 10727 6791 10733
rect 6733 10724 6745 10727
rect 3200 10696 6745 10724
rect 3200 10684 3206 10696
rect 6733 10693 6745 10696
rect 6779 10693 6791 10727
rect 7193 10727 7251 10733
rect 7193 10724 7205 10727
rect 6733 10687 6791 10693
rect 7024 10696 7205 10724
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10656 1458 10668
rect 1673 10659 1731 10665
rect 1673 10656 1685 10659
rect 1452 10628 1685 10656
rect 1452 10616 1458 10628
rect 1673 10625 1685 10628
rect 1719 10625 1731 10659
rect 1673 10619 1731 10625
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4430 10656 4436 10668
rect 4212 10628 4436 10656
rect 4212 10616 4218 10628
rect 4430 10616 4436 10628
rect 4488 10656 4494 10668
rect 4709 10659 4767 10665
rect 4709 10656 4721 10659
rect 4488 10628 4721 10656
rect 4488 10616 4494 10628
rect 4709 10625 4721 10628
rect 4755 10625 4767 10659
rect 4709 10619 4767 10625
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10656 5595 10659
rect 5997 10659 6055 10665
rect 5997 10656 6009 10659
rect 5583 10628 6009 10656
rect 5583 10625 5595 10628
rect 5537 10619 5595 10625
rect 5997 10625 6009 10628
rect 6043 10625 6055 10659
rect 7024 10656 7052 10696
rect 7193 10693 7205 10696
rect 7239 10693 7251 10727
rect 8570 10724 8576 10736
rect 8531 10696 8576 10724
rect 7193 10687 7251 10693
rect 8570 10684 8576 10696
rect 8628 10684 8634 10736
rect 10594 10724 10600 10736
rect 9508 10696 10600 10724
rect 5997 10619 6055 10625
rect 6288 10628 7052 10656
rect 1578 10548 1584 10600
rect 1636 10588 1642 10600
rect 2314 10588 2320 10600
rect 1636 10560 2320 10588
rect 1636 10548 1642 10560
rect 2314 10548 2320 10560
rect 2372 10588 2378 10600
rect 4062 10588 4068 10600
rect 2372 10560 4068 10588
rect 2372 10548 2378 10560
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 4525 10591 4583 10597
rect 4525 10557 4537 10591
rect 4571 10557 4583 10591
rect 4525 10551 4583 10557
rect 4617 10591 4675 10597
rect 4617 10557 4629 10591
rect 4663 10588 4675 10591
rect 4890 10588 4896 10600
rect 4663 10560 4896 10588
rect 4663 10557 4675 10560
rect 4617 10551 4675 10557
rect 4540 10520 4568 10551
rect 4890 10548 4896 10560
rect 4948 10548 4954 10600
rect 5353 10591 5411 10597
rect 5353 10557 5365 10591
rect 5399 10588 5411 10591
rect 5718 10588 5724 10600
rect 5399 10560 5724 10588
rect 5399 10557 5411 10560
rect 5353 10551 5411 10557
rect 5718 10548 5724 10560
rect 5776 10588 5782 10600
rect 6288 10588 6316 10628
rect 7098 10616 7104 10668
rect 7156 10656 7162 10668
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 7156 10628 7849 10656
rect 7156 10616 7162 10628
rect 7837 10625 7849 10628
rect 7883 10625 7895 10659
rect 9508 10656 9536 10696
rect 10594 10684 10600 10696
rect 10652 10684 10658 10736
rect 10781 10727 10839 10733
rect 10781 10693 10793 10727
rect 10827 10724 10839 10727
rect 10962 10724 10968 10736
rect 10827 10696 10968 10724
rect 10827 10693 10839 10696
rect 10781 10687 10839 10693
rect 10962 10684 10968 10696
rect 11020 10684 11026 10736
rect 11238 10684 11244 10736
rect 11296 10724 11302 10736
rect 11296 10696 12940 10724
rect 11296 10684 11302 10696
rect 7837 10619 7895 10625
rect 8496 10628 9536 10656
rect 9585 10659 9643 10665
rect 6454 10588 6460 10600
rect 5776 10560 6316 10588
rect 6415 10560 6460 10588
rect 5776 10548 5782 10560
rect 6454 10548 6460 10560
rect 6512 10548 6518 10600
rect 6641 10591 6699 10597
rect 6641 10588 6653 10591
rect 6564 10560 6653 10588
rect 4798 10520 4804 10532
rect 4540 10492 4804 10520
rect 4798 10480 4804 10492
rect 4856 10480 4862 10532
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 2958 10412 2964 10464
rect 3016 10452 3022 10464
rect 6564 10452 6592 10560
rect 6641 10557 6653 10560
rect 6687 10557 6699 10591
rect 6641 10551 6699 10557
rect 6822 10548 6828 10600
rect 6880 10588 6886 10600
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 6880 10560 7573 10588
rect 6880 10548 6886 10560
rect 7561 10557 7573 10560
rect 7607 10557 7619 10591
rect 7561 10551 7619 10557
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10588 7803 10591
rect 7926 10588 7932 10600
rect 7791 10560 7932 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 7926 10548 7932 10560
rect 7984 10548 7990 10600
rect 8496 10597 8524 10628
rect 9585 10625 9597 10659
rect 9631 10656 9643 10659
rect 9766 10656 9772 10668
rect 9631 10628 9772 10656
rect 9631 10625 9643 10628
rect 9585 10619 9643 10625
rect 9766 10616 9772 10628
rect 9824 10616 9830 10668
rect 10689 10659 10747 10665
rect 10689 10625 10701 10659
rect 10735 10656 10747 10659
rect 11149 10659 11207 10665
rect 11149 10656 11161 10659
rect 10735 10628 11161 10656
rect 10735 10625 10747 10628
rect 10689 10619 10747 10625
rect 11149 10625 11161 10628
rect 11195 10625 11207 10659
rect 11149 10619 11207 10625
rect 12641 10659 12699 10665
rect 12641 10625 12653 10659
rect 12687 10656 12699 10659
rect 12802 10656 12808 10668
rect 12687 10628 12808 10656
rect 12687 10625 12699 10628
rect 12641 10619 12699 10625
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 12912 10665 12940 10696
rect 15194 10684 15200 10736
rect 15252 10724 15258 10736
rect 15749 10727 15807 10733
rect 15749 10724 15761 10727
rect 15252 10696 15761 10724
rect 15252 10684 15258 10696
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 13173 10659 13231 10665
rect 13173 10625 13185 10659
rect 13219 10656 13231 10659
rect 15102 10656 15108 10668
rect 13219 10628 15108 10656
rect 13219 10625 13231 10628
rect 13173 10619 13231 10625
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10557 8539 10591
rect 8481 10551 8539 10557
rect 9490 10548 9496 10600
rect 9548 10588 9554 10600
rect 9677 10591 9735 10597
rect 9677 10588 9689 10591
rect 9548 10560 9689 10588
rect 9548 10548 9554 10560
rect 9677 10557 9689 10560
rect 9723 10557 9735 10591
rect 9950 10588 9956 10600
rect 9911 10560 9956 10588
rect 9677 10551 9735 10557
rect 9950 10548 9956 10560
rect 10008 10548 10014 10600
rect 10870 10548 10876 10600
rect 10928 10588 10934 10600
rect 12912 10588 12940 10619
rect 15102 10616 15108 10628
rect 15160 10616 15166 10668
rect 15378 10656 15384 10668
rect 15436 10665 15442 10668
rect 15672 10665 15700 10696
rect 15749 10693 15761 10696
rect 15795 10724 15807 10727
rect 15933 10727 15991 10733
rect 15933 10724 15945 10727
rect 15795 10696 15945 10724
rect 15795 10693 15807 10696
rect 15749 10687 15807 10693
rect 15933 10693 15945 10696
rect 15979 10724 15991 10727
rect 15979 10696 16712 10724
rect 15979 10693 15991 10696
rect 15933 10687 15991 10693
rect 16684 10665 16712 10696
rect 17494 10684 17500 10736
rect 17552 10724 17558 10736
rect 21094 10727 21152 10733
rect 21094 10724 21106 10727
rect 17552 10696 21106 10724
rect 17552 10684 17558 10696
rect 21094 10693 21106 10696
rect 21140 10693 21152 10727
rect 21094 10687 21152 10693
rect 15348 10628 15384 10656
rect 15378 10616 15384 10628
rect 15436 10619 15448 10665
rect 15657 10659 15715 10665
rect 15657 10625 15669 10659
rect 15703 10625 15715 10659
rect 15657 10619 15715 10625
rect 16669 10659 16727 10665
rect 16669 10625 16681 10659
rect 16715 10625 16727 10659
rect 16925 10659 16983 10665
rect 16925 10656 16937 10659
rect 16669 10619 16727 10625
rect 16776 10628 16937 10656
rect 15436 10616 15442 10619
rect 13262 10588 13268 10600
rect 10928 10560 10973 10588
rect 12912 10560 13268 10588
rect 10928 10548 10934 10560
rect 13262 10548 13268 10560
rect 13320 10588 13326 10600
rect 13357 10591 13415 10597
rect 13357 10588 13369 10591
rect 13320 10560 13369 10588
rect 13320 10548 13326 10560
rect 13357 10557 13369 10560
rect 13403 10557 13415 10591
rect 16776 10588 16804 10628
rect 16925 10625 16937 10628
rect 16971 10625 16983 10659
rect 16925 10619 16983 10625
rect 17862 10616 17868 10668
rect 17920 10656 17926 10668
rect 18673 10659 18731 10665
rect 18673 10656 18685 10659
rect 17920 10628 18685 10656
rect 17920 10616 17926 10628
rect 18673 10625 18685 10628
rect 18719 10625 18731 10659
rect 18673 10619 18731 10625
rect 18414 10588 18420 10600
rect 13357 10551 13415 10557
rect 15672 10560 16804 10588
rect 18375 10560 18420 10588
rect 7282 10480 7288 10532
rect 7340 10520 7346 10532
rect 11054 10520 11060 10532
rect 7340 10492 11060 10520
rect 7340 10480 7346 10492
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 12986 10520 12992 10532
rect 12947 10492 12992 10520
rect 12986 10480 12992 10492
rect 13044 10480 13050 10532
rect 13464 10492 14412 10520
rect 3016 10424 6592 10452
rect 7101 10455 7159 10461
rect 3016 10412 3022 10424
rect 7101 10421 7113 10455
rect 7147 10452 7159 10455
rect 9766 10452 9772 10464
rect 7147 10424 9772 10452
rect 7147 10421 7159 10424
rect 7101 10415 7159 10421
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 9858 10412 9864 10464
rect 9916 10452 9922 10464
rect 11517 10455 11575 10461
rect 11517 10452 11529 10455
rect 9916 10424 11529 10452
rect 9916 10412 9922 10424
rect 11517 10421 11529 10424
rect 11563 10452 11575 10455
rect 13078 10452 13084 10464
rect 11563 10424 13084 10452
rect 11563 10421 11575 10424
rect 11517 10415 11575 10421
rect 13078 10412 13084 10424
rect 13136 10452 13142 10464
rect 13464 10452 13492 10492
rect 13136 10424 13492 10452
rect 13136 10412 13142 10424
rect 13814 10412 13820 10464
rect 13872 10452 13878 10464
rect 14277 10455 14335 10461
rect 14277 10452 14289 10455
rect 13872 10424 14289 10452
rect 13872 10412 13878 10424
rect 14277 10421 14289 10424
rect 14323 10421 14335 10455
rect 14384 10452 14412 10492
rect 15672 10452 15700 10560
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 21358 10588 21364 10600
rect 21319 10560 21364 10588
rect 21358 10548 21364 10560
rect 21416 10588 21422 10600
rect 21453 10591 21511 10597
rect 21453 10588 21465 10591
rect 21416 10560 21465 10588
rect 21416 10548 21422 10560
rect 21453 10557 21465 10560
rect 21499 10557 21511 10591
rect 21453 10551 21511 10557
rect 18141 10523 18199 10529
rect 18141 10520 18153 10523
rect 17604 10492 18153 10520
rect 14384 10424 15700 10452
rect 14277 10415 14335 10421
rect 16482 10412 16488 10464
rect 16540 10452 16546 10464
rect 17604 10452 17632 10492
rect 18141 10489 18153 10492
rect 18187 10489 18199 10523
rect 19702 10520 19708 10532
rect 18141 10483 18199 10489
rect 19628 10492 19708 10520
rect 16540 10424 17632 10452
rect 16540 10412 16546 10424
rect 17770 10412 17776 10464
rect 17828 10452 17834 10464
rect 18049 10455 18107 10461
rect 18049 10452 18061 10455
rect 17828 10424 18061 10452
rect 17828 10412 17834 10424
rect 18049 10421 18061 10424
rect 18095 10421 18107 10455
rect 18156 10452 18184 10483
rect 19628 10452 19656 10492
rect 19702 10480 19708 10492
rect 19760 10480 19766 10532
rect 19794 10452 19800 10464
rect 18156 10424 19656 10452
rect 19755 10424 19800 10452
rect 18049 10415 18107 10421
rect 19794 10412 19800 10424
rect 19852 10412 19858 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 2038 10208 2044 10260
rect 2096 10248 2102 10260
rect 2133 10251 2191 10257
rect 2133 10248 2145 10251
rect 2096 10220 2145 10248
rect 2096 10208 2102 10220
rect 2133 10217 2145 10220
rect 2179 10217 2191 10251
rect 3142 10248 3148 10260
rect 3103 10220 3148 10248
rect 2133 10211 2191 10217
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 3329 10251 3387 10257
rect 3329 10217 3341 10251
rect 3375 10248 3387 10251
rect 3418 10248 3424 10260
rect 3375 10220 3424 10248
rect 3375 10217 3387 10220
rect 3329 10211 3387 10217
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 4338 10208 4344 10260
rect 4396 10248 4402 10260
rect 4801 10251 4859 10257
rect 4801 10248 4813 10251
rect 4396 10220 4813 10248
rect 4396 10208 4402 10220
rect 4801 10217 4813 10220
rect 4847 10217 4859 10251
rect 4801 10211 4859 10217
rect 5629 10251 5687 10257
rect 5629 10217 5641 10251
rect 5675 10248 5687 10251
rect 5810 10248 5816 10260
rect 5675 10220 5816 10248
rect 5675 10217 5687 10220
rect 5629 10211 5687 10217
rect 5810 10208 5816 10220
rect 5868 10208 5874 10260
rect 6822 10208 6828 10260
rect 6880 10248 6886 10260
rect 7190 10248 7196 10260
rect 6880 10220 7052 10248
rect 7151 10220 7196 10248
rect 6880 10208 6886 10220
rect 1581 10183 1639 10189
rect 1581 10149 1593 10183
rect 1627 10180 1639 10183
rect 4890 10180 4896 10192
rect 1627 10152 4896 10180
rect 1627 10149 1639 10152
rect 1581 10143 1639 10149
rect 4890 10140 4896 10152
rect 4948 10140 4954 10192
rect 6914 10180 6920 10192
rect 6288 10152 6920 10180
rect 2593 10115 2651 10121
rect 2593 10081 2605 10115
rect 2639 10112 2651 10115
rect 3326 10112 3332 10124
rect 2639 10084 3332 10112
rect 2639 10081 2651 10084
rect 2593 10075 2651 10081
rect 3326 10072 3332 10084
rect 3384 10072 3390 10124
rect 3786 10072 3792 10124
rect 3844 10112 3850 10124
rect 3881 10115 3939 10121
rect 3881 10112 3893 10115
rect 3844 10084 3893 10112
rect 3844 10072 3850 10084
rect 3881 10081 3893 10084
rect 3927 10081 3939 10115
rect 4062 10112 4068 10124
rect 4023 10084 4068 10112
rect 3881 10075 3939 10081
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 5537 10115 5595 10121
rect 4172 10084 5120 10112
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 1670 10044 1676 10056
rect 1631 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10044 1734 10056
rect 1949 10047 2007 10053
rect 1949 10044 1961 10047
rect 1728 10016 1961 10044
rect 1728 10004 1734 10016
rect 1949 10013 1961 10016
rect 1995 10013 2007 10047
rect 1949 10007 2007 10013
rect 2317 10047 2375 10053
rect 2317 10013 2329 10047
rect 2363 10044 2375 10047
rect 3418 10044 3424 10056
rect 2363 10016 3424 10044
rect 2363 10013 2375 10016
rect 2317 10007 2375 10013
rect 3418 10004 3424 10016
rect 3476 10004 3482 10056
rect 3970 10004 3976 10056
rect 4028 10044 4034 10056
rect 4172 10044 4200 10084
rect 4706 10044 4712 10056
rect 4028 10016 4200 10044
rect 4667 10016 4712 10044
rect 4028 10004 4034 10016
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 4982 10044 4988 10056
rect 4943 10016 4988 10044
rect 4982 10004 4988 10016
rect 5040 10004 5046 10056
rect 5092 10044 5120 10084
rect 5537 10081 5549 10115
rect 5583 10112 5595 10115
rect 5626 10112 5632 10124
rect 5583 10084 5632 10112
rect 5583 10081 5595 10084
rect 5537 10075 5595 10081
rect 5626 10072 5632 10084
rect 5684 10112 5690 10124
rect 6086 10112 6092 10124
rect 5684 10084 6092 10112
rect 5684 10072 5690 10084
rect 6086 10072 6092 10084
rect 6144 10072 6150 10124
rect 6288 10121 6316 10152
rect 6914 10140 6920 10152
rect 6972 10140 6978 10192
rect 7024 10180 7052 10220
rect 7190 10208 7196 10220
rect 7248 10208 7254 10260
rect 7285 10251 7343 10257
rect 7285 10217 7297 10251
rect 7331 10248 7343 10251
rect 7558 10248 7564 10260
rect 7331 10220 7564 10248
rect 7331 10217 7343 10220
rect 7285 10211 7343 10217
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 7926 10208 7932 10260
rect 7984 10248 7990 10260
rect 8297 10251 8355 10257
rect 8297 10248 8309 10251
rect 7984 10220 8309 10248
rect 7984 10208 7990 10220
rect 8297 10217 8309 10220
rect 8343 10217 8355 10251
rect 8297 10211 8355 10217
rect 8662 10208 8668 10260
rect 8720 10248 8726 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 8720 10220 8953 10248
rect 8720 10208 8726 10220
rect 8941 10217 8953 10220
rect 8987 10217 8999 10251
rect 8941 10211 8999 10217
rect 11701 10251 11759 10257
rect 11701 10217 11713 10251
rect 11747 10248 11759 10251
rect 14458 10248 14464 10260
rect 11747 10220 14464 10248
rect 11747 10217 11759 10220
rect 11701 10211 11759 10217
rect 14458 10208 14464 10220
rect 14516 10208 14522 10260
rect 7024 10152 9536 10180
rect 6273 10115 6331 10121
rect 6273 10081 6285 10115
rect 6319 10081 6331 10115
rect 6638 10112 6644 10124
rect 6599 10084 6644 10112
rect 6273 10075 6331 10081
rect 6638 10072 6644 10084
rect 6696 10072 6702 10124
rect 6822 10072 6828 10124
rect 6880 10072 6886 10124
rect 7006 10072 7012 10124
rect 7064 10112 7070 10124
rect 9508 10121 9536 10152
rect 7837 10115 7895 10121
rect 7837 10112 7849 10115
rect 7064 10084 7849 10112
rect 7064 10072 7070 10084
rect 7837 10081 7849 10084
rect 7883 10081 7895 10115
rect 7837 10075 7895 10081
rect 9493 10115 9551 10121
rect 9493 10081 9505 10115
rect 9539 10081 9551 10115
rect 9493 10075 9551 10081
rect 13081 10115 13139 10121
rect 13081 10081 13093 10115
rect 13127 10112 13139 10115
rect 13262 10112 13268 10124
rect 13127 10084 13268 10112
rect 13127 10081 13139 10084
rect 13081 10075 13139 10081
rect 13262 10072 13268 10084
rect 13320 10072 13326 10124
rect 13446 10072 13452 10124
rect 13504 10112 13510 10124
rect 13504 10084 14320 10112
rect 13504 10072 13510 10084
rect 6733 10047 6791 10053
rect 6733 10044 6745 10047
rect 5092 10016 6745 10044
rect 6733 10013 6745 10016
rect 6779 10013 6791 10047
rect 6840 10044 6868 10072
rect 7653 10047 7711 10053
rect 7653 10044 7665 10047
rect 6840 10016 7665 10044
rect 6733 10007 6791 10013
rect 7653 10013 7665 10016
rect 7699 10013 7711 10047
rect 7653 10007 7711 10013
rect 8018 10004 8024 10056
rect 8076 10044 8082 10056
rect 8205 10047 8263 10053
rect 8205 10044 8217 10047
rect 8076 10016 8217 10044
rect 8076 10004 8082 10016
rect 8205 10013 8217 10016
rect 8251 10044 8263 10047
rect 8570 10044 8576 10056
rect 8251 10016 8576 10044
rect 8251 10013 8263 10016
rect 8205 10007 8263 10013
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10044 9367 10047
rect 9950 10044 9956 10056
rect 9355 10016 9956 10044
rect 9355 10013 9367 10016
rect 9309 10007 9367 10013
rect 9950 10004 9956 10016
rect 10008 10004 10014 10056
rect 10137 10047 10195 10053
rect 10137 10013 10149 10047
rect 10183 10044 10195 10047
rect 11238 10044 11244 10056
rect 10183 10016 11244 10044
rect 10183 10013 10195 10016
rect 10137 10007 10195 10013
rect 11238 10004 11244 10016
rect 11296 10004 11302 10056
rect 13280 10044 13308 10072
rect 14185 10047 14243 10053
rect 14185 10044 14197 10047
rect 13280 10016 14197 10044
rect 14185 10013 14197 10016
rect 14231 10013 14243 10047
rect 14292 10044 14320 10084
rect 18708 10084 19380 10112
rect 14441 10047 14499 10053
rect 14441 10044 14453 10047
rect 14292 10016 14453 10044
rect 14185 10007 14243 10013
rect 14441 10013 14453 10016
rect 14487 10013 14499 10047
rect 17034 10044 17040 10056
rect 16995 10016 17040 10044
rect 14441 10007 14499 10013
rect 17034 10004 17040 10016
rect 17092 10044 17098 10056
rect 17129 10047 17187 10053
rect 17129 10044 17141 10047
rect 17092 10016 17141 10044
rect 17092 10004 17098 10016
rect 17129 10013 17141 10016
rect 17175 10013 17187 10047
rect 17129 10007 17187 10013
rect 17770 10004 17776 10056
rect 17828 10044 17834 10056
rect 18708 10044 18736 10084
rect 19245 10047 19303 10053
rect 19245 10044 19257 10047
rect 17828 10016 18736 10044
rect 18800 10016 19257 10044
rect 17828 10004 17834 10016
rect 3605 9979 3663 9985
rect 1872 9948 3556 9976
rect 1872 9917 1900 9948
rect 1857 9911 1915 9917
rect 1857 9877 1869 9911
rect 1903 9877 1915 9911
rect 2682 9908 2688 9920
rect 2643 9880 2688 9908
rect 1857 9871 1915 9877
rect 2682 9868 2688 9880
rect 2740 9868 2746 9920
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 3528 9908 3556 9948
rect 3605 9945 3617 9979
rect 3651 9976 3663 9979
rect 4157 9979 4215 9985
rect 4157 9976 4169 9979
rect 3651 9948 4169 9976
rect 3651 9945 3663 9948
rect 3605 9939 3663 9945
rect 4157 9945 4169 9948
rect 4203 9945 4215 9979
rect 6825 9979 6883 9985
rect 6825 9976 6837 9979
rect 4157 9939 4215 9945
rect 4540 9948 6837 9976
rect 4430 9908 4436 9920
rect 2832 9880 2877 9908
rect 3528 9880 4436 9908
rect 2832 9868 2838 9880
rect 4430 9868 4436 9880
rect 4488 9868 4494 9920
rect 4540 9917 4568 9948
rect 6825 9945 6837 9948
rect 6871 9945 6883 9979
rect 6825 9939 6883 9945
rect 6932 9948 9996 9976
rect 4525 9911 4583 9917
rect 4525 9877 4537 9911
rect 4571 9877 4583 9911
rect 4525 9871 4583 9877
rect 5902 9868 5908 9920
rect 5960 9908 5966 9920
rect 5997 9911 6055 9917
rect 5997 9908 6009 9911
rect 5960 9880 6009 9908
rect 5960 9868 5966 9880
rect 5997 9877 6009 9880
rect 6043 9877 6055 9911
rect 5997 9871 6055 9877
rect 6454 9868 6460 9920
rect 6512 9908 6518 9920
rect 6932 9908 6960 9948
rect 6512 9880 6960 9908
rect 7745 9911 7803 9917
rect 6512 9868 6518 9880
rect 7745 9877 7757 9911
rect 7791 9908 7803 9911
rect 8478 9908 8484 9920
rect 7791 9880 8484 9908
rect 7791 9877 7803 9880
rect 7745 9871 7803 9877
rect 8478 9868 8484 9880
rect 8536 9908 8542 9920
rect 8573 9911 8631 9917
rect 8573 9908 8585 9911
rect 8536 9880 8585 9908
rect 8536 9868 8542 9880
rect 8573 9877 8585 9880
rect 8619 9908 8631 9911
rect 9030 9908 9036 9920
rect 8619 9880 9036 9908
rect 8619 9877 8631 9880
rect 8573 9871 8631 9877
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 9398 9908 9404 9920
rect 9359 9880 9404 9908
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 9766 9908 9772 9920
rect 9727 9880 9772 9908
rect 9766 9868 9772 9880
rect 9824 9868 9830 9920
rect 9968 9908 9996 9948
rect 10042 9936 10048 9988
rect 10100 9976 10106 9988
rect 10382 9979 10440 9985
rect 10382 9976 10394 9979
rect 10100 9948 10394 9976
rect 10100 9936 10106 9948
rect 10382 9945 10394 9948
rect 10428 9945 10440 9979
rect 10382 9939 10440 9945
rect 12836 9979 12894 9985
rect 12836 9945 12848 9979
rect 12882 9976 12894 9979
rect 14274 9976 14280 9988
rect 12882 9948 14280 9976
rect 12882 9945 12894 9948
rect 12836 9939 12894 9945
rect 14274 9936 14280 9948
rect 14332 9936 14338 9988
rect 15930 9936 15936 9988
rect 15988 9976 15994 9988
rect 16482 9976 16488 9988
rect 15988 9948 16488 9976
rect 15988 9936 15994 9948
rect 16482 9936 16488 9948
rect 16540 9976 16546 9988
rect 16770 9979 16828 9985
rect 16770 9976 16782 9979
rect 16540 9948 16782 9976
rect 16540 9936 16546 9948
rect 16770 9945 16782 9948
rect 16816 9945 16828 9979
rect 17374 9979 17432 9985
rect 17374 9976 17386 9979
rect 16770 9939 16828 9945
rect 16868 9948 17386 9976
rect 10502 9908 10508 9920
rect 9968 9880 10508 9908
rect 10502 9868 10508 9880
rect 10560 9868 10566 9920
rect 10686 9868 10692 9920
rect 10744 9908 10750 9920
rect 11517 9911 11575 9917
rect 11517 9908 11529 9911
rect 10744 9880 11529 9908
rect 10744 9868 10750 9880
rect 11517 9877 11529 9880
rect 11563 9908 11575 9911
rect 13722 9908 13728 9920
rect 11563 9880 13728 9908
rect 11563 9877 11575 9880
rect 11517 9871 11575 9877
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 15562 9908 15568 9920
rect 15523 9880 15568 9908
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 15654 9868 15660 9920
rect 15712 9908 15718 9920
rect 15712 9880 15757 9908
rect 15712 9868 15718 9880
rect 16390 9868 16396 9920
rect 16448 9908 16454 9920
rect 16868 9908 16896 9948
rect 17374 9945 17386 9948
rect 17420 9945 17432 9979
rect 17374 9939 17432 9945
rect 18046 9936 18052 9988
rect 18104 9976 18110 9988
rect 18414 9976 18420 9988
rect 18104 9948 18420 9976
rect 18104 9936 18110 9948
rect 18414 9936 18420 9948
rect 18472 9976 18478 9988
rect 18800 9985 18828 10016
rect 19245 10013 19257 10016
rect 19291 10013 19303 10047
rect 19352 10044 19380 10084
rect 19501 10047 19559 10053
rect 19501 10044 19513 10047
rect 19352 10016 19513 10044
rect 19245 10007 19303 10013
rect 19501 10013 19513 10016
rect 19547 10013 19559 10047
rect 19501 10007 19559 10013
rect 18601 9979 18659 9985
rect 18601 9976 18613 9979
rect 18472 9948 18613 9976
rect 18472 9936 18478 9948
rect 18601 9945 18613 9948
rect 18647 9976 18659 9979
rect 18785 9979 18843 9985
rect 18785 9976 18797 9979
rect 18647 9948 18797 9976
rect 18647 9945 18659 9948
rect 18601 9939 18659 9945
rect 18785 9945 18797 9948
rect 18831 9945 18843 9979
rect 18785 9939 18843 9945
rect 18506 9908 18512 9920
rect 16448 9880 16896 9908
rect 18467 9880 18512 9908
rect 16448 9868 16454 9880
rect 18506 9868 18512 9880
rect 18564 9908 18570 9920
rect 19886 9908 19892 9920
rect 18564 9880 19892 9908
rect 18564 9868 18570 9880
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 20530 9868 20536 9920
rect 20588 9908 20594 9920
rect 20625 9911 20683 9917
rect 20625 9908 20637 9911
rect 20588 9880 20637 9908
rect 20588 9868 20594 9880
rect 20625 9877 20637 9880
rect 20671 9877 20683 9911
rect 20806 9908 20812 9920
rect 20767 9880 20812 9908
rect 20625 9871 20683 9877
rect 20806 9868 20812 9880
rect 20864 9908 20870 9920
rect 21358 9908 21364 9920
rect 20864 9880 21364 9908
rect 20864 9868 20870 9880
rect 21358 9868 21364 9880
rect 21416 9908 21422 9920
rect 21453 9911 21511 9917
rect 21453 9908 21465 9911
rect 21416 9880 21465 9908
rect 21416 9868 21422 9880
rect 21453 9877 21465 9880
rect 21499 9877 21511 9911
rect 21453 9871 21511 9877
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 1394 9704 1400 9716
rect 1355 9676 1400 9704
rect 1394 9664 1400 9676
rect 1452 9664 1458 9716
rect 2774 9664 2780 9716
rect 2832 9704 2838 9716
rect 2869 9707 2927 9713
rect 2869 9704 2881 9707
rect 2832 9676 2881 9704
rect 2832 9664 2838 9676
rect 2869 9673 2881 9676
rect 2915 9673 2927 9707
rect 2869 9667 2927 9673
rect 10410 9664 10416 9716
rect 10468 9704 10474 9716
rect 10468 9676 10824 9704
rect 10468 9664 10474 9676
rect 4430 9596 4436 9648
rect 4488 9636 4494 9648
rect 4893 9639 4951 9645
rect 4893 9636 4905 9639
rect 4488 9608 4905 9636
rect 4488 9596 4494 9608
rect 4893 9605 4905 9608
rect 4939 9605 4951 9639
rect 5442 9636 5448 9648
rect 5403 9608 5448 9636
rect 4893 9599 4951 9605
rect 5442 9596 5448 9608
rect 5500 9596 5506 9648
rect 5534 9596 5540 9648
rect 5592 9636 5598 9648
rect 5592 9608 5856 9636
rect 5592 9596 5598 9608
rect 1762 9568 1768 9580
rect 1723 9540 1768 9568
rect 1762 9528 1768 9540
rect 1820 9528 1826 9580
rect 2038 9568 2044 9580
rect 1999 9540 2044 9568
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 2130 9528 2136 9580
rect 2188 9568 2194 9580
rect 2317 9571 2375 9577
rect 2317 9568 2329 9571
rect 2188 9540 2329 9568
rect 2188 9528 2194 9540
rect 2317 9537 2329 9540
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9537 2651 9571
rect 5460 9568 5488 9596
rect 5828 9580 5856 9608
rect 6086 9596 6092 9648
rect 6144 9636 6150 9648
rect 6641 9639 6699 9645
rect 6641 9636 6653 9639
rect 6144 9608 6653 9636
rect 6144 9596 6150 9608
rect 6641 9605 6653 9608
rect 6687 9605 6699 9639
rect 6641 9599 6699 9605
rect 6914 9596 6920 9648
rect 6972 9636 6978 9648
rect 7193 9639 7251 9645
rect 7193 9636 7205 9639
rect 6972 9608 7205 9636
rect 6972 9596 6978 9608
rect 7193 9605 7205 9608
rect 7239 9605 7251 9639
rect 7193 9599 7251 9605
rect 9309 9639 9367 9645
rect 9309 9605 9321 9639
rect 9355 9636 9367 9639
rect 9766 9636 9772 9648
rect 9355 9608 9772 9636
rect 9355 9605 9367 9608
rect 9309 9599 9367 9605
rect 9766 9596 9772 9608
rect 9824 9596 9830 9648
rect 10796 9645 10824 9676
rect 12526 9664 12532 9716
rect 12584 9704 12590 9716
rect 13170 9704 13176 9716
rect 12584 9676 13176 9704
rect 12584 9664 12590 9676
rect 13170 9664 13176 9676
rect 13228 9664 13234 9716
rect 13814 9704 13820 9716
rect 13740 9676 13820 9704
rect 10781 9639 10839 9645
rect 10781 9605 10793 9639
rect 10827 9636 10839 9639
rect 10827 9608 10861 9636
rect 10827 9605 10839 9608
rect 10781 9599 10839 9605
rect 10962 9596 10968 9648
rect 11020 9636 11026 9648
rect 13480 9639 13538 9645
rect 13480 9636 13492 9639
rect 11020 9608 13492 9636
rect 11020 9596 11026 9608
rect 13480 9605 13492 9608
rect 13526 9636 13538 9639
rect 13740 9636 13768 9676
rect 13814 9664 13820 9676
rect 13872 9664 13878 9716
rect 20806 9664 20812 9716
rect 20864 9704 20870 9716
rect 21177 9707 21235 9713
rect 21177 9704 21189 9707
rect 20864 9676 21189 9704
rect 20864 9664 20870 9676
rect 13906 9636 13912 9648
rect 13526 9608 13768 9636
rect 13832 9608 13912 9636
rect 13526 9605 13538 9608
rect 13480 9599 13538 9605
rect 2593 9531 2651 9537
rect 4632 9540 5488 9568
rect 2222 9460 2228 9512
rect 2280 9500 2286 9512
rect 2608 9500 2636 9531
rect 4632 9509 4660 9540
rect 5810 9528 5816 9580
rect 5868 9528 5874 9580
rect 6733 9571 6791 9577
rect 6733 9568 6745 9571
rect 5920 9540 6745 9568
rect 2280 9472 2636 9500
rect 4617 9503 4675 9509
rect 2280 9460 2286 9472
rect 4617 9469 4629 9503
rect 4663 9469 4675 9503
rect 4798 9500 4804 9512
rect 4759 9472 4804 9500
rect 4617 9463 4675 9469
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 5350 9500 5356 9512
rect 5276 9472 5356 9500
rect 1486 9392 1492 9444
rect 1544 9432 1550 9444
rect 1581 9435 1639 9441
rect 1581 9432 1593 9435
rect 1544 9404 1593 9432
rect 1544 9392 1550 9404
rect 1581 9401 1593 9404
rect 1627 9401 1639 9435
rect 1854 9432 1860 9444
rect 1815 9404 1860 9432
rect 1581 9395 1639 9401
rect 1854 9392 1860 9404
rect 1912 9392 1918 9444
rect 1946 9392 1952 9444
rect 2004 9432 2010 9444
rect 2133 9435 2191 9441
rect 2133 9432 2145 9435
rect 2004 9404 2145 9432
rect 2004 9392 2010 9404
rect 2133 9401 2145 9404
rect 2179 9401 2191 9435
rect 2406 9432 2412 9444
rect 2367 9404 2412 9432
rect 2133 9395 2191 9401
rect 2406 9392 2412 9404
rect 2464 9392 2470 9444
rect 2498 9392 2504 9444
rect 2556 9432 2562 9444
rect 5166 9432 5172 9444
rect 2556 9404 5172 9432
rect 2556 9392 2562 9404
rect 5166 9392 5172 9404
rect 5224 9392 5230 9444
rect 5276 9441 5304 9472
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 5442 9460 5448 9512
rect 5500 9500 5506 9512
rect 5537 9503 5595 9509
rect 5537 9500 5549 9503
rect 5500 9472 5549 9500
rect 5500 9460 5506 9472
rect 5537 9469 5549 9472
rect 5583 9469 5595 9503
rect 5537 9463 5595 9469
rect 5261 9435 5319 9441
rect 5261 9401 5273 9435
rect 5307 9401 5319 9435
rect 5920 9432 5948 9540
rect 6733 9537 6745 9540
rect 6779 9537 6791 9571
rect 9490 9568 9496 9580
rect 6733 9531 6791 9537
rect 9140 9540 9496 9568
rect 9140 9509 9168 9540
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9537 10379 9571
rect 10321 9531 10379 9537
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9568 10471 9571
rect 11149 9571 11207 9577
rect 11149 9568 11161 9571
rect 10459 9540 11161 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 11149 9537 11161 9540
rect 11195 9568 11207 9571
rect 12526 9568 12532 9580
rect 11195 9540 12532 9568
rect 11195 9537 11207 9540
rect 11149 9531 11207 9537
rect 6457 9503 6515 9509
rect 6457 9469 6469 9503
rect 6503 9469 6515 9503
rect 6457 9463 6515 9469
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9469 9183 9503
rect 9125 9463 9183 9469
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9500 9275 9503
rect 9766 9500 9772 9512
rect 9263 9472 9772 9500
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 5261 9395 5319 9401
rect 5460 9404 5948 9432
rect 6472 9432 6500 9463
rect 7006 9432 7012 9444
rect 6472 9404 7012 9432
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 2832 9336 2877 9364
rect 2832 9324 2838 9336
rect 4522 9324 4528 9376
rect 4580 9364 4586 9376
rect 5460 9364 5488 9404
rect 7006 9392 7012 9404
rect 7064 9392 7070 9444
rect 7101 9435 7159 9441
rect 7101 9401 7113 9435
rect 7147 9432 7159 9435
rect 7650 9432 7656 9444
rect 7147 9404 7656 9432
rect 7147 9401 7159 9404
rect 7101 9395 7159 9401
rect 7650 9392 7656 9404
rect 7708 9392 7714 9444
rect 9232 9432 9260 9463
rect 9766 9460 9772 9472
rect 9824 9460 9830 9512
rect 10336 9500 10364 9531
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 13832 9568 13860 9608
rect 13906 9596 13912 9608
rect 13964 9596 13970 9648
rect 15654 9596 15660 9648
rect 15712 9636 15718 9648
rect 18386 9639 18444 9645
rect 18386 9636 18398 9639
rect 15712 9608 18398 9636
rect 15712 9596 15718 9608
rect 18386 9605 18398 9608
rect 18432 9605 18444 9639
rect 18386 9599 18444 9605
rect 14930 9571 14988 9577
rect 14930 9568 14942 9571
rect 12676 9540 13860 9568
rect 13924 9540 14942 9568
rect 12676 9528 12682 9540
rect 10597 9503 10655 9509
rect 10336 9472 10425 9500
rect 8772 9404 9260 9432
rect 4580 9336 5488 9364
rect 4580 9324 4586 9336
rect 5534 9324 5540 9376
rect 5592 9364 5598 9376
rect 6730 9364 6736 9376
rect 5592 9336 6736 9364
rect 5592 9324 5598 9336
rect 6730 9324 6736 9336
rect 6788 9324 6794 9376
rect 8478 9324 8484 9376
rect 8536 9364 8542 9376
rect 8772 9373 8800 9404
rect 9306 9392 9312 9444
rect 9364 9432 9370 9444
rect 9677 9435 9735 9441
rect 9677 9432 9689 9435
rect 9364 9404 9689 9432
rect 9364 9392 9370 9404
rect 9677 9401 9689 9404
rect 9723 9401 9735 9435
rect 10397 9432 10425 9472
rect 10597 9469 10609 9503
rect 10643 9500 10655 9503
rect 10870 9500 10876 9512
rect 10643 9472 10876 9500
rect 10643 9469 10655 9472
rect 10597 9463 10655 9469
rect 10870 9460 10876 9472
rect 10928 9460 10934 9512
rect 11882 9500 11888 9512
rect 11795 9472 11888 9500
rect 11882 9460 11888 9472
rect 11940 9500 11946 9512
rect 12342 9500 12348 9512
rect 11940 9472 12348 9500
rect 11940 9460 11946 9472
rect 12342 9460 12348 9472
rect 12400 9460 12406 9512
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9500 13783 9503
rect 13814 9500 13820 9512
rect 13771 9472 13820 9500
rect 13771 9469 13783 9472
rect 13725 9463 13783 9469
rect 13814 9460 13820 9472
rect 13872 9460 13878 9512
rect 11900 9432 11928 9460
rect 13924 9432 13952 9540
rect 14930 9537 14942 9540
rect 14976 9537 14988 9571
rect 14930 9531 14988 9537
rect 15102 9528 15108 9580
rect 15160 9528 15166 9580
rect 15194 9528 15200 9580
rect 15252 9568 15258 9580
rect 16025 9571 16083 9577
rect 16025 9568 16037 9571
rect 15252 9540 16037 9568
rect 15252 9528 15258 9540
rect 16025 9537 16037 9540
rect 16071 9568 16083 9571
rect 17034 9568 17040 9580
rect 16071 9540 17040 9568
rect 16071 9537 16083 9540
rect 16025 9531 16083 9537
rect 17034 9528 17040 9540
rect 17092 9528 17098 9580
rect 17793 9571 17851 9577
rect 17793 9537 17805 9571
rect 17839 9568 17851 9571
rect 18230 9568 18236 9580
rect 17839 9540 18236 9568
rect 17839 9537 17851 9540
rect 17793 9531 17851 9537
rect 18230 9528 18236 9540
rect 18288 9528 18294 9580
rect 20829 9571 20887 9577
rect 20829 9537 20841 9571
rect 20875 9568 20887 9571
rect 20990 9568 20996 9580
rect 20875 9540 20996 9568
rect 20875 9537 20887 9540
rect 20829 9531 20887 9537
rect 20990 9528 20996 9540
rect 21048 9528 21054 9580
rect 21100 9577 21128 9676
rect 21177 9673 21189 9676
rect 21223 9704 21235 9707
rect 21361 9707 21419 9713
rect 21361 9704 21373 9707
rect 21223 9676 21373 9704
rect 21223 9673 21235 9676
rect 21177 9667 21235 9673
rect 21361 9673 21373 9676
rect 21407 9673 21419 9707
rect 21361 9667 21419 9673
rect 21085 9571 21143 9577
rect 21085 9537 21097 9571
rect 21131 9537 21143 9571
rect 21085 9531 21143 9537
rect 15120 9500 15148 9528
rect 15841 9503 15899 9509
rect 15841 9500 15853 9503
rect 15120 9472 15853 9500
rect 15841 9469 15853 9472
rect 15887 9469 15899 9503
rect 18046 9500 18052 9512
rect 18007 9472 18052 9500
rect 15841 9463 15899 9469
rect 18046 9460 18052 9472
rect 18104 9500 18110 9512
rect 18141 9503 18199 9509
rect 18141 9500 18153 9503
rect 18104 9472 18153 9500
rect 18104 9460 18110 9472
rect 18141 9469 18153 9472
rect 18187 9469 18199 9503
rect 18141 9463 18199 9469
rect 16666 9432 16672 9444
rect 10397 9404 11928 9432
rect 13740 9404 13952 9432
rect 16627 9404 16672 9432
rect 9677 9395 9735 9401
rect 8757 9367 8815 9373
rect 8757 9364 8769 9367
rect 8536 9336 8769 9364
rect 8536 9324 8542 9336
rect 8757 9333 8769 9336
rect 8803 9333 8815 9367
rect 8757 9327 8815 9333
rect 9030 9324 9036 9376
rect 9088 9364 9094 9376
rect 9490 9364 9496 9376
rect 9088 9336 9496 9364
rect 9088 9324 9094 9336
rect 9490 9324 9496 9336
rect 9548 9324 9554 9376
rect 9766 9364 9772 9376
rect 9727 9336 9772 9364
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 9953 9367 10011 9373
rect 9953 9333 9965 9367
rect 9999 9364 10011 9367
rect 10134 9364 10140 9376
rect 9999 9336 10140 9364
rect 9999 9333 10011 9336
rect 9953 9327 10011 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10502 9324 10508 9376
rect 10560 9364 10566 9376
rect 10778 9364 10784 9376
rect 10560 9336 10784 9364
rect 10560 9324 10566 9336
rect 10778 9324 10784 9336
rect 10836 9364 10842 9376
rect 11057 9367 11115 9373
rect 11057 9364 11069 9367
rect 10836 9336 11069 9364
rect 10836 9324 10842 9336
rect 11057 9333 11069 9336
rect 11103 9333 11115 9367
rect 11698 9364 11704 9376
rect 11659 9336 11704 9364
rect 11057 9327 11115 9333
rect 11698 9324 11704 9336
rect 11756 9324 11762 9376
rect 12158 9324 12164 9376
rect 12216 9364 12222 9376
rect 12345 9367 12403 9373
rect 12345 9364 12357 9367
rect 12216 9336 12357 9364
rect 12216 9324 12222 9336
rect 12345 9333 12357 9336
rect 12391 9333 12403 9367
rect 12345 9327 12403 9333
rect 13446 9324 13452 9376
rect 13504 9364 13510 9376
rect 13740 9364 13768 9404
rect 16666 9392 16672 9404
rect 16724 9392 16730 9444
rect 19521 9435 19579 9441
rect 19521 9401 19533 9435
rect 19567 9432 19579 9435
rect 19567 9404 19840 9432
rect 19567 9401 19579 9404
rect 19521 9395 19579 9401
rect 13504 9336 13768 9364
rect 13817 9367 13875 9373
rect 13504 9324 13510 9336
rect 13817 9333 13829 9367
rect 13863 9364 13875 9367
rect 13906 9364 13912 9376
rect 13863 9336 13912 9364
rect 13863 9333 13875 9336
rect 13817 9327 13875 9333
rect 13906 9324 13912 9336
rect 13964 9324 13970 9376
rect 14274 9324 14280 9376
rect 14332 9364 14338 9376
rect 15289 9367 15347 9373
rect 15289 9364 15301 9367
rect 14332 9336 15301 9364
rect 14332 9324 14338 9336
rect 15289 9333 15301 9336
rect 15335 9333 15347 9367
rect 15289 9327 15347 9333
rect 17862 9324 17868 9376
rect 17920 9364 17926 9376
rect 19705 9367 19763 9373
rect 19705 9364 19717 9367
rect 17920 9336 19717 9364
rect 17920 9324 17926 9336
rect 19705 9333 19717 9336
rect 19751 9333 19763 9367
rect 19812 9364 19840 9404
rect 20714 9364 20720 9376
rect 19812 9336 20720 9364
rect 19705 9327 19763 9333
rect 20714 9324 20720 9336
rect 20772 9324 20778 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 2130 9160 2136 9172
rect 2091 9132 2136 9160
rect 2130 9120 2136 9132
rect 2188 9120 2194 9172
rect 2590 9160 2596 9172
rect 2240 9132 2596 9160
rect 1581 9095 1639 9101
rect 1581 9061 1593 9095
rect 1627 9092 1639 9095
rect 2240 9092 2268 9132
rect 2590 9120 2596 9132
rect 2648 9120 2654 9172
rect 3050 9160 3056 9172
rect 3011 9132 3056 9160
rect 3050 9120 3056 9132
rect 3108 9120 3114 9172
rect 3326 9160 3332 9172
rect 3160 9132 3332 9160
rect 2958 9092 2964 9104
rect 1627 9064 2268 9092
rect 2919 9064 2964 9092
rect 1627 9061 1639 9064
rect 1581 9055 1639 9061
rect 2958 9052 2964 9064
rect 3016 9052 3022 9104
rect 2409 9027 2467 9033
rect 2409 8993 2421 9027
rect 2455 9024 2467 9027
rect 3160 9024 3188 9132
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 3881 9163 3939 9169
rect 3881 9160 3893 9163
rect 3476 9132 3893 9160
rect 3476 9120 3482 9132
rect 3881 9129 3893 9132
rect 3927 9129 3939 9163
rect 5442 9160 5448 9172
rect 3881 9123 3939 9129
rect 4632 9132 5448 9160
rect 2455 8996 3188 9024
rect 2455 8993 2467 8996
rect 2409 8987 2467 8993
rect 4338 8984 4344 9036
rect 4396 9024 4402 9036
rect 4632 9033 4660 9132
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 6089 9163 6147 9169
rect 6089 9129 6101 9163
rect 6135 9160 6147 9163
rect 6546 9160 6552 9172
rect 6135 9132 6552 9160
rect 6135 9129 6147 9132
rect 6089 9123 6147 9129
rect 6546 9120 6552 9132
rect 6604 9120 6610 9172
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 8018 9160 8024 9172
rect 7800 9132 8024 9160
rect 7800 9120 7806 9132
rect 8018 9120 8024 9132
rect 8076 9160 8082 9172
rect 8076 9132 9536 9160
rect 8076 9120 8082 9132
rect 7009 9095 7067 9101
rect 7009 9092 7021 9095
rect 4724 9064 7021 9092
rect 4617 9027 4675 9033
rect 4617 9024 4629 9027
rect 4396 8996 4629 9024
rect 4396 8984 4402 8996
rect 4617 8993 4629 8996
rect 4663 8993 4675 9027
rect 4617 8987 4675 8993
rect 1394 8956 1400 8968
rect 1307 8928 1400 8956
rect 1394 8916 1400 8928
rect 1452 8916 1458 8968
rect 1670 8956 1676 8968
rect 1631 8928 1676 8956
rect 1670 8916 1676 8928
rect 1728 8916 1734 8968
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8956 2007 8959
rect 2498 8956 2504 8968
rect 1995 8928 2504 8956
rect 1995 8925 2007 8928
rect 1949 8919 2007 8925
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 2590 8916 2596 8968
rect 2648 8956 2654 8968
rect 3237 8959 3295 8965
rect 2648 8928 2693 8956
rect 2648 8916 2654 8928
rect 3237 8925 3249 8959
rect 3283 8925 3295 8959
rect 4062 8956 4068 8968
rect 4023 8928 4068 8956
rect 3237 8919 3295 8925
rect 1412 8888 1440 8916
rect 2774 8888 2780 8900
rect 1412 8860 2780 8888
rect 2774 8848 2780 8860
rect 2832 8848 2838 8900
rect 3252 8888 3280 8919
rect 4062 8916 4068 8928
rect 4120 8916 4126 8968
rect 4724 8888 4752 9064
rect 7009 9061 7021 9064
rect 7055 9061 7067 9095
rect 7009 9055 7067 9061
rect 8110 9052 8116 9104
rect 8168 9092 8174 9104
rect 9508 9092 9536 9132
rect 9582 9120 9588 9172
rect 9640 9160 9646 9172
rect 9677 9163 9735 9169
rect 9677 9160 9689 9163
rect 9640 9132 9689 9160
rect 9640 9120 9646 9132
rect 9677 9129 9689 9132
rect 9723 9129 9735 9163
rect 9677 9123 9735 9129
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 13630 9160 13636 9172
rect 9824 9132 13636 9160
rect 9824 9120 9830 9132
rect 13630 9120 13636 9132
rect 13688 9120 13694 9172
rect 16114 9160 16120 9172
rect 14108 9132 16120 9160
rect 10502 9092 10508 9104
rect 8168 9064 8524 9092
rect 9508 9064 10508 9092
rect 8168 9052 8174 9064
rect 8496 9036 8524 9064
rect 10502 9052 10508 9064
rect 10560 9052 10566 9104
rect 13446 9092 13452 9104
rect 13407 9064 13452 9092
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 13538 9052 13544 9104
rect 13596 9092 13602 9104
rect 14108 9092 14136 9132
rect 16114 9120 16120 9132
rect 16172 9120 16178 9172
rect 13596 9064 14136 9092
rect 13596 9052 13602 9064
rect 4801 9027 4859 9033
rect 4801 8993 4813 9027
rect 4847 9024 4859 9027
rect 5074 9024 5080 9036
rect 4847 8996 5080 9024
rect 4847 8993 4859 8996
rect 4801 8987 4859 8993
rect 5074 8984 5080 8996
rect 5132 8984 5138 9036
rect 5537 9027 5595 9033
rect 5537 8993 5549 9027
rect 5583 9024 5595 9027
rect 5718 9024 5724 9036
rect 5583 8996 5724 9024
rect 5583 8993 5595 8996
rect 5537 8987 5595 8993
rect 5718 8984 5724 8996
rect 5776 9024 5782 9036
rect 5902 9024 5908 9036
rect 5776 8996 5908 9024
rect 5776 8984 5782 8996
rect 5902 8984 5908 8996
rect 5960 8984 5966 9036
rect 6822 9024 6828 9036
rect 6783 8996 6828 9024
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 7653 9027 7711 9033
rect 7653 8993 7665 9027
rect 7699 9024 7711 9027
rect 8202 9024 8208 9036
rect 7699 8996 8208 9024
rect 7699 8993 7711 8996
rect 7653 8987 7711 8993
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 8478 9024 8484 9036
rect 8439 8996 8484 9024
rect 8478 8984 8484 8996
rect 8536 8984 8542 9036
rect 8570 8984 8576 9036
rect 8628 9024 8634 9036
rect 8754 9024 8760 9036
rect 8628 8996 8760 9024
rect 8628 8984 8634 8996
rect 8754 8984 8760 8996
rect 8812 8984 8818 9036
rect 10134 9024 10140 9036
rect 10095 8996 10140 9024
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 10318 9024 10324 9036
rect 10279 8996 10324 9024
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 10778 8984 10784 9036
rect 10836 9024 10842 9036
rect 11057 9027 11115 9033
rect 11057 9024 11069 9027
rect 10836 8996 11069 9024
rect 10836 8984 10842 8996
rect 11057 8993 11069 8996
rect 11103 8993 11115 9027
rect 11057 8987 11115 8993
rect 11698 8984 11704 9036
rect 11756 9024 11762 9036
rect 12069 9027 12127 9033
rect 12069 9024 12081 9027
rect 11756 8996 12081 9024
rect 11756 8984 11762 8996
rect 12069 8993 12081 8996
rect 12115 8993 12127 9027
rect 12069 8987 12127 8993
rect 4890 8956 4896 8968
rect 4851 8928 4896 8956
rect 4890 8916 4896 8928
rect 4948 8916 4954 8968
rect 9950 8956 9956 8968
rect 5092 8928 9956 8956
rect 3252 8860 4752 8888
rect 1857 8823 1915 8829
rect 1857 8789 1869 8823
rect 1903 8820 1915 8823
rect 1946 8820 1952 8832
rect 1903 8792 1952 8820
rect 1903 8789 1915 8792
rect 1857 8783 1915 8789
rect 1946 8780 1952 8792
rect 2004 8780 2010 8832
rect 2498 8820 2504 8832
rect 2459 8792 2504 8820
rect 2498 8780 2504 8792
rect 2556 8780 2562 8832
rect 5092 8820 5120 8928
rect 9950 8916 9956 8928
rect 10008 8916 10014 8968
rect 10502 8916 10508 8968
rect 10560 8956 10566 8968
rect 10965 8959 11023 8965
rect 10965 8956 10977 8959
rect 10560 8928 10977 8956
rect 10560 8916 10566 8928
rect 10965 8925 10977 8928
rect 11011 8925 11023 8959
rect 12084 8956 12112 8987
rect 13814 8956 13820 8968
rect 12084 8928 13820 8956
rect 10965 8919 11023 8925
rect 13814 8916 13820 8928
rect 13872 8956 13878 8968
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13872 8928 14105 8956
rect 13872 8916 13878 8928
rect 14093 8925 14105 8928
rect 14139 8956 14151 8959
rect 15194 8956 15200 8968
rect 14139 8928 15200 8956
rect 14139 8925 14151 8928
rect 14093 8919 14151 8925
rect 15194 8916 15200 8928
rect 15252 8956 15258 8968
rect 15565 8959 15623 8965
rect 15565 8956 15577 8959
rect 15252 8928 15577 8956
rect 15252 8916 15258 8928
rect 15565 8925 15577 8928
rect 15611 8956 15623 8959
rect 15746 8956 15752 8968
rect 15611 8928 15752 8956
rect 15611 8925 15623 8928
rect 15565 8919 15623 8925
rect 15746 8916 15752 8928
rect 15804 8956 15810 8968
rect 16301 8959 16359 8965
rect 16301 8956 16313 8959
rect 15804 8928 16313 8956
rect 15804 8916 15810 8928
rect 16301 8925 16313 8928
rect 16347 8956 16359 8959
rect 17773 8959 17831 8965
rect 17773 8956 17785 8959
rect 16347 8928 17785 8956
rect 16347 8925 16359 8928
rect 16301 8919 16359 8925
rect 17773 8925 17785 8928
rect 17819 8956 17831 8959
rect 18046 8956 18052 8968
rect 17819 8928 18052 8956
rect 17819 8925 17831 8928
rect 17773 8919 17831 8925
rect 18046 8916 18052 8928
rect 18104 8956 18110 8968
rect 18141 8959 18199 8965
rect 18141 8956 18153 8959
rect 18104 8928 18153 8956
rect 18104 8916 18110 8928
rect 18141 8925 18153 8928
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 20622 8916 20628 8968
rect 20680 8965 20686 8968
rect 20680 8956 20692 8965
rect 20680 8928 20725 8956
rect 20680 8919 20692 8928
rect 20680 8916 20686 8919
rect 20806 8916 20812 8968
rect 20864 8956 20870 8968
rect 20901 8959 20959 8965
rect 20901 8956 20913 8959
rect 20864 8928 20913 8956
rect 20864 8916 20870 8928
rect 20901 8925 20913 8928
rect 20947 8956 20959 8959
rect 20993 8959 21051 8965
rect 20993 8956 21005 8959
rect 20947 8928 21005 8956
rect 20947 8925 20959 8928
rect 20901 8919 20959 8925
rect 20993 8925 21005 8928
rect 21039 8925 21051 8959
rect 20993 8919 21051 8925
rect 5166 8848 5172 8900
rect 5224 8888 5230 8900
rect 5224 8860 6224 8888
rect 5224 8848 5230 8860
rect 5261 8823 5319 8829
rect 5261 8820 5273 8823
rect 5092 8792 5273 8820
rect 5261 8789 5273 8792
rect 5307 8789 5319 8823
rect 5261 8783 5319 8789
rect 5350 8780 5356 8832
rect 5408 8820 5414 8832
rect 5629 8823 5687 8829
rect 5629 8820 5641 8823
rect 5408 8792 5641 8820
rect 5408 8780 5414 8792
rect 5629 8789 5641 8792
rect 5675 8789 5687 8823
rect 5629 8783 5687 8789
rect 5718 8780 5724 8832
rect 5776 8820 5782 8832
rect 6196 8829 6224 8860
rect 7006 8848 7012 8900
rect 7064 8888 7070 8900
rect 7282 8888 7288 8900
rect 7064 8860 7288 8888
rect 7064 8848 7070 8860
rect 7282 8848 7288 8860
rect 7340 8848 7346 8900
rect 7377 8891 7435 8897
rect 7377 8857 7389 8891
rect 7423 8888 7435 8891
rect 7423 8860 7880 8888
rect 7423 8857 7435 8860
rect 7377 8851 7435 8857
rect 6181 8823 6239 8829
rect 5776 8792 5821 8820
rect 5776 8780 5782 8792
rect 6181 8789 6193 8823
rect 6227 8789 6239 8823
rect 6546 8820 6552 8832
rect 6507 8792 6552 8820
rect 6181 8783 6239 8789
rect 6546 8780 6552 8792
rect 6604 8780 6610 8832
rect 6638 8780 6644 8832
rect 6696 8820 6702 8832
rect 7469 8823 7527 8829
rect 6696 8792 6741 8820
rect 6696 8780 6702 8792
rect 7469 8789 7481 8823
rect 7515 8820 7527 8823
rect 7742 8820 7748 8832
rect 7515 8792 7748 8820
rect 7515 8789 7527 8792
rect 7469 8783 7527 8789
rect 7742 8780 7748 8792
rect 7800 8780 7806 8832
rect 7852 8829 7880 8860
rect 7926 8848 7932 8900
rect 7984 8888 7990 8900
rect 9766 8888 9772 8900
rect 7984 8860 9772 8888
rect 7984 8848 7990 8860
rect 9766 8848 9772 8860
rect 9824 8848 9830 8900
rect 10873 8891 10931 8897
rect 10873 8857 10885 8891
rect 10919 8888 10931 8891
rect 11333 8891 11391 8897
rect 11333 8888 11345 8891
rect 10919 8860 11345 8888
rect 10919 8857 10931 8860
rect 10873 8851 10931 8857
rect 11333 8857 11345 8860
rect 11379 8857 11391 8891
rect 11333 8851 11391 8857
rect 12336 8891 12394 8897
rect 12336 8857 12348 8891
rect 12382 8888 12394 8891
rect 12526 8888 12532 8900
rect 12382 8860 12532 8888
rect 12382 8857 12394 8860
rect 12336 8851 12394 8857
rect 12526 8848 12532 8860
rect 12584 8848 12590 8900
rect 14360 8891 14418 8897
rect 14360 8857 14372 8891
rect 14406 8888 14418 8891
rect 14458 8888 14464 8900
rect 14406 8860 14464 8888
rect 14406 8857 14418 8860
rect 14360 8851 14418 8857
rect 14458 8848 14464 8860
rect 14516 8848 14522 8900
rect 16568 8891 16626 8897
rect 16568 8857 16580 8891
rect 16614 8888 16626 8891
rect 16942 8888 16948 8900
rect 16614 8860 16948 8888
rect 16614 8857 16626 8860
rect 16568 8851 16626 8857
rect 16942 8848 16948 8860
rect 17000 8848 17006 8900
rect 7837 8823 7895 8829
rect 7837 8789 7849 8823
rect 7883 8789 7895 8823
rect 8202 8820 8208 8832
rect 8163 8792 8208 8820
rect 7837 8783 7895 8789
rect 8202 8780 8208 8792
rect 8260 8780 8266 8832
rect 8297 8823 8355 8829
rect 8297 8789 8309 8823
rect 8343 8820 8355 8823
rect 8570 8820 8576 8832
rect 8343 8792 8576 8820
rect 8343 8789 8355 8792
rect 8297 8783 8355 8789
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 8754 8820 8760 8832
rect 8715 8792 8760 8820
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 10042 8820 10048 8832
rect 10003 8792 10048 8820
rect 10042 8780 10048 8792
rect 10100 8780 10106 8832
rect 10502 8820 10508 8832
rect 10463 8792 10508 8820
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 13630 8820 13636 8832
rect 13591 8792 13636 8820
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 15194 8780 15200 8832
rect 15252 8820 15258 8832
rect 15473 8823 15531 8829
rect 15473 8820 15485 8823
rect 15252 8792 15485 8820
rect 15252 8780 15258 8792
rect 15473 8789 15485 8792
rect 15519 8820 15531 8823
rect 16390 8820 16396 8832
rect 15519 8792 16396 8820
rect 15519 8789 15531 8792
rect 15473 8783 15531 8789
rect 16390 8780 16396 8792
rect 16448 8780 16454 8832
rect 17494 8780 17500 8832
rect 17552 8820 17558 8832
rect 17681 8823 17739 8829
rect 17681 8820 17693 8823
rect 17552 8792 17693 8820
rect 17552 8780 17558 8792
rect 17681 8789 17693 8792
rect 17727 8789 17739 8823
rect 19518 8820 19524 8832
rect 19479 8792 19524 8820
rect 17681 8783 17739 8789
rect 19518 8780 19524 8792
rect 19576 8780 19582 8832
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 1670 8616 1676 8628
rect 1631 8588 1676 8616
rect 1670 8576 1676 8588
rect 1728 8576 1734 8628
rect 2038 8576 2044 8628
rect 2096 8616 2102 8628
rect 2685 8619 2743 8625
rect 2685 8616 2697 8619
rect 2096 8588 2697 8616
rect 2096 8576 2102 8588
rect 2685 8585 2697 8588
rect 2731 8585 2743 8619
rect 2685 8579 2743 8585
rect 2774 8576 2780 8628
rect 2832 8616 2838 8628
rect 3970 8616 3976 8628
rect 2832 8588 3976 8616
rect 2832 8576 2838 8588
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4341 8619 4399 8625
rect 4341 8616 4353 8619
rect 4212 8588 4353 8616
rect 4212 8576 4218 8588
rect 4341 8585 4353 8588
rect 4387 8585 4399 8619
rect 5994 8616 6000 8628
rect 4341 8579 4399 8585
rect 4724 8588 6000 8616
rect 4724 8548 4752 8588
rect 5994 8576 6000 8588
rect 6052 8576 6058 8628
rect 6181 8619 6239 8625
rect 6181 8585 6193 8619
rect 6227 8616 6239 8619
rect 6546 8616 6552 8628
rect 6227 8588 6552 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 6914 8576 6920 8628
rect 6972 8616 6978 8628
rect 8018 8616 8024 8628
rect 6972 8588 8024 8616
rect 6972 8576 6978 8588
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 8570 8616 8576 8628
rect 8531 8588 8576 8616
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 9950 8616 9956 8628
rect 9911 8588 9956 8616
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 10042 8576 10048 8628
rect 10100 8616 10106 8628
rect 10505 8619 10563 8625
rect 10505 8616 10517 8619
rect 10100 8588 10517 8616
rect 10100 8576 10106 8588
rect 10505 8585 10517 8588
rect 10551 8585 10563 8619
rect 10505 8579 10563 8585
rect 10778 8576 10784 8628
rect 10836 8616 10842 8628
rect 13538 8616 13544 8628
rect 10836 8588 13544 8616
rect 10836 8576 10842 8588
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 13814 8616 13820 8628
rect 13775 8588 13820 8616
rect 13814 8576 13820 8588
rect 13872 8616 13878 8628
rect 13909 8619 13967 8625
rect 13909 8616 13921 8619
rect 13872 8588 13921 8616
rect 13872 8576 13878 8588
rect 13909 8585 13921 8588
rect 13955 8585 13967 8619
rect 13909 8579 13967 8585
rect 15102 8576 15108 8628
rect 15160 8616 15166 8628
rect 15565 8619 15623 8625
rect 15565 8616 15577 8619
rect 15160 8588 15577 8616
rect 15160 8576 15166 8588
rect 15565 8585 15577 8588
rect 15611 8585 15623 8619
rect 15746 8616 15752 8628
rect 15707 8588 15752 8616
rect 15565 8579 15623 8585
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 16114 8576 16120 8628
rect 16172 8616 16178 8628
rect 17954 8616 17960 8628
rect 16172 8588 17960 8616
rect 16172 8576 16178 8588
rect 17954 8576 17960 8588
rect 18012 8576 18018 8628
rect 20622 8616 20628 8628
rect 18064 8588 20628 8616
rect 7285 8551 7343 8557
rect 1964 8520 3096 8548
rect 1394 8480 1400 8492
rect 1355 8452 1400 8480
rect 1394 8440 1400 8452
rect 1452 8440 1458 8492
rect 1964 8421 1992 8520
rect 2038 8440 2044 8492
rect 2096 8480 2102 8492
rect 2225 8483 2283 8489
rect 2225 8480 2237 8483
rect 2096 8452 2237 8480
rect 2096 8440 2102 8452
rect 2225 8449 2237 8452
rect 2271 8449 2283 8483
rect 2866 8480 2872 8492
rect 2827 8452 2872 8480
rect 2225 8443 2283 8449
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3068 8489 3096 8520
rect 4172 8520 4752 8548
rect 5092 8520 7236 8548
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3142 8480 3148 8492
rect 3099 8452 3148 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 1949 8415 2007 8421
rect 1949 8381 1961 8415
rect 1995 8381 2007 8415
rect 2130 8412 2136 8424
rect 2091 8384 2136 8412
rect 1949 8375 2007 8381
rect 2130 8372 2136 8384
rect 2188 8372 2194 8424
rect 2593 8347 2651 8353
rect 2593 8313 2605 8347
rect 2639 8344 2651 8347
rect 2774 8344 2780 8356
rect 2639 8316 2780 8344
rect 2639 8313 2651 8316
rect 2593 8307 2651 8313
rect 2774 8304 2780 8316
rect 2832 8304 2838 8356
rect 1581 8279 1639 8285
rect 1581 8245 1593 8279
rect 1627 8276 1639 8279
rect 4172 8276 4200 8520
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8449 4491 8483
rect 4433 8443 4491 8449
rect 4249 8415 4307 8421
rect 4249 8381 4261 8415
rect 4295 8412 4307 8415
rect 4338 8412 4344 8424
rect 4295 8384 4344 8412
rect 4295 8381 4307 8384
rect 4249 8375 4307 8381
rect 4338 8372 4344 8384
rect 4396 8372 4402 8424
rect 4448 8412 4476 8443
rect 4893 8415 4951 8421
rect 4893 8412 4905 8415
rect 4448 8384 4905 8412
rect 4893 8381 4905 8384
rect 4939 8381 4951 8415
rect 4893 8375 4951 8381
rect 1627 8248 4200 8276
rect 4801 8279 4859 8285
rect 1627 8245 1639 8248
rect 1581 8239 1639 8245
rect 4801 8245 4813 8279
rect 4847 8276 4859 8279
rect 5092 8276 5120 8520
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 5994 8480 6000 8492
rect 5859 8452 6000 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 6086 8440 6092 8492
rect 6144 8480 6150 8492
rect 6730 8480 6736 8492
rect 6144 8452 6736 8480
rect 6144 8440 6150 8452
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 7208 8480 7236 8520
rect 7285 8517 7297 8551
rect 7331 8548 7343 8551
rect 7466 8548 7472 8560
rect 7331 8520 7472 8548
rect 7331 8517 7343 8520
rect 7285 8511 7343 8517
rect 7466 8508 7472 8520
rect 7524 8508 7530 8560
rect 8113 8551 8171 8557
rect 8113 8517 8125 8551
rect 8159 8548 8171 8551
rect 9401 8551 9459 8557
rect 9401 8548 9413 8551
rect 8159 8520 9413 8548
rect 8159 8517 8171 8520
rect 8113 8511 8171 8517
rect 9401 8517 9413 8520
rect 9447 8517 9459 8551
rect 9401 8511 9459 8517
rect 9674 8508 9680 8560
rect 9732 8548 9738 8560
rect 9732 8520 9996 8548
rect 9732 8508 9738 8520
rect 8941 8483 8999 8489
rect 7208 8452 8616 8480
rect 5534 8412 5540 8424
rect 5495 8384 5540 8412
rect 5534 8372 5540 8384
rect 5592 8372 5598 8424
rect 5718 8412 5724 8424
rect 5679 8384 5724 8412
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 5902 8372 5908 8424
rect 5960 8412 5966 8424
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 5960 8384 6377 8412
rect 5960 8372 5966 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 7374 8412 7380 8424
rect 7335 8384 7380 8412
rect 6365 8375 6423 8381
rect 7374 8372 7380 8384
rect 7432 8372 7438 8424
rect 7561 8415 7619 8421
rect 7561 8381 7573 8415
rect 7607 8381 7619 8415
rect 7926 8412 7932 8424
rect 7887 8384 7932 8412
rect 7561 8375 7619 8381
rect 5166 8304 5172 8356
rect 5224 8344 5230 8356
rect 6917 8347 6975 8353
rect 6917 8344 6929 8347
rect 5224 8316 6929 8344
rect 5224 8304 5230 8316
rect 6917 8313 6929 8316
rect 6963 8313 6975 8347
rect 7576 8344 7604 8375
rect 7926 8372 7932 8384
rect 7984 8372 7990 8424
rect 8294 8412 8300 8424
rect 8128 8384 8300 8412
rect 8128 8344 8156 8384
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 7576 8316 8156 8344
rect 6917 8307 6975 8313
rect 8202 8304 8208 8356
rect 8260 8344 8266 8356
rect 8481 8347 8539 8353
rect 8481 8344 8493 8347
rect 8260 8316 8493 8344
rect 8260 8304 8266 8316
rect 8481 8313 8493 8316
rect 8527 8313 8539 8347
rect 8588 8344 8616 8452
rect 8941 8449 8953 8483
rect 8987 8449 8999 8483
rect 9766 8480 9772 8492
rect 8941 8443 8999 8449
rect 9232 8452 9772 8480
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 8956 8412 8984 8443
rect 8720 8384 8984 8412
rect 9033 8415 9091 8421
rect 8720 8372 8726 8384
rect 9033 8381 9045 8415
rect 9079 8412 9091 8415
rect 9122 8412 9128 8424
rect 9079 8384 9128 8412
rect 9079 8381 9091 8384
rect 9033 8375 9091 8381
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 9232 8421 9260 8452
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 9217 8415 9275 8421
rect 9217 8381 9229 8415
rect 9263 8381 9275 8415
rect 9858 8412 9864 8424
rect 9819 8384 9864 8412
rect 9217 8375 9275 8381
rect 9858 8372 9864 8384
rect 9916 8372 9922 8424
rect 9968 8412 9996 8520
rect 10134 8508 10140 8560
rect 10192 8548 10198 8560
rect 10192 8520 11652 8548
rect 10192 8508 10198 8520
rect 10042 8440 10048 8492
rect 10100 8480 10106 8492
rect 10873 8483 10931 8489
rect 10100 8452 10145 8480
rect 10100 8440 10106 8452
rect 10873 8449 10885 8483
rect 10919 8480 10931 8483
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 10919 8452 11529 8480
rect 10919 8449 10931 8452
rect 10873 8443 10931 8449
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 10965 8415 11023 8421
rect 10965 8412 10977 8415
rect 9968 8384 10977 8412
rect 10965 8381 10977 8384
rect 11011 8381 11023 8415
rect 10965 8375 11023 8381
rect 11057 8415 11115 8421
rect 11057 8381 11069 8415
rect 11103 8381 11115 8415
rect 11057 8375 11115 8381
rect 10042 8344 10048 8356
rect 8588 8316 10048 8344
rect 8481 8307 8539 8313
rect 10042 8304 10048 8316
rect 10100 8304 10106 8356
rect 10410 8344 10416 8356
rect 10371 8316 10416 8344
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 10870 8304 10876 8356
rect 10928 8344 10934 8356
rect 11072 8344 11100 8375
rect 10928 8316 11100 8344
rect 11624 8344 11652 8520
rect 12158 8440 12164 8492
rect 12216 8480 12222 8492
rect 13366 8483 13424 8489
rect 13366 8480 13378 8483
rect 12216 8452 13378 8480
rect 12216 8440 12222 8452
rect 13366 8449 13378 8452
rect 13412 8449 13424 8483
rect 13366 8443 13424 8449
rect 13633 8483 13691 8489
rect 13633 8449 13645 8483
rect 13679 8480 13691 8483
rect 13832 8480 13860 8576
rect 14918 8508 14924 8560
rect 14976 8548 14982 8560
rect 18064 8548 18092 8588
rect 20622 8576 20628 8588
rect 20680 8576 20686 8628
rect 20717 8551 20775 8557
rect 20717 8548 20729 8551
rect 14976 8520 18092 8548
rect 19168 8520 20729 8548
rect 14976 8508 14982 8520
rect 14185 8483 14243 8489
rect 14185 8480 14197 8483
rect 13679 8452 14197 8480
rect 13679 8449 13691 8452
rect 13633 8443 13691 8449
rect 14185 8449 14197 8452
rect 14231 8449 14243 8483
rect 14441 8483 14499 8489
rect 14441 8480 14453 8483
rect 14185 8443 14243 8449
rect 14292 8452 14453 8480
rect 13722 8372 13728 8424
rect 13780 8412 13786 8424
rect 14292 8412 14320 8452
rect 14441 8449 14453 8452
rect 14487 8449 14499 8483
rect 14441 8443 14499 8449
rect 18046 8440 18052 8492
rect 18104 8480 18110 8492
rect 19168 8489 19196 8520
rect 20717 8517 20729 8520
rect 20763 8548 20775 8551
rect 20806 8548 20812 8560
rect 20763 8520 20812 8548
rect 20763 8517 20775 8520
rect 20717 8511 20775 8517
rect 20806 8508 20812 8520
rect 20864 8508 20870 8560
rect 19426 8489 19432 8492
rect 19153 8483 19211 8489
rect 19153 8480 19165 8483
rect 18104 8452 19165 8480
rect 18104 8440 18110 8452
rect 19153 8449 19165 8452
rect 19199 8449 19211 8483
rect 19420 8480 19432 8489
rect 19387 8452 19432 8480
rect 19153 8443 19211 8449
rect 19420 8443 19432 8452
rect 19426 8440 19432 8443
rect 19484 8440 19490 8492
rect 13780 8384 14320 8412
rect 13780 8372 13786 8384
rect 12253 8347 12311 8353
rect 12253 8344 12265 8347
rect 11624 8316 12265 8344
rect 10928 8304 10934 8316
rect 12253 8313 12265 8316
rect 12299 8313 12311 8347
rect 12253 8307 12311 8313
rect 13630 8304 13636 8356
rect 13688 8344 13694 8356
rect 18506 8344 18512 8356
rect 13688 8316 14228 8344
rect 13688 8304 13694 8316
rect 4847 8248 5120 8276
rect 5261 8279 5319 8285
rect 4847 8245 4859 8248
rect 4801 8239 4859 8245
rect 5261 8245 5273 8279
rect 5307 8276 5319 8279
rect 5442 8276 5448 8288
rect 5307 8248 5448 8276
rect 5307 8245 5319 8248
rect 5261 8239 5319 8245
rect 5442 8236 5448 8248
rect 5500 8276 5506 8288
rect 7650 8276 7656 8288
rect 5500 8248 7656 8276
rect 5500 8236 5506 8248
rect 7650 8236 7656 8248
rect 7708 8236 7714 8288
rect 8110 8236 8116 8288
rect 8168 8276 8174 8288
rect 12710 8276 12716 8288
rect 8168 8248 12716 8276
rect 8168 8236 8174 8248
rect 12710 8236 12716 8248
rect 12768 8236 12774 8288
rect 14200 8276 14228 8316
rect 15120 8316 18512 8344
rect 15120 8276 15148 8316
rect 18506 8304 18512 8316
rect 18564 8304 18570 8356
rect 14200 8248 15148 8276
rect 20438 8236 20444 8288
rect 20496 8276 20502 8288
rect 20533 8279 20591 8285
rect 20533 8276 20545 8279
rect 20496 8248 20545 8276
rect 20496 8236 20502 8248
rect 20533 8245 20545 8248
rect 20579 8245 20591 8279
rect 20533 8239 20591 8245
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 1762 8032 1768 8084
rect 1820 8072 1826 8084
rect 2593 8075 2651 8081
rect 2593 8072 2605 8075
rect 1820 8044 2605 8072
rect 1820 8032 1826 8044
rect 2593 8041 2605 8044
rect 2639 8041 2651 8075
rect 2593 8035 2651 8041
rect 3878 8032 3884 8084
rect 3936 8072 3942 8084
rect 5445 8075 5503 8081
rect 5445 8072 5457 8075
rect 3936 8044 5457 8072
rect 3936 8032 3942 8044
rect 5445 8041 5457 8044
rect 5491 8041 5503 8075
rect 5445 8035 5503 8041
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 6457 8075 6515 8081
rect 6457 8072 6469 8075
rect 5776 8044 6469 8072
rect 5776 8032 5782 8044
rect 6457 8041 6469 8044
rect 6503 8041 6515 8075
rect 6457 8035 6515 8041
rect 6914 8032 6920 8084
rect 6972 8072 6978 8084
rect 7561 8075 7619 8081
rect 7561 8072 7573 8075
rect 6972 8044 7573 8072
rect 6972 8032 6978 8044
rect 7561 8041 7573 8044
rect 7607 8041 7619 8075
rect 7561 8035 7619 8041
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 7837 8075 7895 8081
rect 7837 8072 7849 8075
rect 7800 8044 7849 8072
rect 7800 8032 7806 8044
rect 7837 8041 7849 8044
rect 7883 8041 7895 8075
rect 7837 8035 7895 8041
rect 8018 8032 8024 8084
rect 8076 8072 8082 8084
rect 8665 8075 8723 8081
rect 8665 8072 8677 8075
rect 8076 8044 8677 8072
rect 8076 8032 8082 8044
rect 8665 8041 8677 8044
rect 8711 8072 8723 8075
rect 9122 8072 9128 8084
rect 8711 8044 9128 8072
rect 8711 8041 8723 8044
rect 8665 8035 8723 8041
rect 9122 8032 9128 8044
rect 9180 8032 9186 8084
rect 12802 8072 12808 8084
rect 11992 8044 12808 8072
rect 1581 8007 1639 8013
rect 1581 7973 1593 8007
rect 1627 8004 1639 8007
rect 2406 8004 2412 8016
rect 1627 7976 2412 8004
rect 1627 7973 1639 7976
rect 1581 7967 1639 7973
rect 2406 7964 2412 7976
rect 2464 7964 2470 8016
rect 2501 8007 2559 8013
rect 2501 7973 2513 8007
rect 2547 8004 2559 8007
rect 4890 8004 4896 8016
rect 2547 7976 4896 8004
rect 2547 7973 2559 7976
rect 2501 7967 2559 7973
rect 4890 7964 4896 7976
rect 4948 7964 4954 8016
rect 4982 7964 4988 8016
rect 5040 8004 5046 8016
rect 6086 8004 6092 8016
rect 5040 7976 5672 8004
rect 6047 7976 6092 8004
rect 5040 7964 5046 7976
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7936 2007 7939
rect 2869 7939 2927 7945
rect 2869 7936 2881 7939
rect 1995 7908 2881 7936
rect 1995 7905 2007 7908
rect 1949 7899 2007 7905
rect 2869 7905 2881 7908
rect 2915 7936 2927 7939
rect 5442 7936 5448 7948
rect 2915 7908 5448 7936
rect 2915 7905 2927 7908
rect 2869 7899 2927 7905
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 5644 7936 5672 7976
rect 6086 7964 6092 7976
rect 6144 7964 6150 8016
rect 11885 8007 11943 8013
rect 11885 8004 11897 8007
rect 7024 7976 11897 8004
rect 5718 7936 5724 7948
rect 5631 7908 5724 7936
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 7024 7936 7052 7976
rect 11885 7973 11897 7976
rect 11931 7973 11943 8007
rect 11885 7967 11943 7973
rect 6104 7908 7052 7936
rect 7101 7939 7159 7945
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 2590 7868 2596 7880
rect 2056 7840 2596 7868
rect 2056 7809 2084 7840
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7837 2835 7871
rect 2777 7831 2835 7837
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7837 5687 7871
rect 6104 7844 6132 7908
rect 7101 7905 7113 7939
rect 7147 7936 7159 7939
rect 7190 7936 7196 7948
rect 7147 7908 7196 7936
rect 7147 7905 7159 7908
rect 7101 7899 7159 7905
rect 7190 7896 7196 7908
rect 7248 7936 7254 7948
rect 8202 7936 8208 7948
rect 7248 7908 8208 7936
rect 7248 7896 7254 7908
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 8478 7936 8484 7948
rect 8439 7908 8484 7936
rect 8478 7896 8484 7908
rect 8536 7896 8542 7948
rect 10042 7896 10048 7948
rect 10100 7936 10106 7948
rect 10318 7936 10324 7948
rect 10100 7908 10324 7936
rect 10100 7896 10106 7908
rect 10318 7896 10324 7908
rect 10376 7896 10382 7948
rect 10413 7939 10471 7945
rect 10413 7905 10425 7939
rect 10459 7936 10471 7939
rect 10962 7936 10968 7948
rect 10459 7908 10968 7936
rect 10459 7905 10471 7908
rect 10413 7899 10471 7905
rect 10962 7896 10968 7908
rect 11020 7896 11026 7948
rect 11241 7939 11299 7945
rect 11241 7936 11253 7939
rect 11072 7908 11253 7936
rect 11072 7880 11100 7908
rect 11241 7905 11253 7908
rect 11287 7936 11299 7939
rect 11992 7936 12020 8044
rect 12802 8032 12808 8044
rect 12860 8032 12866 8084
rect 14550 8032 14556 8084
rect 14608 8072 14614 8084
rect 14829 8075 14887 8081
rect 14829 8072 14841 8075
rect 14608 8044 14841 8072
rect 14608 8032 14614 8044
rect 14829 8041 14841 8044
rect 14875 8072 14887 8075
rect 15102 8072 15108 8084
rect 14875 8044 15108 8072
rect 14875 8041 14887 8044
rect 14829 8035 14887 8041
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 17586 8032 17592 8084
rect 17644 8072 17650 8084
rect 19429 8075 19487 8081
rect 19429 8072 19441 8075
rect 17644 8044 19441 8072
rect 17644 8032 17650 8044
rect 19429 8041 19441 8044
rect 19475 8072 19487 8075
rect 20162 8072 20168 8084
rect 19475 8044 20168 8072
rect 19475 8041 19487 8044
rect 19429 8035 19487 8041
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 20806 8032 20812 8084
rect 20864 8072 20870 8084
rect 20901 8075 20959 8081
rect 20901 8072 20913 8075
rect 20864 8044 20913 8072
rect 20864 8032 20870 8044
rect 20901 8041 20913 8044
rect 20947 8041 20959 8075
rect 20901 8035 20959 8041
rect 14369 8007 14427 8013
rect 14369 8004 14381 8007
rect 11287 7908 12020 7936
rect 12268 7976 14381 8004
rect 11287 7905 11299 7908
rect 11241 7899 11299 7905
rect 5629 7831 5687 7837
rect 2041 7803 2099 7809
rect 2041 7769 2053 7803
rect 2087 7769 2099 7803
rect 2041 7763 2099 7769
rect 2133 7803 2191 7809
rect 2133 7769 2145 7803
rect 2179 7800 2191 7803
rect 2682 7800 2688 7812
rect 2179 7772 2688 7800
rect 2179 7769 2191 7772
rect 2133 7763 2191 7769
rect 2682 7760 2688 7772
rect 2740 7760 2746 7812
rect 2792 7800 2820 7831
rect 5166 7800 5172 7812
rect 2792 7772 5172 7800
rect 5166 7760 5172 7772
rect 5224 7760 5230 7812
rect 5644 7800 5672 7831
rect 6012 7816 6132 7844
rect 6273 7871 6331 7877
rect 6273 7837 6285 7871
rect 6319 7868 6331 7871
rect 6546 7868 6552 7880
rect 6319 7840 6552 7868
rect 6319 7837 6331 7840
rect 6273 7831 6331 7837
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 8662 7868 8668 7880
rect 6840 7840 8668 7868
rect 6012 7800 6040 7816
rect 5644 7772 6040 7800
rect 6362 7760 6368 7812
rect 6420 7800 6426 7812
rect 6840 7809 6868 7840
rect 8662 7828 8668 7840
rect 8720 7828 8726 7880
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 10137 7871 10195 7877
rect 9180 7840 9674 7868
rect 9180 7828 9186 7840
rect 6825 7803 6883 7809
rect 6825 7800 6837 7803
rect 6420 7772 6837 7800
rect 6420 7760 6426 7772
rect 6825 7769 6837 7772
rect 6871 7769 6883 7803
rect 8018 7800 8024 7812
rect 6825 7763 6883 7769
rect 6932 7772 8024 7800
rect 1946 7692 1952 7744
rect 2004 7732 2010 7744
rect 4982 7732 4988 7744
rect 2004 7704 4988 7732
rect 2004 7692 2010 7704
rect 4982 7692 4988 7704
rect 5040 7692 5046 7744
rect 5902 7692 5908 7744
rect 5960 7732 5966 7744
rect 6932 7741 6960 7772
rect 8018 7760 8024 7772
rect 8076 7760 8082 7812
rect 8205 7803 8263 7809
rect 8205 7769 8217 7803
rect 8251 7800 8263 7803
rect 9306 7800 9312 7812
rect 8251 7772 9312 7800
rect 8251 7769 8263 7772
rect 8205 7763 8263 7769
rect 9306 7760 9312 7772
rect 9364 7760 9370 7812
rect 9646 7800 9674 7840
rect 10137 7837 10149 7871
rect 10183 7868 10195 7871
rect 10502 7868 10508 7880
rect 10183 7840 10508 7868
rect 10183 7837 10195 7840
rect 10137 7831 10195 7837
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 11054 7828 11060 7880
rect 11112 7828 11118 7880
rect 11330 7868 11336 7880
rect 11291 7840 11336 7868
rect 11330 7828 11336 7840
rect 11388 7828 11394 7880
rect 12268 7868 12296 7976
rect 14369 7973 14381 7976
rect 14415 8004 14427 8007
rect 14734 8004 14740 8016
rect 14415 7976 14740 8004
rect 14415 7973 14427 7976
rect 14369 7967 14427 7973
rect 14734 7964 14740 7976
rect 14792 7964 14798 8016
rect 19794 8004 19800 8016
rect 16684 7976 19800 8004
rect 12342 7896 12348 7948
rect 12400 7936 12406 7948
rect 12437 7939 12495 7945
rect 12437 7936 12449 7939
rect 12400 7908 12449 7936
rect 12400 7896 12406 7908
rect 12437 7905 12449 7908
rect 12483 7905 12495 7939
rect 12802 7936 12808 7948
rect 12715 7908 12808 7936
rect 12437 7899 12495 7905
rect 12802 7896 12808 7908
rect 12860 7936 12866 7948
rect 16684 7945 16712 7976
rect 19794 7964 19800 7976
rect 19852 7964 19858 8016
rect 20824 7945 20852 8032
rect 16669 7939 16727 7945
rect 12860 7908 16611 7936
rect 12860 7896 12866 7908
rect 11624 7840 12296 7868
rect 9646 7772 11100 7800
rect 6917 7735 6975 7741
rect 6917 7732 6929 7735
rect 5960 7704 6929 7732
rect 5960 7692 5966 7704
rect 6917 7701 6929 7704
rect 6963 7701 6975 7735
rect 7282 7732 7288 7744
rect 7243 7704 7288 7732
rect 6917 7695 6975 7701
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 8297 7735 8355 7741
rect 8297 7701 8309 7735
rect 8343 7732 8355 7735
rect 8386 7732 8392 7744
rect 8343 7704 8392 7732
rect 8343 7701 8355 7704
rect 8297 7695 8355 7701
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 9766 7732 9772 7744
rect 9727 7704 9772 7732
rect 9766 7692 9772 7704
rect 9824 7692 9830 7744
rect 10226 7692 10232 7744
rect 10284 7732 10290 7744
rect 11072 7732 11100 7772
rect 11146 7760 11152 7812
rect 11204 7800 11210 7812
rect 11425 7803 11483 7809
rect 11425 7800 11437 7803
rect 11204 7772 11437 7800
rect 11204 7760 11210 7772
rect 11425 7769 11437 7772
rect 11471 7769 11483 7803
rect 11425 7763 11483 7769
rect 11624 7732 11652 7840
rect 12526 7828 12532 7880
rect 12584 7828 12590 7880
rect 12710 7828 12716 7880
rect 12768 7868 12774 7880
rect 15286 7868 15292 7880
rect 12768 7840 15292 7868
rect 12768 7828 12774 7840
rect 15286 7828 15292 7840
rect 15344 7828 15350 7880
rect 15749 7871 15807 7877
rect 15749 7837 15761 7871
rect 15795 7868 15807 7871
rect 16583 7868 16611 7908
rect 16669 7905 16681 7939
rect 16715 7905 16727 7939
rect 18509 7939 18567 7945
rect 16669 7899 16727 7905
rect 16776 7908 18460 7936
rect 16776 7868 16804 7908
rect 18325 7871 18383 7877
rect 18325 7868 18337 7871
rect 15795 7840 16528 7868
rect 16583 7840 16804 7868
rect 17512 7840 18337 7868
rect 15795 7837 15807 7840
rect 15749 7831 15807 7837
rect 12544 7800 12572 7828
rect 13722 7800 13728 7812
rect 12544 7772 13728 7800
rect 13722 7760 13728 7772
rect 13780 7760 13786 7812
rect 16393 7803 16451 7809
rect 16393 7800 16405 7803
rect 15856 7772 16405 7800
rect 11790 7732 11796 7744
rect 10284 7704 10329 7732
rect 11072 7704 11652 7732
rect 11751 7704 11796 7732
rect 10284 7692 10290 7704
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 12066 7692 12072 7744
rect 12124 7732 12130 7744
rect 12253 7735 12311 7741
rect 12253 7732 12265 7735
rect 12124 7704 12265 7732
rect 12124 7692 12130 7704
rect 12253 7701 12265 7704
rect 12299 7701 12311 7735
rect 12253 7695 12311 7701
rect 12345 7735 12403 7741
rect 12345 7701 12357 7735
rect 12391 7732 12403 7735
rect 12526 7732 12532 7744
rect 12391 7704 12532 7732
rect 12391 7701 12403 7704
rect 12345 7695 12403 7701
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 14274 7732 14280 7744
rect 14235 7704 14280 7732
rect 14274 7692 14280 7704
rect 14332 7692 14338 7744
rect 15746 7692 15752 7744
rect 15804 7732 15810 7744
rect 15856 7741 15884 7772
rect 16393 7769 16405 7772
rect 16439 7769 16451 7803
rect 16393 7763 16451 7769
rect 15841 7735 15899 7741
rect 15841 7732 15853 7735
rect 15804 7704 15853 7732
rect 15804 7692 15810 7704
rect 15841 7701 15853 7704
rect 15887 7701 15899 7735
rect 16022 7732 16028 7744
rect 15983 7704 16028 7732
rect 15841 7695 15899 7701
rect 16022 7692 16028 7704
rect 16080 7692 16086 7744
rect 16500 7741 16528 7840
rect 16485 7735 16543 7741
rect 16485 7701 16497 7735
rect 16531 7732 16543 7735
rect 17310 7732 17316 7744
rect 16531 7704 17316 7732
rect 16531 7701 16543 7704
rect 16485 7695 16543 7701
rect 17310 7692 17316 7704
rect 17368 7692 17374 7744
rect 17402 7692 17408 7744
rect 17460 7732 17466 7744
rect 17512 7741 17540 7840
rect 18325 7837 18337 7840
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 18233 7803 18291 7809
rect 18233 7800 18245 7803
rect 17696 7772 18245 7800
rect 17696 7744 17724 7772
rect 18233 7769 18245 7772
rect 18279 7769 18291 7803
rect 18432 7800 18460 7908
rect 18509 7905 18521 7939
rect 18555 7905 18567 7939
rect 18509 7899 18567 7905
rect 20809 7939 20867 7945
rect 20809 7905 20821 7939
rect 20855 7905 20867 7939
rect 20809 7899 20867 7905
rect 18524 7868 18552 7899
rect 21542 7868 21548 7880
rect 18524 7840 21548 7868
rect 21542 7828 21548 7840
rect 21600 7828 21606 7880
rect 18506 7800 18512 7812
rect 18432 7772 18512 7800
rect 18233 7763 18291 7769
rect 18506 7760 18512 7772
rect 18564 7800 18570 7812
rect 20530 7800 20536 7812
rect 20588 7809 20594 7812
rect 18564 7772 20536 7800
rect 18564 7760 18570 7772
rect 20530 7760 20536 7772
rect 20588 7800 20600 7809
rect 21085 7803 21143 7809
rect 21085 7800 21097 7803
rect 20588 7772 21097 7800
rect 20588 7763 20600 7772
rect 21085 7769 21097 7772
rect 21131 7769 21143 7803
rect 21085 7763 21143 7769
rect 20588 7760 20594 7763
rect 17497 7735 17555 7741
rect 17497 7732 17509 7735
rect 17460 7704 17509 7732
rect 17460 7692 17466 7704
rect 17497 7701 17509 7704
rect 17543 7701 17555 7735
rect 17678 7732 17684 7744
rect 17639 7704 17684 7732
rect 17497 7695 17555 7701
rect 17678 7692 17684 7704
rect 17736 7692 17742 7744
rect 17862 7732 17868 7744
rect 17823 7704 17868 7732
rect 17862 7692 17868 7704
rect 17920 7692 17926 7744
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 1486 7488 1492 7540
rect 1544 7528 1550 7540
rect 2133 7531 2191 7537
rect 2133 7528 2145 7531
rect 1544 7500 2145 7528
rect 1544 7488 1550 7500
rect 2133 7497 2145 7500
rect 2179 7497 2191 7531
rect 2133 7491 2191 7497
rect 2406 7488 2412 7540
rect 2464 7528 2470 7540
rect 4893 7531 4951 7537
rect 4893 7528 4905 7531
rect 2464 7500 4905 7528
rect 2464 7488 2470 7500
rect 4893 7497 4905 7500
rect 4939 7528 4951 7531
rect 5626 7528 5632 7540
rect 4939 7500 5632 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 6181 7531 6239 7537
rect 6181 7497 6193 7531
rect 6227 7528 6239 7531
rect 6638 7528 6644 7540
rect 6227 7500 6644 7528
rect 6227 7497 6239 7500
rect 6181 7491 6239 7497
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 6825 7531 6883 7537
rect 6825 7497 6837 7531
rect 6871 7528 6883 7531
rect 7282 7528 7288 7540
rect 6871 7500 7288 7528
rect 6871 7497 6883 7500
rect 6825 7491 6883 7497
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 7466 7528 7472 7540
rect 7427 7500 7472 7528
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 9033 7531 9091 7537
rect 9033 7497 9045 7531
rect 9079 7528 9091 7531
rect 9585 7531 9643 7537
rect 9585 7528 9597 7531
rect 9079 7500 9597 7528
rect 9079 7497 9091 7500
rect 9033 7491 9091 7497
rect 9585 7497 9597 7500
rect 9631 7497 9643 7531
rect 10505 7531 10563 7537
rect 10505 7528 10517 7531
rect 9585 7491 9643 7497
rect 10336 7500 10517 7528
rect 1578 7420 1584 7472
rect 1636 7460 1642 7472
rect 1949 7463 2007 7469
rect 1949 7460 1961 7463
rect 1636 7432 1961 7460
rect 1636 7420 1642 7432
rect 1949 7429 1961 7432
rect 1995 7429 2007 7463
rect 1949 7423 2007 7429
rect 4985 7463 5043 7469
rect 4985 7429 4997 7463
rect 5031 7460 5043 7463
rect 5258 7460 5264 7472
rect 5031 7432 5264 7460
rect 5031 7429 5043 7432
rect 4985 7423 5043 7429
rect 5258 7420 5264 7432
rect 5316 7420 5322 7472
rect 5442 7420 5448 7472
rect 5500 7460 5506 7472
rect 8202 7460 8208 7472
rect 5500 7432 8208 7460
rect 5500 7420 5506 7432
rect 8202 7420 8208 7432
rect 8260 7420 8266 7472
rect 9493 7463 9551 7469
rect 8496 7432 9444 7460
rect 1394 7392 1400 7404
rect 1355 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7352 1458 7404
rect 1670 7392 1676 7404
rect 1631 7364 1676 7392
rect 1670 7352 1676 7364
rect 1728 7392 1734 7404
rect 2317 7395 2375 7401
rect 2317 7392 2329 7395
rect 1728 7364 2329 7392
rect 1728 7352 1734 7364
rect 2317 7361 2329 7364
rect 2363 7361 2375 7395
rect 2317 7355 2375 7361
rect 4890 7352 4896 7404
rect 4948 7392 4954 7404
rect 5626 7392 5632 7404
rect 4948 7364 5632 7392
rect 4948 7352 4954 7364
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 5810 7392 5816 7404
rect 5771 7364 5816 7392
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 7190 7392 7196 7404
rect 7116 7364 7196 7392
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7324 4859 7327
rect 4982 7324 4988 7336
rect 4847 7296 4988 7324
rect 4847 7293 4859 7296
rect 4801 7287 4859 7293
rect 4982 7284 4988 7296
rect 5040 7284 5046 7336
rect 5534 7324 5540 7336
rect 5495 7296 5540 7324
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7324 5779 7327
rect 5902 7324 5908 7336
rect 5767 7296 5908 7324
rect 5767 7293 5779 7296
rect 5721 7287 5779 7293
rect 5902 7284 5908 7296
rect 5960 7284 5966 7336
rect 6270 7284 6276 7336
rect 6328 7324 6334 7336
rect 6914 7324 6920 7336
rect 6328 7296 6920 7324
rect 6328 7284 6334 7296
rect 6914 7284 6920 7296
rect 6972 7284 6978 7336
rect 7116 7333 7144 7364
rect 7190 7352 7196 7364
rect 7248 7392 7254 7404
rect 7285 7395 7343 7401
rect 7285 7392 7297 7395
rect 7248 7364 7297 7392
rect 7248 7352 7254 7364
rect 7285 7361 7297 7364
rect 7331 7361 7343 7395
rect 7834 7392 7840 7404
rect 7795 7364 7840 7392
rect 7285 7355 7343 7361
rect 7834 7352 7840 7364
rect 7892 7352 7898 7404
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7392 7987 7395
rect 8294 7392 8300 7404
rect 7975 7364 8300 7392
rect 7975 7361 7987 7364
rect 7929 7355 7987 7361
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7293 7159 7327
rect 8110 7324 8116 7336
rect 8071 7296 8116 7324
rect 7101 7287 7159 7293
rect 8110 7284 8116 7296
rect 8168 7284 8174 7336
rect 8496 7333 8524 7432
rect 8662 7392 8668 7404
rect 8623 7364 8668 7392
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 9416 7392 9444 7432
rect 9493 7429 9505 7463
rect 9539 7460 9551 7463
rect 10336 7460 10364 7500
rect 10505 7497 10517 7500
rect 10551 7497 10563 7531
rect 12066 7528 12072 7540
rect 12027 7500 12072 7528
rect 10505 7491 10563 7497
rect 12066 7488 12072 7500
rect 12124 7488 12130 7540
rect 13446 7528 13452 7540
rect 13407 7500 13452 7528
rect 13446 7488 13452 7500
rect 13504 7488 13510 7540
rect 14274 7488 14280 7540
rect 14332 7528 14338 7540
rect 14645 7531 14703 7537
rect 14645 7528 14657 7531
rect 14332 7500 14657 7528
rect 14332 7488 14338 7500
rect 14645 7497 14657 7500
rect 14691 7497 14703 7531
rect 14645 7491 14703 7497
rect 14734 7488 14740 7540
rect 14792 7528 14798 7540
rect 14792 7500 14837 7528
rect 14792 7488 14798 7500
rect 15102 7488 15108 7540
rect 15160 7528 15166 7540
rect 15565 7531 15623 7537
rect 15565 7528 15577 7531
rect 15160 7500 15577 7528
rect 15160 7488 15166 7500
rect 15565 7497 15577 7500
rect 15611 7528 15623 7531
rect 17218 7528 17224 7540
rect 15611 7500 17224 7528
rect 15611 7497 15623 7500
rect 15565 7491 15623 7497
rect 17218 7488 17224 7500
rect 17276 7488 17282 7540
rect 19337 7531 19395 7537
rect 19337 7497 19349 7531
rect 19383 7497 19395 7531
rect 20806 7528 20812 7540
rect 20767 7500 20812 7528
rect 19337 7491 19395 7497
rect 10962 7460 10968 7472
rect 9539 7432 10364 7460
rect 10923 7432 10968 7460
rect 9539 7429 9551 7432
rect 9493 7423 9551 7429
rect 10962 7420 10968 7432
rect 11020 7420 11026 7472
rect 18230 7460 18236 7472
rect 11624 7432 18236 7460
rect 10873 7395 10931 7401
rect 9416 7364 10824 7392
rect 8481 7327 8539 7333
rect 8481 7293 8493 7327
rect 8527 7293 8539 7327
rect 8481 7287 8539 7293
rect 8573 7327 8631 7333
rect 8573 7293 8585 7327
rect 8619 7293 8631 7327
rect 8573 7287 8631 7293
rect 1578 7256 1584 7268
rect 1539 7228 1584 7256
rect 1578 7216 1584 7228
rect 1636 7216 1642 7268
rect 1857 7259 1915 7265
rect 1857 7225 1869 7259
rect 1903 7256 1915 7259
rect 5074 7256 5080 7268
rect 1903 7228 5080 7256
rect 1903 7225 1915 7228
rect 1857 7219 1915 7225
rect 5074 7216 5080 7228
rect 5132 7216 5138 7268
rect 5166 7216 5172 7268
rect 5224 7256 5230 7268
rect 5224 7228 5948 7256
rect 5224 7216 5230 7228
rect 5353 7191 5411 7197
rect 5353 7157 5365 7191
rect 5399 7188 5411 7191
rect 5442 7188 5448 7200
rect 5399 7160 5448 7188
rect 5399 7157 5411 7160
rect 5353 7151 5411 7157
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 5920 7188 5948 7228
rect 5994 7216 6000 7268
rect 6052 7256 6058 7268
rect 6457 7259 6515 7265
rect 6457 7256 6469 7259
rect 6052 7228 6469 7256
rect 6052 7216 6058 7228
rect 6457 7225 6469 7228
rect 6503 7225 6515 7259
rect 8588 7256 8616 7287
rect 9398 7284 9404 7336
rect 9456 7324 9462 7336
rect 9677 7327 9735 7333
rect 9677 7324 9689 7327
rect 9456 7296 9689 7324
rect 9456 7284 9462 7296
rect 9677 7293 9689 7296
rect 9723 7293 9735 7327
rect 10796 7324 10824 7364
rect 10873 7361 10885 7395
rect 10919 7392 10931 7395
rect 11517 7395 11575 7401
rect 11517 7392 11529 7395
rect 10919 7364 11529 7392
rect 10919 7361 10931 7364
rect 10873 7355 10931 7361
rect 11517 7361 11529 7364
rect 11563 7361 11575 7395
rect 11517 7355 11575 7361
rect 11057 7327 11115 7333
rect 11057 7324 11069 7327
rect 10796 7296 11069 7324
rect 9677 7287 9735 7293
rect 11057 7293 11069 7296
rect 11103 7324 11115 7327
rect 11624 7324 11652 7432
rect 18230 7420 18236 7432
rect 18288 7460 18294 7472
rect 19352 7460 19380 7491
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 18288 7432 19380 7460
rect 18288 7420 18294 7432
rect 12437 7395 12495 7401
rect 12437 7361 12449 7395
rect 12483 7392 12495 7395
rect 12897 7395 12955 7401
rect 12897 7392 12909 7395
rect 12483 7364 12909 7392
rect 12483 7361 12495 7364
rect 12437 7355 12495 7361
rect 12897 7361 12909 7364
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 13817 7395 13875 7401
rect 13817 7361 13829 7395
rect 13863 7392 13875 7395
rect 13863 7364 14044 7392
rect 13863 7361 13875 7364
rect 13817 7355 13875 7361
rect 11103 7296 11652 7324
rect 11103 7293 11115 7296
rect 11057 7287 11115 7293
rect 11698 7284 11704 7336
rect 11756 7324 11762 7336
rect 12529 7327 12587 7333
rect 12529 7324 12541 7327
rect 11756 7296 12541 7324
rect 11756 7284 11762 7296
rect 12529 7293 12541 7296
rect 12575 7293 12587 7327
rect 12710 7324 12716 7336
rect 12671 7296 12716 7324
rect 12529 7287 12587 7293
rect 12710 7284 12716 7296
rect 12768 7284 12774 7336
rect 13909 7327 13967 7333
rect 13909 7293 13921 7327
rect 13955 7293 13967 7327
rect 13909 7287 13967 7293
rect 8588 7228 13768 7256
rect 6457 7219 6515 7225
rect 9125 7191 9183 7197
rect 9125 7188 9137 7191
rect 5920 7160 9137 7188
rect 9125 7157 9137 7160
rect 9171 7157 9183 7191
rect 9125 7151 9183 7157
rect 9858 7148 9864 7200
rect 9916 7188 9922 7200
rect 10045 7191 10103 7197
rect 10045 7188 10057 7191
rect 9916 7160 10057 7188
rect 9916 7148 9922 7160
rect 10045 7157 10057 7160
rect 10091 7188 10103 7191
rect 10594 7188 10600 7200
rect 10091 7160 10600 7188
rect 10091 7157 10103 7160
rect 10045 7151 10103 7157
rect 10594 7148 10600 7160
rect 10652 7148 10658 7200
rect 11698 7148 11704 7200
rect 11756 7188 11762 7200
rect 11885 7191 11943 7197
rect 11885 7188 11897 7191
rect 11756 7160 11897 7188
rect 11756 7148 11762 7160
rect 11885 7157 11897 7160
rect 11931 7157 11943 7191
rect 11885 7151 11943 7157
rect 12158 7148 12164 7200
rect 12216 7188 12222 7200
rect 12434 7188 12440 7200
rect 12216 7160 12440 7188
rect 12216 7148 12222 7160
rect 12434 7148 12440 7160
rect 12492 7148 12498 7200
rect 13740 7188 13768 7228
rect 13814 7216 13820 7268
rect 13872 7256 13878 7268
rect 13924 7256 13952 7287
rect 13872 7228 13952 7256
rect 14016 7256 14044 7364
rect 14734 7352 14740 7404
rect 14792 7392 14798 7404
rect 14792 7364 14964 7392
rect 14792 7352 14798 7364
rect 14936 7336 14964 7364
rect 15194 7352 15200 7404
rect 15252 7392 15258 7404
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 15252 7364 15485 7392
rect 15252 7352 15258 7364
rect 15473 7361 15485 7364
rect 15519 7361 15531 7395
rect 20438 7392 20444 7404
rect 20496 7401 20502 7404
rect 15473 7355 15531 7361
rect 15764 7364 20444 7392
rect 14093 7327 14151 7333
rect 14093 7293 14105 7327
rect 14139 7324 14151 7327
rect 14918 7324 14924 7336
rect 14139 7296 14780 7324
rect 14879 7296 14924 7324
rect 14139 7293 14151 7296
rect 14093 7287 14151 7293
rect 14277 7259 14335 7265
rect 14277 7256 14289 7259
rect 14016 7228 14289 7256
rect 13872 7216 13878 7228
rect 14277 7225 14289 7228
rect 14323 7225 14335 7259
rect 14752 7256 14780 7296
rect 14918 7284 14924 7296
rect 14976 7284 14982 7336
rect 15764 7333 15792 7364
rect 20438 7352 20444 7364
rect 20496 7355 20508 7401
rect 20717 7395 20775 7401
rect 20717 7361 20729 7395
rect 20763 7392 20775 7395
rect 20824 7392 20852 7488
rect 20763 7364 20852 7392
rect 20763 7361 20775 7364
rect 20717 7355 20775 7361
rect 20496 7352 20502 7355
rect 15749 7327 15807 7333
rect 15749 7293 15761 7327
rect 15795 7293 15807 7327
rect 15749 7287 15807 7293
rect 19518 7256 19524 7268
rect 14752 7228 19524 7256
rect 14277 7219 14335 7225
rect 19518 7216 19524 7228
rect 19576 7216 19582 7268
rect 15105 7191 15163 7197
rect 15105 7188 15117 7191
rect 13740 7160 15117 7188
rect 15105 7157 15117 7160
rect 15151 7157 15163 7191
rect 15105 7151 15163 7157
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 1394 6944 1400 6996
rect 1452 6984 1458 6996
rect 1949 6987 2007 6993
rect 1949 6984 1961 6987
rect 1452 6956 1961 6984
rect 1452 6944 1458 6956
rect 1949 6953 1961 6956
rect 1995 6953 2007 6987
rect 1949 6947 2007 6953
rect 5810 6944 5816 6996
rect 5868 6984 5874 6996
rect 6457 6987 6515 6993
rect 6457 6984 6469 6987
rect 5868 6956 6469 6984
rect 5868 6944 5874 6956
rect 6457 6953 6469 6956
rect 6503 6953 6515 6987
rect 6457 6947 6515 6953
rect 7190 6944 7196 6996
rect 7248 6984 7254 6996
rect 7285 6987 7343 6993
rect 7285 6984 7297 6987
rect 7248 6956 7297 6984
rect 7248 6944 7254 6956
rect 7285 6953 7297 6956
rect 7331 6953 7343 6987
rect 8386 6984 8392 6996
rect 8347 6956 8392 6984
rect 7285 6947 7343 6953
rect 8386 6944 8392 6956
rect 8444 6944 8450 6996
rect 9306 6984 9312 6996
rect 9267 6956 9312 6984
rect 9306 6944 9312 6956
rect 9364 6944 9370 6996
rect 9950 6984 9956 6996
rect 9600 6956 9956 6984
rect 1581 6919 1639 6925
rect 1581 6885 1593 6919
rect 1627 6914 1639 6919
rect 7208 6916 7236 6944
rect 1627 6886 1661 6914
rect 7208 6888 8064 6916
rect 1627 6885 1639 6886
rect 1581 6879 1639 6885
rect 1596 6848 1624 6879
rect 4062 6848 4068 6860
rect 1596 6820 2774 6848
rect 4023 6820 4068 6848
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 1670 6780 1676 6792
rect 1631 6752 1676 6780
rect 1670 6740 1676 6752
rect 1728 6780 1734 6792
rect 2133 6783 2191 6789
rect 2133 6780 2145 6783
rect 1728 6752 2145 6780
rect 1728 6740 1734 6752
rect 2133 6749 2145 6752
rect 2179 6749 2191 6783
rect 2746 6780 2774 6820
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 4157 6851 4215 6857
rect 4157 6817 4169 6851
rect 4203 6848 4215 6851
rect 4798 6848 4804 6860
rect 4203 6820 4804 6848
rect 4203 6817 4215 6820
rect 4157 6811 4215 6817
rect 4172 6780 4200 6811
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 4890 6808 4896 6860
rect 4948 6848 4954 6860
rect 4948 6820 6960 6848
rect 4948 6808 4954 6820
rect 2746 6752 4200 6780
rect 4249 6783 4307 6789
rect 2133 6743 2191 6749
rect 4249 6749 4261 6783
rect 4295 6780 4307 6783
rect 4430 6780 4436 6792
rect 4295 6752 4436 6780
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 4430 6740 4436 6752
rect 4488 6740 4494 6792
rect 5718 6740 5724 6792
rect 5776 6780 5782 6792
rect 5994 6780 6000 6792
rect 5776 6752 6000 6780
rect 5776 6740 5782 6752
rect 5994 6740 6000 6752
rect 6052 6780 6058 6792
rect 6089 6783 6147 6789
rect 6089 6780 6101 6783
rect 6052 6752 6101 6780
rect 6052 6740 6058 6752
rect 6089 6749 6101 6752
rect 6135 6780 6147 6783
rect 6638 6780 6644 6792
rect 6135 6752 6644 6780
rect 6135 6749 6147 6752
rect 6089 6743 6147 6749
rect 6638 6740 6644 6752
rect 6696 6740 6702 6792
rect 6822 6780 6828 6792
rect 6783 6752 6828 6780
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 6932 6780 6960 6820
rect 7098 6808 7104 6860
rect 7156 6848 7162 6860
rect 7208 6848 7236 6888
rect 7837 6851 7895 6857
rect 7156 6820 7249 6848
rect 7156 6808 7162 6820
rect 7837 6817 7849 6851
rect 7883 6848 7895 6851
rect 7926 6848 7932 6860
rect 7883 6820 7932 6848
rect 7883 6817 7895 6820
rect 7837 6811 7895 6817
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 8036 6848 8064 6888
rect 8202 6876 8208 6928
rect 8260 6916 8266 6928
rect 9600 6916 9628 6956
rect 9950 6944 9956 6956
rect 10008 6944 10014 6996
rect 10137 6987 10195 6993
rect 10137 6953 10149 6987
rect 10183 6984 10195 6987
rect 10226 6984 10232 6996
rect 10183 6956 10232 6984
rect 10183 6953 10195 6956
rect 10137 6947 10195 6953
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 10410 6944 10416 6996
rect 10468 6984 10474 6996
rect 12066 6984 12072 6996
rect 10468 6956 12072 6984
rect 10468 6944 10474 6956
rect 12066 6944 12072 6956
rect 12124 6944 12130 6996
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 14093 6987 14151 6993
rect 14093 6984 14105 6987
rect 13872 6956 14105 6984
rect 13872 6944 13878 6956
rect 14093 6953 14105 6956
rect 14139 6953 14151 6987
rect 14093 6947 14151 6953
rect 8260 6888 9628 6916
rect 8260 6876 8266 6888
rect 9674 6876 9680 6928
rect 9732 6916 9738 6928
rect 9732 6888 9904 6916
rect 9732 6876 9738 6888
rect 8941 6851 8999 6857
rect 8941 6848 8953 6851
rect 8036 6820 8953 6848
rect 8941 6817 8953 6820
rect 8987 6817 8999 6851
rect 9214 6848 9220 6860
rect 9175 6820 9220 6848
rect 8941 6811 8999 6817
rect 9214 6808 9220 6820
rect 9272 6848 9278 6860
rect 9876 6857 9904 6888
rect 10612 6888 10916 6916
rect 9769 6851 9827 6857
rect 9769 6848 9781 6851
rect 9272 6820 9781 6848
rect 9272 6808 9278 6820
rect 9769 6817 9781 6820
rect 9815 6817 9827 6851
rect 9769 6811 9827 6817
rect 9861 6851 9919 6857
rect 9861 6817 9873 6851
rect 9907 6817 9919 6851
rect 9861 6811 9919 6817
rect 10318 6808 10324 6860
rect 10376 6848 10382 6860
rect 10612 6848 10640 6888
rect 10778 6848 10784 6860
rect 10376 6820 10640 6848
rect 10739 6820 10784 6848
rect 10376 6808 10382 6820
rect 10778 6808 10784 6820
rect 10836 6808 10842 6860
rect 10888 6848 10916 6888
rect 13998 6876 14004 6928
rect 14056 6916 14062 6928
rect 17770 6916 17776 6928
rect 14056 6888 17776 6916
rect 14056 6876 14062 6888
rect 17770 6876 17776 6888
rect 17828 6876 17834 6928
rect 11698 6848 11704 6860
rect 10888 6820 11704 6848
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 11977 6851 12035 6857
rect 11977 6817 11989 6851
rect 12023 6848 12035 6851
rect 12710 6848 12716 6860
rect 12023 6820 12716 6848
rect 12023 6817 12035 6820
rect 11977 6811 12035 6817
rect 12710 6808 12716 6820
rect 12768 6808 12774 6860
rect 14734 6848 14740 6860
rect 14695 6820 14740 6848
rect 14734 6808 14740 6820
rect 14792 6808 14798 6860
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 6932 6752 8033 6780
rect 8021 6749 8033 6752
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 10962 6780 10968 6792
rect 9732 6752 10968 6780
rect 9732 6740 9738 6752
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6780 14611 6783
rect 17862 6780 17868 6792
rect 14599 6752 17868 6780
rect 14599 6749 14611 6752
rect 14553 6743 14611 6749
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 1412 6712 1440 6740
rect 2317 6715 2375 6721
rect 2317 6712 2329 6715
rect 1412 6684 2329 6712
rect 2317 6681 2329 6684
rect 2363 6681 2375 6715
rect 9950 6712 9956 6724
rect 2317 6675 2375 6681
rect 4632 6684 9956 6712
rect 1857 6647 1915 6653
rect 1857 6613 1869 6647
rect 1903 6644 1915 6647
rect 2498 6644 2504 6656
rect 1903 6616 2504 6644
rect 1903 6613 1915 6616
rect 1857 6607 1915 6613
rect 2498 6604 2504 6616
rect 2556 6644 2562 6656
rect 3970 6644 3976 6656
rect 2556 6616 3976 6644
rect 2556 6604 2562 6616
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 4632 6653 4660 6684
rect 9950 6672 9956 6684
rect 10008 6672 10014 6724
rect 10502 6712 10508 6724
rect 10463 6684 10508 6712
rect 10502 6672 10508 6684
rect 10560 6672 10566 6724
rect 12069 6715 12127 6721
rect 12069 6681 12081 6715
rect 12115 6712 12127 6715
rect 16022 6712 16028 6724
rect 12115 6684 16028 6712
rect 12115 6681 12127 6684
rect 12069 6675 12127 6681
rect 16022 6672 16028 6684
rect 16080 6672 16086 6724
rect 4617 6647 4675 6653
rect 4617 6613 4629 6647
rect 4663 6613 4675 6647
rect 4617 6607 4675 6613
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 4764 6616 4809 6644
rect 4764 6604 4770 6616
rect 4982 6604 4988 6656
rect 5040 6644 5046 6656
rect 5445 6647 5503 6653
rect 5445 6644 5457 6647
rect 5040 6616 5457 6644
rect 5040 6604 5046 6616
rect 5445 6613 5457 6616
rect 5491 6613 5503 6647
rect 5445 6607 5503 6613
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 6270 6644 6276 6656
rect 5592 6616 6276 6644
rect 5592 6604 5598 6616
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 6638 6604 6644 6656
rect 6696 6644 6702 6656
rect 6917 6647 6975 6653
rect 6917 6644 6929 6647
rect 6696 6616 6929 6644
rect 6696 6604 6702 6616
rect 6917 6613 6929 6616
rect 6963 6613 6975 6647
rect 6917 6607 6975 6613
rect 7561 6647 7619 6653
rect 7561 6613 7573 6647
rect 7607 6644 7619 6647
rect 7926 6644 7932 6656
rect 7607 6616 7932 6644
rect 7607 6613 7619 6616
rect 7561 6607 7619 6613
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 8386 6604 8392 6656
rect 8444 6644 8450 6656
rect 8573 6647 8631 6653
rect 8573 6644 8585 6647
rect 8444 6616 8585 6644
rect 8444 6604 8450 6616
rect 8573 6613 8585 6616
rect 8619 6644 8631 6647
rect 9030 6644 9036 6656
rect 8619 6616 9036 6644
rect 8619 6613 8631 6616
rect 8573 6607 8631 6613
rect 9030 6604 9036 6616
rect 9088 6644 9094 6656
rect 9582 6644 9588 6656
rect 9088 6616 9588 6644
rect 9088 6604 9094 6616
rect 9582 6604 9588 6616
rect 9640 6604 9646 6656
rect 10594 6644 10600 6656
rect 10555 6616 10600 6644
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 12161 6647 12219 6653
rect 12161 6644 12173 6647
rect 11204 6616 12173 6644
rect 11204 6604 11210 6616
rect 12161 6613 12173 6616
rect 12207 6613 12219 6647
rect 12161 6607 12219 6613
rect 12434 6604 12440 6656
rect 12492 6644 12498 6656
rect 12529 6647 12587 6653
rect 12529 6644 12541 6647
rect 12492 6616 12541 6644
rect 12492 6604 12498 6616
rect 12529 6613 12541 6616
rect 12575 6613 12587 6647
rect 12529 6607 12587 6613
rect 12986 6604 12992 6656
rect 13044 6644 13050 6656
rect 13262 6644 13268 6656
rect 13044 6616 13268 6644
rect 13044 6604 13050 6616
rect 13262 6604 13268 6616
rect 13320 6604 13326 6656
rect 14274 6604 14280 6656
rect 14332 6644 14338 6656
rect 14461 6647 14519 6653
rect 14461 6644 14473 6647
rect 14332 6616 14473 6644
rect 14332 6604 14338 6616
rect 14461 6613 14473 6616
rect 14507 6613 14519 6647
rect 14461 6607 14519 6613
rect 14826 6604 14832 6656
rect 14884 6644 14890 6656
rect 14921 6647 14979 6653
rect 14921 6644 14933 6647
rect 14884 6616 14933 6644
rect 14884 6604 14890 6616
rect 14921 6613 14933 6616
rect 14967 6644 14979 6647
rect 15010 6644 15016 6656
rect 14967 6616 15016 6644
rect 14967 6613 14979 6616
rect 14921 6607 14979 6613
rect 15010 6604 15016 6616
rect 15068 6604 15074 6656
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6409 1639 6443
rect 2038 6440 2044 6452
rect 1999 6412 2044 6440
rect 1581 6403 1639 6409
rect 1596 6372 1624 6403
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 4341 6443 4399 6449
rect 4341 6409 4353 6443
rect 4387 6440 4399 6443
rect 4614 6440 4620 6452
rect 4387 6412 4620 6440
rect 4387 6409 4399 6412
rect 4341 6403 4399 6409
rect 4614 6400 4620 6412
rect 4672 6400 4678 6452
rect 4801 6443 4859 6449
rect 4801 6409 4813 6443
rect 4847 6440 4859 6443
rect 7101 6443 7159 6449
rect 4847 6412 7052 6440
rect 4847 6409 4859 6412
rect 4801 6403 4859 6409
rect 1949 6375 2007 6381
rect 1949 6372 1961 6375
rect 1596 6344 1961 6372
rect 1949 6341 1961 6344
rect 1995 6372 2007 6375
rect 2130 6372 2136 6384
rect 1995 6344 2136 6372
rect 1995 6341 2007 6344
rect 1949 6335 2007 6341
rect 2130 6332 2136 6344
rect 2188 6332 2194 6384
rect 4433 6375 4491 6381
rect 4433 6341 4445 6375
rect 4479 6372 4491 6375
rect 5721 6375 5779 6381
rect 5721 6372 5733 6375
rect 4479 6344 5733 6372
rect 4479 6341 4491 6344
rect 4433 6335 4491 6341
rect 5721 6341 5733 6344
rect 5767 6341 5779 6375
rect 7024 6372 7052 6412
rect 7101 6409 7113 6443
rect 7147 6440 7159 6443
rect 7374 6440 7380 6452
rect 7147 6412 7380 6440
rect 7147 6409 7159 6412
rect 7101 6403 7159 6409
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 7469 6443 7527 6449
rect 7469 6409 7481 6443
rect 7515 6440 7527 6443
rect 7929 6443 7987 6449
rect 7929 6440 7941 6443
rect 7515 6412 7941 6440
rect 7515 6409 7527 6412
rect 7469 6403 7527 6409
rect 7929 6409 7941 6412
rect 7975 6409 7987 6443
rect 7929 6403 7987 6409
rect 8294 6400 8300 6452
rect 8352 6440 8358 6452
rect 8757 6443 8815 6449
rect 8757 6440 8769 6443
rect 8352 6412 8769 6440
rect 8352 6400 8358 6412
rect 8757 6409 8769 6412
rect 8803 6409 8815 6443
rect 8757 6403 8815 6409
rect 9030 6400 9036 6452
rect 9088 6440 9094 6452
rect 9217 6443 9275 6449
rect 9217 6440 9229 6443
rect 9088 6412 9229 6440
rect 9088 6400 9094 6412
rect 9217 6409 9229 6412
rect 9263 6409 9275 6443
rect 9950 6440 9956 6452
rect 9911 6412 9956 6440
rect 9217 6403 9275 6409
rect 9950 6400 9956 6412
rect 10008 6400 10014 6452
rect 10594 6400 10600 6452
rect 10652 6440 10658 6452
rect 12253 6443 12311 6449
rect 12253 6440 12265 6443
rect 10652 6412 12265 6440
rect 10652 6400 10658 6412
rect 12253 6409 12265 6412
rect 12299 6409 12311 6443
rect 15562 6440 15568 6452
rect 12253 6403 12311 6409
rect 12912 6412 15568 6440
rect 10045 6375 10103 6381
rect 10045 6372 10057 6375
rect 7024 6344 10057 6372
rect 5721 6335 5779 6341
rect 10045 6341 10057 6344
rect 10091 6341 10103 6375
rect 10045 6335 10103 6341
rect 1394 6304 1400 6316
rect 1355 6276 1400 6304
rect 1394 6264 1400 6276
rect 1452 6264 1458 6316
rect 5261 6307 5319 6313
rect 2746 6276 5212 6304
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6236 1915 6239
rect 2038 6236 2044 6248
rect 1903 6208 2044 6236
rect 1903 6205 1915 6208
rect 1857 6199 1915 6205
rect 2038 6196 2044 6208
rect 2096 6196 2102 6248
rect 2409 6103 2467 6109
rect 2409 6069 2421 6103
rect 2455 6100 2467 6103
rect 2746 6100 2774 6276
rect 4154 6196 4160 6248
rect 4212 6236 4218 6248
rect 4249 6239 4307 6245
rect 4249 6236 4261 6239
rect 4212 6208 4261 6236
rect 4212 6196 4218 6208
rect 4249 6205 4261 6208
rect 4295 6236 4307 6239
rect 4706 6236 4712 6248
rect 4295 6208 4712 6236
rect 4295 6205 4307 6208
rect 4249 6199 4307 6205
rect 4706 6196 4712 6208
rect 4764 6196 4770 6248
rect 5184 6245 5212 6276
rect 5261 6273 5273 6307
rect 5307 6273 5319 6307
rect 5261 6267 5319 6273
rect 7009 6307 7067 6313
rect 7009 6273 7021 6307
rect 7055 6304 7067 6307
rect 7466 6304 7472 6316
rect 7055 6276 7472 6304
rect 7055 6273 7067 6276
rect 7009 6267 7067 6273
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6205 5135 6239
rect 5077 6199 5135 6205
rect 5169 6239 5227 6245
rect 5169 6205 5181 6239
rect 5215 6205 5227 6239
rect 5169 6199 5227 6205
rect 2455 6072 2774 6100
rect 5092 6100 5120 6199
rect 5276 6180 5304 6267
rect 7466 6264 7472 6276
rect 7524 6304 7530 6316
rect 8294 6304 8300 6316
rect 7524 6276 8156 6304
rect 8255 6276 8300 6304
rect 7524 6264 7530 6276
rect 7190 6196 7196 6248
rect 7248 6236 7254 6248
rect 7561 6239 7619 6245
rect 7561 6236 7573 6239
rect 7248 6208 7573 6236
rect 7248 6196 7254 6208
rect 7561 6205 7573 6208
rect 7607 6205 7619 6239
rect 7561 6199 7619 6205
rect 7745 6239 7803 6245
rect 7745 6205 7757 6239
rect 7791 6236 7803 6239
rect 8018 6236 8024 6248
rect 7791 6208 8024 6236
rect 7791 6205 7803 6208
rect 7745 6199 7803 6205
rect 8018 6196 8024 6208
rect 8076 6196 8082 6248
rect 8128 6236 8156 6276
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 9122 6304 9128 6316
rect 9083 6276 9128 6304
rect 9122 6264 9128 6276
rect 9180 6264 9186 6316
rect 10965 6307 11023 6313
rect 10965 6304 10977 6307
rect 9508 6276 10977 6304
rect 8389 6239 8447 6245
rect 8389 6236 8401 6239
rect 8128 6208 8401 6236
rect 8389 6205 8401 6208
rect 8435 6205 8447 6239
rect 8389 6199 8447 6205
rect 8478 6196 8484 6248
rect 8536 6236 8542 6248
rect 8573 6239 8631 6245
rect 8573 6236 8585 6239
rect 8536 6208 8585 6236
rect 8536 6196 8542 6208
rect 8573 6205 8585 6208
rect 8619 6236 8631 6239
rect 9306 6236 9312 6248
rect 8619 6208 9312 6236
rect 8619 6205 8631 6208
rect 8573 6199 8631 6205
rect 9306 6196 9312 6208
rect 9364 6236 9370 6248
rect 9364 6208 9409 6236
rect 9364 6196 9370 6208
rect 5258 6128 5264 6180
rect 5316 6128 5322 6180
rect 5629 6171 5687 6177
rect 5629 6137 5641 6171
rect 5675 6168 5687 6171
rect 9508 6168 9536 6276
rect 10965 6273 10977 6276
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 11514 6264 11520 6316
rect 11572 6304 11578 6316
rect 12618 6304 12624 6316
rect 11572 6276 12020 6304
rect 12579 6276 12624 6304
rect 11572 6264 11578 6276
rect 9861 6239 9919 6245
rect 9861 6205 9873 6239
rect 9907 6205 9919 6239
rect 10686 6236 10692 6248
rect 10647 6208 10692 6236
rect 9861 6199 9919 6205
rect 5675 6140 9536 6168
rect 9876 6168 9904 6199
rect 10686 6196 10692 6208
rect 10744 6196 10750 6248
rect 10870 6236 10876 6248
rect 10831 6208 10876 6236
rect 10870 6196 10876 6208
rect 10928 6196 10934 6248
rect 11790 6196 11796 6248
rect 11848 6236 11854 6248
rect 11885 6239 11943 6245
rect 11885 6236 11897 6239
rect 11848 6208 11897 6236
rect 11848 6196 11854 6208
rect 11885 6205 11897 6208
rect 11931 6205 11943 6239
rect 11992 6236 12020 6276
rect 12618 6264 12624 6276
rect 12676 6264 12682 6316
rect 12710 6236 12716 6248
rect 11992 6208 12572 6236
rect 12671 6208 12716 6236
rect 11885 6199 11943 6205
rect 11054 6168 11060 6180
rect 9876 6140 11060 6168
rect 5675 6137 5687 6140
rect 5629 6131 5687 6137
rect 11054 6128 11060 6140
rect 11112 6128 11118 6180
rect 12434 6168 12440 6180
rect 11256 6140 12440 6168
rect 8110 6100 8116 6112
rect 5092 6072 8116 6100
rect 2455 6069 2467 6072
rect 2409 6063 2467 6069
rect 8110 6060 8116 6072
rect 8168 6100 8174 6112
rect 10134 6100 10140 6112
rect 8168 6072 10140 6100
rect 8168 6060 8174 6072
rect 10134 6060 10140 6072
rect 10192 6060 10198 6112
rect 10413 6103 10471 6109
rect 10413 6069 10425 6103
rect 10459 6100 10471 6103
rect 11256 6100 11284 6140
rect 12434 6128 12440 6140
rect 12492 6128 12498 6180
rect 12544 6168 12572 6208
rect 12710 6196 12716 6208
rect 12768 6196 12774 6248
rect 12912 6245 12940 6412
rect 15562 6400 15568 6412
rect 15620 6400 15626 6452
rect 21174 6400 21180 6452
rect 21232 6440 21238 6452
rect 21361 6443 21419 6449
rect 21361 6440 21373 6443
rect 21232 6412 21373 6440
rect 21232 6400 21238 6412
rect 21361 6409 21373 6412
rect 21407 6409 21419 6443
rect 21361 6403 21419 6409
rect 13262 6264 13268 6316
rect 13320 6304 13326 6316
rect 14277 6307 14335 6313
rect 13320 6276 14228 6304
rect 13320 6264 13326 6276
rect 12897 6239 12955 6245
rect 12897 6205 12909 6239
rect 12943 6205 12955 6239
rect 13998 6236 14004 6248
rect 13959 6208 14004 6236
rect 12897 6199 12955 6205
rect 13998 6196 14004 6208
rect 14056 6196 14062 6248
rect 14200 6245 14228 6276
rect 14277 6273 14289 6307
rect 14323 6273 14335 6307
rect 14277 6267 14335 6273
rect 21269 6307 21327 6313
rect 21269 6273 21281 6307
rect 21315 6304 21327 6307
rect 21542 6304 21548 6316
rect 21315 6276 21548 6304
rect 21315 6273 21327 6276
rect 21269 6267 21327 6273
rect 14185 6239 14243 6245
rect 14185 6205 14197 6239
rect 14231 6205 14243 6239
rect 14185 6199 14243 6205
rect 12544 6140 12848 6168
rect 10459 6072 11284 6100
rect 11333 6103 11391 6109
rect 10459 6069 10471 6072
rect 10413 6063 10471 6069
rect 11333 6069 11345 6103
rect 11379 6100 11391 6103
rect 11606 6100 11612 6112
rect 11379 6072 11612 6100
rect 11379 6069 11391 6072
rect 11333 6063 11391 6069
rect 11606 6060 11612 6072
rect 11664 6060 11670 6112
rect 11698 6060 11704 6112
rect 11756 6100 11762 6112
rect 12710 6100 12716 6112
rect 11756 6072 12716 6100
rect 11756 6060 11762 6072
rect 12710 6060 12716 6072
rect 12768 6060 12774 6112
rect 12820 6100 12848 6140
rect 13538 6128 13544 6180
rect 13596 6168 13602 6180
rect 14292 6168 14320 6267
rect 21542 6264 21548 6276
rect 21600 6264 21606 6316
rect 15654 6168 15660 6180
rect 13596 6140 14320 6168
rect 14375 6140 15660 6168
rect 13596 6128 13602 6140
rect 14375 6100 14403 6140
rect 15654 6128 15660 6140
rect 15712 6128 15718 6180
rect 12820 6072 14403 6100
rect 14645 6103 14703 6109
rect 14645 6069 14657 6103
rect 14691 6100 14703 6103
rect 15838 6100 15844 6112
rect 14691 6072 15844 6100
rect 14691 6069 14703 6072
rect 14645 6063 14703 6069
rect 15838 6060 15844 6072
rect 15896 6060 15902 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 1394 5856 1400 5908
rect 1452 5896 1458 5908
rect 1949 5899 2007 5905
rect 1949 5896 1961 5899
rect 1452 5868 1961 5896
rect 1452 5856 1458 5868
rect 1949 5865 1961 5868
rect 1995 5865 2007 5899
rect 7190 5896 7196 5908
rect 7151 5868 7196 5896
rect 1949 5859 2007 5865
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 7282 5856 7288 5908
rect 7340 5896 7346 5908
rect 8478 5896 8484 5908
rect 7340 5868 8484 5896
rect 7340 5856 7346 5868
rect 8478 5856 8484 5868
rect 8536 5856 8542 5908
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 8757 5899 8815 5905
rect 8628 5868 8708 5896
rect 8628 5856 8634 5868
rect 1578 5828 1584 5840
rect 1539 5800 1584 5828
rect 1578 5788 1584 5800
rect 1636 5788 1642 5840
rect 1857 5831 1915 5837
rect 1857 5797 1869 5831
rect 1903 5828 1915 5831
rect 1903 5800 2774 5828
rect 1903 5797 1915 5800
rect 1857 5791 1915 5797
rect 2746 5760 2774 5800
rect 5074 5788 5080 5840
rect 5132 5828 5138 5840
rect 8680 5828 8708 5868
rect 8757 5865 8769 5899
rect 8803 5896 8815 5899
rect 10870 5896 10876 5908
rect 8803 5868 10876 5896
rect 8803 5865 8815 5868
rect 8757 5859 8815 5865
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 12894 5896 12900 5908
rect 10980 5868 12900 5896
rect 10980 5828 11008 5868
rect 12894 5856 12900 5868
rect 12952 5856 12958 5908
rect 13262 5896 13268 5908
rect 13223 5868 13268 5896
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 20714 5896 20720 5908
rect 16684 5868 20720 5896
rect 5132 5800 8524 5828
rect 8680 5800 11008 5828
rect 11149 5831 11207 5837
rect 5132 5788 5138 5800
rect 5350 5760 5356 5772
rect 2746 5732 5356 5760
rect 5350 5720 5356 5732
rect 5408 5720 5414 5772
rect 5810 5760 5816 5772
rect 5771 5732 5816 5760
rect 5810 5720 5816 5732
rect 5868 5720 5874 5772
rect 5905 5763 5963 5769
rect 5905 5729 5917 5763
rect 5951 5760 5963 5763
rect 6546 5760 6552 5772
rect 5951 5732 6552 5760
rect 5951 5729 5963 5732
rect 5905 5723 5963 5729
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 6641 5763 6699 5769
rect 6641 5729 6653 5763
rect 6687 5760 6699 5763
rect 7282 5760 7288 5772
rect 6687 5732 7288 5760
rect 6687 5729 6699 5732
rect 6641 5723 6699 5729
rect 7282 5720 7288 5732
rect 7340 5720 7346 5772
rect 8110 5760 8116 5772
rect 8071 5732 8116 5760
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 1394 5692 1400 5704
rect 1355 5664 1400 5692
rect 1394 5652 1400 5664
rect 1452 5652 1458 5704
rect 1670 5692 1676 5704
rect 1631 5664 1676 5692
rect 1670 5652 1676 5664
rect 1728 5692 1734 5704
rect 2501 5695 2559 5701
rect 2501 5692 2513 5695
rect 1728 5664 2513 5692
rect 1728 5652 1734 5664
rect 2501 5661 2513 5664
rect 2547 5661 2559 5695
rect 2501 5655 2559 5661
rect 5166 5652 5172 5704
rect 5224 5692 5230 5704
rect 5828 5692 5856 5720
rect 5224 5664 5856 5692
rect 5997 5695 6055 5701
rect 5224 5652 5230 5664
rect 5997 5661 6009 5695
rect 6043 5692 6055 5695
rect 6730 5692 6736 5704
rect 6043 5664 6736 5692
rect 6043 5661 6055 5664
rect 5997 5655 6055 5661
rect 6730 5652 6736 5664
rect 6788 5652 6794 5704
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 8389 5695 8447 5701
rect 8389 5692 8401 5695
rect 6972 5664 8401 5692
rect 6972 5652 6978 5664
rect 8389 5661 8401 5664
rect 8435 5661 8447 5695
rect 8496 5692 8524 5800
rect 11149 5797 11161 5831
rect 11195 5828 11207 5831
rect 16574 5828 16580 5840
rect 11195 5800 16580 5828
rect 11195 5797 11207 5800
rect 11149 5791 11207 5797
rect 16574 5788 16580 5800
rect 16632 5788 16638 5840
rect 8846 5720 8852 5772
rect 8904 5760 8910 5772
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 8904 5732 9689 5760
rect 8904 5720 8910 5732
rect 9677 5729 9689 5732
rect 9723 5760 9735 5763
rect 10410 5760 10416 5772
rect 9723 5732 10416 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 10410 5720 10416 5732
rect 10468 5720 10474 5772
rect 10597 5763 10655 5769
rect 10597 5729 10609 5763
rect 10643 5760 10655 5763
rect 11514 5760 11520 5772
rect 10643 5732 11520 5760
rect 10643 5729 10655 5732
rect 10597 5723 10655 5729
rect 11514 5720 11520 5732
rect 11572 5720 11578 5772
rect 11606 5720 11612 5772
rect 11664 5760 11670 5772
rect 12713 5763 12771 5769
rect 11664 5732 12434 5760
rect 11664 5720 11670 5732
rect 10781 5695 10839 5701
rect 10781 5692 10793 5695
rect 8496 5664 10793 5692
rect 8389 5655 8447 5661
rect 10781 5661 10793 5664
rect 10827 5661 10839 5695
rect 11790 5692 11796 5704
rect 11751 5664 11796 5692
rect 10781 5655 10839 5661
rect 11790 5652 11796 5664
rect 11848 5652 11854 5704
rect 12406 5692 12434 5732
rect 12713 5729 12725 5763
rect 12759 5760 12771 5763
rect 13078 5760 13084 5772
rect 12759 5732 13084 5760
rect 12759 5729 12771 5732
rect 12713 5723 12771 5729
rect 13078 5720 13084 5732
rect 13136 5720 13142 5772
rect 13262 5720 13268 5772
rect 13320 5760 13326 5772
rect 13630 5760 13636 5772
rect 13320 5732 13636 5760
rect 13320 5720 13326 5732
rect 13630 5720 13636 5732
rect 13688 5720 13694 5772
rect 16684 5769 16712 5868
rect 20714 5856 20720 5868
rect 20772 5856 20778 5908
rect 17313 5831 17371 5837
rect 17313 5797 17325 5831
rect 17359 5828 17371 5831
rect 18782 5828 18788 5840
rect 17359 5800 18788 5828
rect 17359 5797 17371 5800
rect 17313 5791 17371 5797
rect 18782 5788 18788 5800
rect 18840 5788 18846 5840
rect 16669 5763 16727 5769
rect 16669 5729 16681 5763
rect 16715 5729 16727 5763
rect 17586 5760 17592 5772
rect 17547 5732 17592 5760
rect 16669 5723 16727 5729
rect 17586 5720 17592 5732
rect 17644 5720 17650 5772
rect 20070 5760 20076 5772
rect 20031 5732 20076 5760
rect 20070 5720 20076 5732
rect 20128 5720 20134 5772
rect 13357 5695 13415 5701
rect 13357 5692 13369 5695
rect 12406 5664 13369 5692
rect 13357 5661 13369 5664
rect 13403 5661 13415 5695
rect 13357 5655 13415 5661
rect 16482 5652 16488 5704
rect 16540 5692 16546 5704
rect 17681 5695 17739 5701
rect 17681 5692 17693 5695
rect 16540 5664 17693 5692
rect 16540 5652 16546 5664
rect 17681 5661 17693 5664
rect 17727 5661 17739 5695
rect 17681 5655 17739 5661
rect 1412 5624 1440 5652
rect 2685 5627 2743 5633
rect 2685 5624 2697 5627
rect 1412 5596 2697 5624
rect 2685 5593 2697 5596
rect 2731 5593 2743 5627
rect 2685 5587 2743 5593
rect 4798 5584 4804 5636
rect 4856 5624 4862 5636
rect 6825 5627 6883 5633
rect 6825 5624 6837 5627
rect 4856 5596 6837 5624
rect 4856 5584 4862 5596
rect 6825 5593 6837 5596
rect 6871 5593 6883 5627
rect 6825 5587 6883 5593
rect 8297 5627 8355 5633
rect 8297 5593 8309 5627
rect 8343 5624 8355 5627
rect 9493 5627 9551 5633
rect 8343 5596 9168 5624
rect 8343 5593 8355 5596
rect 8297 5587 8355 5593
rect 2222 5556 2228 5568
rect 2183 5528 2228 5556
rect 2222 5516 2228 5528
rect 2280 5516 2286 5568
rect 4706 5516 4712 5568
rect 4764 5556 4770 5568
rect 4893 5559 4951 5565
rect 4893 5556 4905 5559
rect 4764 5528 4905 5556
rect 4764 5516 4770 5528
rect 4893 5525 4905 5528
rect 4939 5525 4951 5559
rect 4893 5519 4951 5525
rect 4982 5516 4988 5568
rect 5040 5556 5046 5568
rect 5261 5559 5319 5565
rect 5261 5556 5273 5559
rect 5040 5528 5273 5556
rect 5040 5516 5046 5528
rect 5261 5525 5273 5528
rect 5307 5556 5319 5559
rect 5718 5556 5724 5568
rect 5307 5528 5724 5556
rect 5307 5525 5319 5528
rect 5261 5519 5319 5525
rect 5718 5516 5724 5528
rect 5776 5516 5782 5568
rect 6365 5559 6423 5565
rect 6365 5525 6377 5559
rect 6411 5556 6423 5559
rect 6638 5556 6644 5568
rect 6411 5528 6644 5556
rect 6411 5525 6423 5528
rect 6365 5519 6423 5525
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 6733 5559 6791 5565
rect 6733 5525 6745 5559
rect 6779 5556 6791 5559
rect 7006 5556 7012 5568
rect 6779 5528 7012 5556
rect 6779 5525 6791 5528
rect 6733 5519 6791 5525
rect 7006 5516 7012 5528
rect 7064 5556 7070 5568
rect 7285 5559 7343 5565
rect 7285 5556 7297 5559
rect 7064 5528 7297 5556
rect 7064 5516 7070 5528
rect 7285 5525 7297 5528
rect 7331 5556 7343 5559
rect 7374 5556 7380 5568
rect 7331 5528 7380 5556
rect 7331 5525 7343 5528
rect 7285 5519 7343 5525
rect 7374 5516 7380 5528
rect 7432 5516 7438 5568
rect 7926 5556 7932 5568
rect 7887 5528 7932 5556
rect 7926 5516 7932 5528
rect 7984 5516 7990 5568
rect 8754 5516 8760 5568
rect 8812 5556 8818 5568
rect 8941 5559 8999 5565
rect 8941 5556 8953 5559
rect 8812 5528 8953 5556
rect 8812 5516 8818 5528
rect 8941 5525 8953 5528
rect 8987 5556 8999 5559
rect 9030 5556 9036 5568
rect 8987 5528 9036 5556
rect 8987 5525 8999 5528
rect 8941 5519 8999 5525
rect 9030 5516 9036 5528
rect 9088 5516 9094 5568
rect 9140 5565 9168 5596
rect 9493 5593 9505 5627
rect 9539 5624 9551 5627
rect 9766 5624 9772 5636
rect 9539 5596 9772 5624
rect 9539 5593 9551 5596
rect 9493 5587 9551 5593
rect 9766 5584 9772 5596
rect 9824 5584 9830 5636
rect 10870 5584 10876 5636
rect 10928 5624 10934 5636
rect 16945 5627 17003 5633
rect 16945 5624 16957 5627
rect 10928 5596 11744 5624
rect 10928 5584 10934 5596
rect 9125 5559 9183 5565
rect 9125 5525 9137 5559
rect 9171 5525 9183 5559
rect 9125 5519 9183 5525
rect 9582 5516 9588 5568
rect 9640 5556 9646 5568
rect 10686 5556 10692 5568
rect 9640 5528 9685 5556
rect 10647 5528 10692 5556
rect 9640 5516 9646 5528
rect 10686 5516 10692 5528
rect 10744 5516 10750 5568
rect 11054 5516 11060 5568
rect 11112 5556 11118 5568
rect 11330 5556 11336 5568
rect 11112 5528 11336 5556
rect 11112 5516 11118 5528
rect 11330 5516 11336 5528
rect 11388 5516 11394 5568
rect 11716 5565 11744 5596
rect 12406 5596 16957 5624
rect 11701 5559 11759 5565
rect 11701 5525 11713 5559
rect 11747 5525 11759 5559
rect 11701 5519 11759 5525
rect 12161 5559 12219 5565
rect 12161 5525 12173 5559
rect 12207 5556 12219 5559
rect 12406 5556 12434 5596
rect 16945 5593 16957 5596
rect 16991 5593 17003 5627
rect 20349 5627 20407 5633
rect 20349 5624 20361 5627
rect 16945 5587 17003 5593
rect 18156 5596 20361 5624
rect 12802 5556 12808 5568
rect 12207 5528 12434 5556
rect 12763 5528 12808 5556
rect 12207 5525 12219 5528
rect 12161 5519 12219 5525
rect 12802 5516 12808 5528
rect 12860 5516 12866 5568
rect 12894 5516 12900 5568
rect 12952 5556 12958 5568
rect 13538 5556 13544 5568
rect 12952 5528 12997 5556
rect 13499 5528 13544 5556
rect 12952 5516 12958 5528
rect 13538 5516 13544 5528
rect 13596 5516 13602 5568
rect 16574 5516 16580 5568
rect 16632 5556 16638 5568
rect 16853 5559 16911 5565
rect 16853 5556 16865 5559
rect 16632 5528 16865 5556
rect 16632 5516 16638 5528
rect 16853 5525 16865 5528
rect 16899 5525 16911 5559
rect 16853 5519 16911 5525
rect 17770 5516 17776 5568
rect 17828 5556 17834 5568
rect 18156 5565 18184 5596
rect 20349 5593 20361 5596
rect 20395 5593 20407 5627
rect 20349 5587 20407 5593
rect 18141 5559 18199 5565
rect 17828 5528 17873 5556
rect 17828 5516 17834 5528
rect 18141 5525 18153 5559
rect 18187 5525 18199 5559
rect 20254 5556 20260 5568
rect 20215 5528 20260 5556
rect 18141 5519 18199 5525
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 20717 5559 20775 5565
rect 20717 5525 20729 5559
rect 20763 5556 20775 5559
rect 20806 5556 20812 5568
rect 20763 5528 20812 5556
rect 20763 5525 20775 5528
rect 20717 5519 20775 5525
rect 20806 5516 20812 5528
rect 20864 5516 20870 5568
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 2222 5352 2228 5364
rect 2183 5324 2228 5352
rect 2222 5312 2228 5324
rect 2280 5312 2286 5364
rect 2593 5355 2651 5361
rect 2593 5321 2605 5355
rect 2639 5352 2651 5355
rect 5258 5352 5264 5364
rect 2639 5324 5264 5352
rect 2639 5321 2651 5324
rect 2593 5315 2651 5321
rect 5258 5312 5264 5324
rect 5316 5312 5322 5364
rect 6638 5352 6644 5364
rect 6599 5324 6644 5352
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 7101 5355 7159 5361
rect 7101 5321 7113 5355
rect 7147 5321 7159 5355
rect 7101 5315 7159 5321
rect 2133 5287 2191 5293
rect 2133 5253 2145 5287
rect 2179 5284 2191 5287
rect 2314 5284 2320 5296
rect 2179 5256 2320 5284
rect 2179 5253 2191 5256
rect 2133 5247 2191 5253
rect 2314 5244 2320 5256
rect 2372 5244 2378 5296
rect 4614 5284 4620 5296
rect 4527 5256 4620 5284
rect 4614 5244 4620 5256
rect 4672 5284 4678 5296
rect 5537 5287 5595 5293
rect 5537 5284 5549 5287
rect 4672 5256 5549 5284
rect 4672 5244 4678 5256
rect 5537 5253 5549 5256
rect 5583 5253 5595 5287
rect 5537 5247 5595 5253
rect 5718 5244 5724 5296
rect 5776 5284 5782 5296
rect 7116 5284 7144 5315
rect 7926 5312 7932 5364
rect 7984 5352 7990 5364
rect 8297 5355 8355 5361
rect 8297 5352 8309 5355
rect 7984 5324 8309 5352
rect 7984 5312 7990 5324
rect 8297 5321 8309 5324
rect 8343 5321 8355 5355
rect 9306 5352 9312 5364
rect 9267 5324 9312 5352
rect 8297 5315 8355 5321
rect 9306 5312 9312 5324
rect 9364 5352 9370 5364
rect 9674 5352 9680 5364
rect 9364 5324 9680 5352
rect 9364 5312 9370 5324
rect 9674 5312 9680 5324
rect 9732 5352 9738 5364
rect 10137 5355 10195 5361
rect 9732 5324 9777 5352
rect 9732 5312 9738 5324
rect 10137 5321 10149 5355
rect 10183 5352 10195 5355
rect 10686 5352 10692 5364
rect 10183 5324 10692 5352
rect 10183 5321 10195 5324
rect 10137 5315 10195 5321
rect 10686 5312 10692 5324
rect 10744 5312 10750 5364
rect 10965 5355 11023 5361
rect 10965 5321 10977 5355
rect 11011 5352 11023 5355
rect 11885 5355 11943 5361
rect 11885 5352 11897 5355
rect 11011 5324 11897 5352
rect 11011 5321 11023 5324
rect 10965 5315 11023 5321
rect 11885 5321 11897 5324
rect 11931 5321 11943 5355
rect 11885 5315 11943 5321
rect 12802 5312 12808 5364
rect 12860 5352 12866 5364
rect 13173 5355 13231 5361
rect 13173 5352 13185 5355
rect 12860 5324 13185 5352
rect 12860 5312 12866 5324
rect 13173 5321 13185 5324
rect 13219 5321 13231 5355
rect 13173 5315 13231 5321
rect 13354 5312 13360 5364
rect 13412 5352 13418 5364
rect 13541 5355 13599 5361
rect 13541 5352 13553 5355
rect 13412 5324 13553 5352
rect 13412 5312 13418 5324
rect 13541 5321 13553 5324
rect 13587 5321 13599 5355
rect 13541 5315 13599 5321
rect 17221 5355 17279 5361
rect 17221 5321 17233 5355
rect 17267 5352 17279 5355
rect 17770 5352 17776 5364
rect 17267 5324 17776 5352
rect 17267 5321 17279 5324
rect 17221 5315 17279 5321
rect 17770 5312 17776 5324
rect 17828 5312 17834 5364
rect 11977 5287 12035 5293
rect 11977 5284 11989 5287
rect 5776 5256 6868 5284
rect 7116 5256 11989 5284
rect 5776 5244 5782 5256
rect 1486 5216 1492 5228
rect 1447 5188 1492 5216
rect 1486 5176 1492 5188
rect 1544 5216 1550 5228
rect 2685 5219 2743 5225
rect 2685 5216 2697 5219
rect 1544 5188 2697 5216
rect 1544 5176 1550 5188
rect 2685 5185 2697 5188
rect 2731 5185 2743 5219
rect 2685 5179 2743 5185
rect 4709 5219 4767 5225
rect 4709 5185 4721 5219
rect 4755 5216 4767 5219
rect 5350 5216 5356 5228
rect 4755 5188 5356 5216
rect 4755 5185 4767 5188
rect 4709 5179 4767 5185
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 5810 5176 5816 5228
rect 5868 5216 5874 5228
rect 6733 5219 6791 5225
rect 6733 5216 6745 5219
rect 5868 5188 6745 5216
rect 5868 5176 5874 5188
rect 6733 5185 6745 5188
rect 6779 5185 6791 5219
rect 6840 5216 6868 5256
rect 11977 5253 11989 5256
rect 12023 5253 12035 5287
rect 11977 5247 12035 5253
rect 12066 5244 12072 5296
rect 12124 5284 12130 5296
rect 15381 5287 15439 5293
rect 15381 5284 15393 5287
rect 12124 5256 15393 5284
rect 12124 5244 12130 5256
rect 15381 5253 15393 5256
rect 15427 5253 15439 5287
rect 15381 5247 15439 5253
rect 6840 5188 8708 5216
rect 6733 5179 6791 5185
rect 2038 5148 2044 5160
rect 1999 5120 2044 5148
rect 2038 5108 2044 5120
rect 2096 5108 2102 5160
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5148 4583 5151
rect 4982 5148 4988 5160
rect 4571 5120 4988 5148
rect 4571 5117 4583 5120
rect 4525 5111 4583 5117
rect 4982 5108 4988 5120
rect 5040 5108 5046 5160
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5117 5319 5151
rect 5261 5111 5319 5117
rect 5445 5151 5503 5157
rect 5445 5117 5457 5151
rect 5491 5148 5503 5151
rect 5718 5148 5724 5160
rect 5491 5120 5724 5148
rect 5491 5117 5503 5120
rect 5445 5111 5503 5117
rect 1673 5083 1731 5089
rect 1673 5049 1685 5083
rect 1719 5080 1731 5083
rect 4706 5080 4712 5092
rect 1719 5052 4712 5080
rect 1719 5049 1731 5052
rect 1673 5043 1731 5049
rect 4706 5040 4712 5052
rect 4764 5040 4770 5092
rect 5074 5080 5080 5092
rect 5035 5052 5080 5080
rect 5074 5040 5080 5052
rect 5132 5040 5138 5092
rect 2038 4972 2044 5024
rect 2096 5012 2102 5024
rect 5276 5012 5304 5111
rect 5718 5108 5724 5120
rect 5776 5108 5782 5160
rect 5994 5148 6000 5160
rect 5955 5120 6000 5148
rect 5994 5108 6000 5120
rect 6052 5108 6058 5160
rect 6546 5148 6552 5160
rect 6507 5120 6552 5148
rect 6546 5108 6552 5120
rect 6604 5108 6610 5160
rect 8389 5151 8447 5157
rect 8389 5117 8401 5151
rect 8435 5117 8447 5151
rect 8389 5111 8447 5117
rect 5905 5083 5963 5089
rect 5905 5049 5917 5083
rect 5951 5080 5963 5083
rect 6914 5080 6920 5092
rect 5951 5052 6920 5080
rect 5951 5049 5963 5052
rect 5905 5043 5963 5049
rect 6914 5040 6920 5052
rect 6972 5040 6978 5092
rect 7834 5040 7840 5092
rect 7892 5080 7898 5092
rect 7929 5083 7987 5089
rect 7929 5080 7941 5083
rect 7892 5052 7941 5080
rect 7892 5040 7898 5052
rect 7929 5049 7941 5052
rect 7975 5049 7987 5083
rect 7929 5043 7987 5049
rect 7006 5012 7012 5024
rect 2096 4984 7012 5012
rect 2096 4972 2102 4984
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 7190 4972 7196 5024
rect 7248 5012 7254 5024
rect 7745 5015 7803 5021
rect 7745 5012 7757 5015
rect 7248 4984 7757 5012
rect 7248 4972 7254 4984
rect 7745 4981 7757 4984
rect 7791 5012 7803 5015
rect 8404 5012 8432 5111
rect 8478 5108 8484 5160
rect 8536 5148 8542 5160
rect 8680 5148 8708 5188
rect 9398 5176 9404 5228
rect 9456 5216 9462 5228
rect 9769 5219 9827 5225
rect 9769 5216 9781 5219
rect 9456 5188 9781 5216
rect 9456 5176 9462 5188
rect 9769 5185 9781 5188
rect 9815 5185 9827 5219
rect 10597 5219 10655 5225
rect 10597 5216 10609 5219
rect 9769 5179 9827 5185
rect 9876 5188 10609 5216
rect 9490 5148 9496 5160
rect 8536 5120 8581 5148
rect 8680 5120 9496 5148
rect 8536 5108 8542 5120
rect 9490 5108 9496 5120
rect 9548 5108 9554 5160
rect 9876 5148 9904 5188
rect 10597 5185 10609 5188
rect 10643 5185 10655 5219
rect 10597 5179 10655 5185
rect 10870 5176 10876 5228
rect 10928 5216 10934 5228
rect 10928 5188 12572 5216
rect 10928 5176 10934 5188
rect 12544 5160 12572 5188
rect 12618 5176 12624 5228
rect 12676 5216 12682 5228
rect 12805 5219 12863 5225
rect 12805 5216 12817 5219
rect 12676 5188 12817 5216
rect 12676 5176 12682 5188
rect 12805 5185 12817 5188
rect 12851 5185 12863 5219
rect 12805 5179 12863 5185
rect 13265 5219 13323 5225
rect 13265 5185 13277 5219
rect 13311 5185 13323 5219
rect 15838 5216 15844 5228
rect 15799 5188 15844 5216
rect 13265 5179 13323 5185
rect 10318 5148 10324 5160
rect 9646 5120 9904 5148
rect 10279 5120 10324 5148
rect 9122 5040 9128 5092
rect 9180 5080 9186 5092
rect 9646 5080 9674 5120
rect 10318 5108 10324 5120
rect 10376 5108 10382 5160
rect 10502 5148 10508 5160
rect 10463 5120 10508 5148
rect 10502 5108 10508 5120
rect 10560 5108 10566 5160
rect 11793 5151 11851 5157
rect 11793 5117 11805 5151
rect 11839 5148 11851 5151
rect 11974 5148 11980 5160
rect 11839 5120 11980 5148
rect 11839 5117 11851 5120
rect 11793 5111 11851 5117
rect 11974 5108 11980 5120
rect 12032 5108 12038 5160
rect 12526 5148 12532 5160
rect 12487 5120 12532 5148
rect 12526 5108 12532 5120
rect 12584 5108 12590 5160
rect 12710 5148 12716 5160
rect 12671 5120 12716 5148
rect 12710 5108 12716 5120
rect 12768 5108 12774 5160
rect 9180 5052 9674 5080
rect 9180 5040 9186 5052
rect 9950 5040 9956 5092
rect 10008 5080 10014 5092
rect 10962 5080 10968 5092
rect 10008 5052 10968 5080
rect 10008 5040 10014 5052
rect 10962 5040 10968 5052
rect 11020 5040 11026 5092
rect 11606 5040 11612 5092
rect 11664 5080 11670 5092
rect 12345 5083 12403 5089
rect 11664 5052 12112 5080
rect 11664 5040 11670 5052
rect 7791 4984 8432 5012
rect 7791 4981 7803 4984
rect 7745 4975 7803 4981
rect 8478 4972 8484 5024
rect 8536 5012 8542 5024
rect 8754 5012 8760 5024
rect 8536 4984 8760 5012
rect 8536 4972 8542 4984
rect 8754 4972 8760 4984
rect 8812 4972 8818 5024
rect 9490 4972 9496 5024
rect 9548 5012 9554 5024
rect 11149 5015 11207 5021
rect 11149 5012 11161 5015
rect 9548 4984 11161 5012
rect 9548 4972 9554 4984
rect 11149 4981 11161 4984
rect 11195 5012 11207 5015
rect 11974 5012 11980 5024
rect 11195 4984 11980 5012
rect 11195 4981 11207 4984
rect 11149 4975 11207 4981
rect 11974 4972 11980 4984
rect 12032 4972 12038 5024
rect 12084 5012 12112 5052
rect 12345 5049 12357 5083
rect 12391 5080 12403 5083
rect 13280 5080 13308 5179
rect 15838 5176 15844 5188
rect 15896 5176 15902 5228
rect 20806 5216 20812 5228
rect 20767 5188 20812 5216
rect 20806 5176 20812 5188
rect 20864 5176 20870 5228
rect 15470 5148 15476 5160
rect 15431 5120 15476 5148
rect 15470 5108 15476 5120
rect 15528 5108 15534 5160
rect 15562 5108 15568 5160
rect 15620 5148 15626 5160
rect 15620 5120 15665 5148
rect 15620 5108 15626 5120
rect 12391 5052 13308 5080
rect 12391 5049 12403 5052
rect 12345 5043 12403 5049
rect 12894 5012 12900 5024
rect 12084 4984 12900 5012
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 13446 5012 13452 5024
rect 13407 4984 13452 5012
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 14826 4972 14832 5024
rect 14884 5012 14890 5024
rect 15013 5015 15071 5021
rect 15013 5012 15025 5015
rect 14884 4984 15025 5012
rect 14884 4972 14890 4984
rect 15013 4981 15025 4984
rect 15059 4981 15071 5015
rect 15013 4975 15071 4981
rect 16025 5015 16083 5021
rect 16025 4981 16037 5015
rect 16071 5012 16083 5015
rect 17034 5012 17040 5024
rect 16071 4984 17040 5012
rect 16071 4981 16083 4984
rect 16025 4975 16083 4981
rect 17034 4972 17040 4984
rect 17092 4972 17098 5024
rect 20625 5015 20683 5021
rect 20625 4981 20637 5015
rect 20671 5012 20683 5015
rect 20714 5012 20720 5024
rect 20671 4984 20720 5012
rect 20671 4981 20683 4984
rect 20625 4975 20683 4981
rect 20714 4972 20720 4984
rect 20772 4972 20778 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 4706 4768 4712 4820
rect 4764 4808 4770 4820
rect 5534 4808 5540 4820
rect 4764 4780 5540 4808
rect 4764 4768 4770 4780
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 5810 4808 5816 4820
rect 5771 4780 5816 4808
rect 5810 4768 5816 4780
rect 5868 4768 5874 4820
rect 5902 4768 5908 4820
rect 5960 4808 5966 4820
rect 6273 4811 6331 4817
rect 6273 4808 6285 4811
rect 5960 4780 6285 4808
rect 5960 4768 5966 4780
rect 6273 4777 6285 4780
rect 6319 4777 6331 4811
rect 7098 4808 7104 4820
rect 7059 4780 7104 4808
rect 6273 4771 6331 4777
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 8481 4811 8539 4817
rect 8481 4777 8493 4811
rect 8527 4808 8539 4811
rect 8570 4808 8576 4820
rect 8527 4780 8576 4808
rect 8527 4777 8539 4780
rect 8481 4771 8539 4777
rect 8570 4768 8576 4780
rect 8628 4768 8634 4820
rect 9033 4811 9091 4817
rect 9033 4777 9045 4811
rect 9079 4808 9091 4811
rect 9306 4808 9312 4820
rect 9079 4780 9312 4808
rect 9079 4777 9091 4780
rect 9033 4771 9091 4777
rect 4246 4740 4252 4752
rect 1964 4712 4252 4740
rect 1964 4681 1992 4712
rect 4246 4700 4252 4712
rect 4304 4740 4310 4752
rect 7006 4740 7012 4752
rect 4304 4712 7012 4740
rect 4304 4700 4310 4712
rect 7006 4700 7012 4712
rect 7064 4700 7070 4752
rect 1949 4675 2007 4681
rect 1949 4641 1961 4675
rect 1995 4641 2007 4675
rect 5166 4672 5172 4684
rect 5127 4644 5172 4672
rect 1949 4635 2007 4641
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5350 4632 5356 4684
rect 5408 4672 5414 4684
rect 6917 4675 6975 4681
rect 5408 4644 6868 4672
rect 5408 4632 5414 4644
rect 2222 4604 2228 4616
rect 2183 4576 2228 4604
rect 2222 4564 2228 4576
rect 2280 4604 2286 4616
rect 2317 4607 2375 4613
rect 2317 4604 2329 4607
rect 2280 4576 2329 4604
rect 2280 4564 2286 4576
rect 2317 4573 2329 4576
rect 2363 4573 2375 4607
rect 2317 4567 2375 4573
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4604 5503 4607
rect 5994 4604 6000 4616
rect 5491 4576 6000 4604
rect 5491 4573 5503 4576
rect 5445 4567 5503 4573
rect 5994 4564 6000 4576
rect 6052 4564 6058 4616
rect 6840 4604 6868 4644
rect 6917 4641 6929 4675
rect 6963 4672 6975 4675
rect 7116 4672 7144 4768
rect 7926 4700 7932 4752
rect 7984 4740 7990 4752
rect 9048 4740 9076 4771
rect 9306 4768 9312 4780
rect 9364 4768 9370 4820
rect 9766 4808 9772 4820
rect 9727 4780 9772 4808
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 10870 4808 10876 4820
rect 9968 4780 10876 4808
rect 9968 4740 9996 4780
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 11422 4808 11428 4820
rect 11383 4780 11428 4808
rect 11422 4768 11428 4780
rect 11480 4808 11486 4820
rect 11882 4808 11888 4820
rect 11480 4780 11888 4808
rect 11480 4768 11486 4780
rect 11882 4768 11888 4780
rect 11940 4768 11946 4820
rect 11974 4768 11980 4820
rect 12032 4808 12038 4820
rect 12345 4811 12403 4817
rect 12032 4780 12112 4808
rect 12032 4768 12038 4780
rect 7984 4712 9076 4740
rect 9140 4712 9996 4740
rect 7984 4700 7990 4712
rect 6963 4644 7144 4672
rect 6963 4641 6975 4644
rect 6917 4635 6975 4641
rect 7650 4632 7656 4684
rect 7708 4672 7714 4684
rect 7837 4675 7895 4681
rect 7837 4672 7849 4675
rect 7708 4644 7849 4672
rect 7708 4632 7714 4644
rect 7837 4641 7849 4644
rect 7883 4672 7895 4675
rect 8665 4675 8723 4681
rect 8665 4672 8677 4675
rect 7883 4644 8677 4672
rect 7883 4641 7895 4644
rect 7837 4635 7895 4641
rect 8665 4641 8677 4644
rect 8711 4672 8723 4675
rect 9140 4672 9168 4712
rect 10042 4700 10048 4752
rect 10100 4740 10106 4752
rect 10100 4712 10272 4740
rect 10100 4700 10106 4712
rect 8711 4644 9168 4672
rect 9677 4675 9735 4681
rect 8711 4641 8723 4644
rect 8665 4635 8723 4641
rect 9677 4641 9689 4675
rect 9723 4672 9735 4675
rect 9950 4672 9956 4684
rect 9723 4644 9956 4672
rect 9723 4641 9735 4644
rect 9677 4635 9735 4641
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 10244 4672 10272 4712
rect 10318 4700 10324 4752
rect 10376 4740 10382 4752
rect 10778 4740 10784 4752
rect 10376 4712 10784 4740
rect 10376 4700 10382 4712
rect 10428 4681 10456 4712
rect 10778 4700 10784 4712
rect 10836 4700 10842 4752
rect 10962 4740 10968 4752
rect 10923 4712 10968 4740
rect 10962 4700 10968 4712
rect 11020 4700 11026 4752
rect 11241 4743 11299 4749
rect 11241 4709 11253 4743
rect 11287 4740 11299 4743
rect 11330 4740 11336 4752
rect 11287 4712 11336 4740
rect 11287 4709 11299 4712
rect 11241 4703 11299 4709
rect 11330 4700 11336 4712
rect 11388 4700 11394 4752
rect 11606 4740 11612 4752
rect 11567 4712 11612 4740
rect 11606 4700 11612 4712
rect 11664 4700 11670 4752
rect 12084 4740 12112 4780
rect 12345 4777 12357 4811
rect 12391 4808 12403 4811
rect 12618 4808 12624 4820
rect 12391 4780 12624 4808
rect 12391 4777 12403 4780
rect 12345 4771 12403 4777
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 15470 4808 15476 4820
rect 15431 4780 15476 4808
rect 15470 4768 15476 4780
rect 15528 4768 15534 4820
rect 17494 4808 17500 4820
rect 16684 4780 17500 4808
rect 16684 4740 16712 4780
rect 17494 4768 17500 4780
rect 17552 4768 17558 4820
rect 18049 4811 18107 4817
rect 18049 4777 18061 4811
rect 18095 4808 18107 4811
rect 20254 4808 20260 4820
rect 18095 4780 20260 4808
rect 18095 4777 18107 4780
rect 18049 4771 18107 4777
rect 20254 4768 20260 4780
rect 20312 4768 20318 4820
rect 12084 4712 14964 4740
rect 10413 4675 10471 4681
rect 10244 4644 10364 4672
rect 8021 4607 8079 4613
rect 8021 4604 8033 4607
rect 6840 4576 8033 4604
rect 8021 4573 8033 4576
rect 8067 4604 8079 4607
rect 9766 4604 9772 4616
rect 8067 4576 9772 4604
rect 8067 4573 8079 4576
rect 8021 4567 8079 4573
rect 9766 4564 9772 4576
rect 9824 4604 9830 4616
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 9824 4576 10241 4604
rect 9824 4564 9830 4576
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 10336 4604 10364 4644
rect 10413 4641 10425 4675
rect 10459 4641 10471 4675
rect 14826 4672 14832 4684
rect 14787 4644 14832 4672
rect 10413 4635 10471 4641
rect 14826 4632 14832 4644
rect 14884 4632 14890 4684
rect 10597 4607 10655 4613
rect 10597 4604 10609 4607
rect 10336 4576 10609 4604
rect 10229 4567 10287 4573
rect 10597 4573 10609 4576
rect 10643 4573 10655 4607
rect 10597 4567 10655 4573
rect 10870 4564 10876 4616
rect 10928 4604 10934 4616
rect 11885 4607 11943 4613
rect 11885 4604 11897 4607
rect 10928 4576 11897 4604
rect 10928 4564 10934 4576
rect 11885 4573 11897 4576
rect 11931 4573 11943 4607
rect 14734 4604 14740 4616
rect 14695 4576 14740 4604
rect 11885 4567 11943 4573
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 14936 4604 14964 4712
rect 15028 4712 16712 4740
rect 16761 4743 16819 4749
rect 15028 4681 15056 4712
rect 16761 4709 16773 4743
rect 16807 4740 16819 4743
rect 16942 4740 16948 4752
rect 16807 4712 16948 4740
rect 16807 4709 16819 4712
rect 16761 4703 16819 4709
rect 16942 4700 16948 4712
rect 17000 4700 17006 4752
rect 15013 4675 15071 4681
rect 15013 4641 15025 4675
rect 15059 4641 15071 4675
rect 16022 4672 16028 4684
rect 15983 4644 16028 4672
rect 15013 4635 15071 4641
rect 16022 4632 16028 4644
rect 16080 4672 16086 4684
rect 16393 4675 16451 4681
rect 16393 4672 16405 4675
rect 16080 4644 16405 4672
rect 16080 4632 16086 4644
rect 16393 4641 16405 4644
rect 16439 4641 16451 4675
rect 16393 4635 16451 4641
rect 17497 4675 17555 4681
rect 17497 4641 17509 4675
rect 17543 4672 17555 4675
rect 17586 4672 17592 4684
rect 17543 4644 17592 4672
rect 17543 4641 17555 4644
rect 17497 4635 17555 4641
rect 17586 4632 17592 4644
rect 17644 4632 17650 4684
rect 15930 4604 15936 4616
rect 14936 4576 15936 4604
rect 15930 4564 15936 4576
rect 15988 4564 15994 4616
rect 16298 4564 16304 4616
rect 16356 4604 16362 4616
rect 16577 4607 16635 4613
rect 16577 4604 16589 4607
rect 16356 4576 16589 4604
rect 16356 4564 16362 4576
rect 16577 4573 16589 4576
rect 16623 4604 16635 4607
rect 16853 4607 16911 4613
rect 16853 4604 16865 4607
rect 16623 4576 16865 4604
rect 16623 4573 16635 4576
rect 16577 4567 16635 4573
rect 16853 4573 16865 4576
rect 16899 4573 16911 4607
rect 18782 4604 18788 4616
rect 18743 4576 18788 4604
rect 16853 4567 16911 4573
rect 18782 4564 18788 4576
rect 18840 4564 18846 4616
rect 4522 4496 4528 4548
rect 4580 4536 4586 4548
rect 5353 4539 5411 4545
rect 5353 4536 5365 4539
rect 4580 4508 5365 4536
rect 4580 4496 4586 4508
rect 5353 4505 5365 4508
rect 5399 4505 5411 4539
rect 5353 4499 5411 4505
rect 5534 4496 5540 4548
rect 5592 4536 5598 4548
rect 6641 4539 6699 4545
rect 6641 4536 6653 4539
rect 5592 4508 6653 4536
rect 5592 4496 5598 4508
rect 6641 4505 6653 4508
rect 6687 4505 6699 4539
rect 6641 4499 6699 4505
rect 6914 4496 6920 4548
rect 6972 4536 6978 4548
rect 8113 4539 8171 4545
rect 8113 4536 8125 4539
rect 6972 4508 8125 4536
rect 6972 4496 6978 4508
rect 8113 4505 8125 4508
rect 8159 4505 8171 4539
rect 10781 4539 10839 4545
rect 10781 4536 10793 4539
rect 8113 4499 8171 4505
rect 9508 4508 10793 4536
rect 9508 4480 9536 4508
rect 10781 4505 10793 4508
rect 10827 4505 10839 4539
rect 10781 4499 10839 4505
rect 11330 4496 11336 4548
rect 11388 4536 11394 4548
rect 11388 4508 11928 4536
rect 11388 4496 11394 4508
rect 5902 4428 5908 4480
rect 5960 4468 5966 4480
rect 6730 4468 6736 4480
rect 5960 4440 6005 4468
rect 6643 4440 6736 4468
rect 5960 4428 5966 4440
rect 6730 4428 6736 4440
rect 6788 4468 6794 4480
rect 7285 4471 7343 4477
rect 7285 4468 7297 4471
rect 6788 4440 7297 4468
rect 6788 4428 6794 4440
rect 7285 4437 7297 4440
rect 7331 4468 7343 4471
rect 8018 4468 8024 4480
rect 7331 4440 8024 4468
rect 7331 4437 7343 4440
rect 7285 4431 7343 4437
rect 8018 4428 8024 4440
rect 8076 4428 8082 4480
rect 8202 4428 8208 4480
rect 8260 4468 8266 4480
rect 9306 4468 9312 4480
rect 8260 4440 9312 4468
rect 8260 4428 8266 4440
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 9401 4471 9459 4477
rect 9401 4437 9413 4471
rect 9447 4468 9459 4471
rect 9490 4468 9496 4480
rect 9447 4440 9496 4468
rect 9447 4437 9459 4440
rect 9401 4431 9459 4437
rect 9490 4428 9496 4440
rect 9548 4428 9554 4480
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 10137 4471 10195 4477
rect 10137 4468 10149 4471
rect 9732 4440 10149 4468
rect 9732 4428 9738 4440
rect 10137 4437 10149 4440
rect 10183 4437 10195 4471
rect 11698 4468 11704 4480
rect 11659 4440 11704 4468
rect 10137 4431 10195 4437
rect 11698 4428 11704 4440
rect 11756 4428 11762 4480
rect 11900 4468 11928 4508
rect 12618 4496 12624 4548
rect 12676 4536 12682 4548
rect 17954 4536 17960 4548
rect 12676 4508 17960 4536
rect 12676 4496 12682 4508
rect 17954 4496 17960 4508
rect 18012 4496 18018 4548
rect 11974 4468 11980 4480
rect 11900 4440 11980 4468
rect 11974 4428 11980 4440
rect 12032 4428 12038 4480
rect 12069 4471 12127 4477
rect 12069 4437 12081 4471
rect 12115 4468 12127 4471
rect 12710 4468 12716 4480
rect 12115 4440 12716 4468
rect 12115 4437 12127 4440
rect 12069 4431 12127 4437
rect 12710 4428 12716 4440
rect 12768 4468 12774 4480
rect 13722 4468 13728 4480
rect 12768 4440 13728 4468
rect 12768 4428 12774 4440
rect 13722 4428 13728 4440
rect 13780 4428 13786 4480
rect 14366 4468 14372 4480
rect 14327 4440 14372 4468
rect 14366 4428 14372 4440
rect 14424 4428 14430 4480
rect 15838 4468 15844 4480
rect 15799 4440 15844 4468
rect 15838 4428 15844 4440
rect 15896 4428 15902 4480
rect 15930 4428 15936 4480
rect 15988 4468 15994 4480
rect 17586 4468 17592 4480
rect 15988 4440 16033 4468
rect 17547 4440 17592 4468
rect 15988 4428 15994 4440
rect 17586 4428 17592 4440
rect 17644 4428 17650 4480
rect 17678 4428 17684 4480
rect 17736 4468 17742 4480
rect 18969 4471 19027 4477
rect 17736 4440 17781 4468
rect 17736 4428 17742 4440
rect 18969 4437 18981 4471
rect 19015 4468 19027 4471
rect 19886 4468 19892 4480
rect 19015 4440 19892 4468
rect 19015 4437 19027 4440
rect 18969 4431 19027 4437
rect 19886 4428 19892 4440
rect 19944 4428 19950 4480
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 5813 4267 5871 4273
rect 5813 4233 5825 4267
rect 5859 4264 5871 4267
rect 5902 4264 5908 4276
rect 5859 4236 5908 4264
rect 5859 4233 5871 4236
rect 5813 4227 5871 4233
rect 5902 4224 5908 4236
rect 5960 4224 5966 4276
rect 8386 4224 8392 4276
rect 8444 4264 8450 4276
rect 8941 4267 8999 4273
rect 8444 4236 8892 4264
rect 8444 4224 8450 4236
rect 2590 4156 2596 4208
rect 2648 4196 2654 4208
rect 5350 4196 5356 4208
rect 2648 4168 5356 4196
rect 2648 4156 2654 4168
rect 5350 4156 5356 4168
rect 5408 4156 5414 4208
rect 5718 4156 5724 4208
rect 5776 4196 5782 4208
rect 6733 4199 6791 4205
rect 6733 4196 6745 4199
rect 5776 4168 6745 4196
rect 5776 4156 5782 4168
rect 6733 4165 6745 4168
rect 6779 4196 6791 4199
rect 6822 4196 6828 4208
rect 6779 4168 6828 4196
rect 6779 4165 6791 4168
rect 6733 4159 6791 4165
rect 6822 4156 6828 4168
rect 6880 4156 6886 4208
rect 7190 4156 7196 4208
rect 7248 4196 7254 4208
rect 7745 4199 7803 4205
rect 7745 4196 7757 4199
rect 7248 4168 7757 4196
rect 7248 4156 7254 4168
rect 7745 4165 7757 4168
rect 7791 4196 7803 4199
rect 7791 4168 8432 4196
rect 7791 4165 7803 4168
rect 7745 4159 7803 4165
rect 1946 4128 1952 4140
rect 1907 4100 1952 4128
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 2038 4088 2044 4140
rect 2096 4128 2102 4140
rect 2682 4128 2688 4140
rect 2096 4100 2688 4128
rect 2096 4088 2102 4100
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 7650 4128 7656 4140
rect 4120 4100 7656 4128
rect 4120 4088 4126 4100
rect 2222 4060 2228 4072
rect 2183 4032 2228 4060
rect 2222 4020 2228 4032
rect 2280 4060 2286 4072
rect 2501 4063 2559 4069
rect 2501 4060 2513 4063
rect 2280 4032 2513 4060
rect 2280 4020 2286 4032
rect 2501 4029 2513 4032
rect 2547 4029 2559 4063
rect 2501 4023 2559 4029
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4029 5687 4063
rect 5629 4023 5687 4029
rect 4246 3952 4252 4004
rect 4304 3992 4310 4004
rect 5644 3992 5672 4023
rect 5718 4020 5724 4072
rect 5776 4060 5782 4072
rect 6840 4069 6868 4100
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 8404 4128 8432 4168
rect 8478 4156 8484 4208
rect 8536 4196 8542 4208
rect 8864 4196 8892 4236
rect 8941 4233 8953 4267
rect 8987 4264 8999 4267
rect 9122 4264 9128 4276
rect 8987 4236 9128 4264
rect 8987 4233 8999 4236
rect 8941 4227 8999 4233
rect 9122 4224 9128 4236
rect 9180 4224 9186 4276
rect 9398 4224 9404 4276
rect 9456 4264 9462 4276
rect 9674 4264 9680 4276
rect 9456 4236 9680 4264
rect 9456 4224 9462 4236
rect 9674 4224 9680 4236
rect 9732 4224 9738 4276
rect 10042 4264 10048 4276
rect 10003 4236 10048 4264
rect 10042 4224 10048 4236
rect 10100 4264 10106 4276
rect 10318 4264 10324 4276
rect 10100 4236 10324 4264
rect 10100 4224 10106 4236
rect 10318 4224 10324 4236
rect 10376 4224 10382 4276
rect 10502 4264 10508 4276
rect 10463 4236 10508 4264
rect 10502 4224 10508 4236
rect 10560 4224 10566 4276
rect 11606 4264 11612 4276
rect 10612 4236 11612 4264
rect 9306 4196 9312 4208
rect 8536 4168 8581 4196
rect 8864 4168 9312 4196
rect 8536 4156 8542 4168
rect 9306 4156 9312 4168
rect 9364 4156 9370 4208
rect 9490 4156 9496 4208
rect 9548 4196 9554 4208
rect 9548 4168 10548 4196
rect 9548 4156 9554 4168
rect 10520 4140 10548 4168
rect 8573 4131 8631 4137
rect 8573 4128 8585 4131
rect 8404 4100 8585 4128
rect 8573 4097 8585 4100
rect 8619 4097 8631 4131
rect 10137 4131 10195 4137
rect 10137 4128 10149 4131
rect 8573 4091 8631 4097
rect 10060 4100 10149 4128
rect 6825 4063 6883 4069
rect 5776 4032 5821 4060
rect 5776 4020 5782 4032
rect 6825 4029 6837 4063
rect 6871 4029 6883 4063
rect 7006 4060 7012 4072
rect 6967 4032 7012 4060
rect 6825 4023 6883 4029
rect 7006 4020 7012 4032
rect 7064 4020 7070 4072
rect 7561 4063 7619 4069
rect 7561 4029 7573 4063
rect 7607 4029 7619 4063
rect 7561 4023 7619 4029
rect 6546 3992 6552 4004
rect 4304 3964 6552 3992
rect 4304 3952 4310 3964
rect 6546 3952 6552 3964
rect 6604 3952 6610 4004
rect 1302 3884 1308 3936
rect 1360 3924 1366 3936
rect 2317 3927 2375 3933
rect 2317 3924 2329 3927
rect 1360 3896 2329 3924
rect 1360 3884 1366 3896
rect 2317 3893 2329 3896
rect 2363 3893 2375 3927
rect 2317 3887 2375 3893
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 2832 3896 2877 3924
rect 2832 3884 2838 3896
rect 2958 3884 2964 3936
rect 3016 3924 3022 3936
rect 6178 3924 6184 3936
rect 3016 3896 3061 3924
rect 6139 3896 6184 3924
rect 3016 3884 3022 3896
rect 6178 3884 6184 3896
rect 6236 3884 6242 3936
rect 6365 3927 6423 3933
rect 6365 3893 6377 3927
rect 6411 3924 6423 3927
rect 6730 3924 6736 3936
rect 6411 3896 6736 3924
rect 6411 3893 6423 3896
rect 6365 3887 6423 3893
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 7576 3924 7604 4023
rect 8018 4020 8024 4072
rect 8076 4060 8082 4072
rect 8389 4063 8447 4069
rect 8076 4032 8340 4060
rect 8076 4020 8082 4032
rect 7926 3924 7932 3936
rect 7576 3896 7932 3924
rect 7926 3884 7932 3896
rect 7984 3884 7990 3936
rect 8110 3924 8116 3936
rect 8071 3896 8116 3924
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 8312 3924 8340 4032
rect 8389 4029 8401 4063
rect 8435 4060 8447 4063
rect 9030 4060 9036 4072
rect 8435 4032 9036 4060
rect 8435 4029 8447 4032
rect 8389 4023 8447 4029
rect 9030 4020 9036 4032
rect 9088 4020 9094 4072
rect 9217 4063 9275 4069
rect 9217 4029 9229 4063
rect 9263 4060 9275 4063
rect 9950 4060 9956 4072
rect 9263 4032 9956 4060
rect 9263 4029 9275 4032
rect 9217 4023 9275 4029
rect 9950 4020 9956 4032
rect 10008 4020 10014 4072
rect 9582 3952 9588 4004
rect 9640 3992 9646 4004
rect 9677 3995 9735 4001
rect 9677 3992 9689 3995
rect 9640 3964 9689 3992
rect 9640 3952 9646 3964
rect 9677 3961 9689 3964
rect 9723 3961 9735 3995
rect 10060 3992 10088 4100
rect 10137 4097 10149 4100
rect 10183 4128 10195 4131
rect 10183 4100 10456 4128
rect 10183 4097 10195 4100
rect 10137 4091 10195 4097
rect 10226 4060 10232 4072
rect 10187 4032 10232 4060
rect 10226 4020 10232 4032
rect 10284 4020 10290 4072
rect 10428 4060 10456 4100
rect 10502 4088 10508 4140
rect 10560 4088 10566 4140
rect 10612 4060 10640 4236
rect 11606 4224 11612 4236
rect 11664 4224 11670 4276
rect 11882 4264 11888 4276
rect 11843 4236 11888 4264
rect 11882 4224 11888 4236
rect 11940 4224 11946 4276
rect 11974 4224 11980 4276
rect 12032 4264 12038 4276
rect 12437 4267 12495 4273
rect 12437 4264 12449 4267
rect 12032 4236 12077 4264
rect 12176 4236 12449 4264
rect 12032 4224 12038 4236
rect 11054 4156 11060 4208
rect 11112 4196 11118 4208
rect 11112 4168 11192 4196
rect 11112 4156 11118 4168
rect 10870 4128 10876 4140
rect 10831 4100 10876 4128
rect 10870 4088 10876 4100
rect 10928 4088 10934 4140
rect 10965 4131 11023 4137
rect 10965 4097 10977 4131
rect 11011 4128 11023 4131
rect 11011 4100 11100 4128
rect 11011 4097 11023 4100
rect 10965 4091 11023 4097
rect 10428 4032 10640 4060
rect 9677 3955 9735 3961
rect 9968 3964 10088 3992
rect 11072 3992 11100 4100
rect 11164 4069 11192 4168
rect 11149 4063 11207 4069
rect 11149 4029 11161 4063
rect 11195 4029 11207 4063
rect 11149 4023 11207 4029
rect 11330 4020 11336 4072
rect 11388 4060 11394 4072
rect 12176 4069 12204 4236
rect 12437 4233 12449 4236
rect 12483 4264 12495 4267
rect 12986 4264 12992 4276
rect 12483 4236 12992 4264
rect 12483 4233 12495 4236
rect 12437 4227 12495 4233
rect 12986 4224 12992 4236
rect 13044 4224 13050 4276
rect 15930 4224 15936 4276
rect 15988 4264 15994 4276
rect 16669 4267 16727 4273
rect 16669 4264 16681 4267
rect 15988 4236 16681 4264
rect 15988 4224 15994 4236
rect 16669 4233 16681 4236
rect 16715 4233 16727 4267
rect 17586 4264 17592 4276
rect 17547 4236 17592 4264
rect 16669 4227 16727 4233
rect 17586 4224 17592 4236
rect 17644 4224 17650 4276
rect 18506 4264 18512 4276
rect 18467 4236 18512 4264
rect 18506 4224 18512 4236
rect 18564 4224 18570 4276
rect 17037 4199 17095 4205
rect 17037 4196 17049 4199
rect 16132 4168 17049 4196
rect 14366 4128 14372 4140
rect 14327 4100 14372 4128
rect 14366 4088 14372 4100
rect 14424 4088 14430 4140
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 11388 4032 12173 4060
rect 11388 4020 11394 4032
rect 12161 4029 12173 4032
rect 12207 4029 12219 4063
rect 12161 4023 12219 4029
rect 12342 4020 12348 4072
rect 12400 4060 12406 4072
rect 12713 4063 12771 4069
rect 12713 4060 12725 4063
rect 12400 4032 12725 4060
rect 12400 4020 12406 4032
rect 12713 4029 12725 4032
rect 12759 4029 12771 4063
rect 12713 4023 12771 4029
rect 13630 4020 13636 4072
rect 13688 4060 13694 4072
rect 16132 4069 16160 4168
rect 17037 4165 17049 4168
rect 17083 4196 17095 4199
rect 17862 4196 17868 4208
rect 17083 4168 17868 4196
rect 17083 4165 17095 4168
rect 17037 4159 17095 4165
rect 17862 4156 17868 4168
rect 17920 4156 17926 4208
rect 16298 4128 16304 4140
rect 16259 4100 16304 4128
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 17218 4088 17224 4140
rect 17276 4128 17282 4140
rect 17276 4100 17448 4128
rect 17276 4088 17282 4100
rect 16117 4063 16175 4069
rect 16117 4060 16129 4063
rect 13688 4032 16129 4060
rect 13688 4020 13694 4032
rect 16117 4029 16129 4032
rect 16163 4029 16175 4063
rect 16316 4060 16344 4088
rect 17129 4063 17187 4069
rect 17129 4060 17141 4063
rect 16316 4032 17141 4060
rect 16117 4023 16175 4029
rect 17129 4029 17141 4032
rect 17175 4029 17187 4063
rect 17129 4023 17187 4029
rect 17313 4063 17371 4069
rect 17313 4029 17325 4063
rect 17359 4029 17371 4063
rect 17420 4060 17448 4100
rect 17586 4088 17592 4140
rect 17644 4128 17650 4140
rect 17957 4131 18015 4137
rect 17957 4128 17969 4131
rect 17644 4100 17969 4128
rect 17644 4088 17650 4100
rect 17957 4097 17969 4100
rect 18003 4097 18015 4131
rect 17957 4091 18015 4097
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 17420 4032 18061 4060
rect 17313 4023 17371 4029
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 18049 4023 18107 4029
rect 18233 4063 18291 4069
rect 18233 4029 18245 4063
rect 18279 4060 18291 4063
rect 18506 4060 18512 4072
rect 18279 4032 18512 4060
rect 18279 4029 18291 4032
rect 18233 4023 18291 4029
rect 11517 3995 11575 4001
rect 11517 3992 11529 3995
rect 11072 3964 11529 3992
rect 9493 3927 9551 3933
rect 9493 3924 9505 3927
rect 8312 3896 9505 3924
rect 9493 3893 9505 3896
rect 9539 3924 9551 3927
rect 9968 3924 9996 3964
rect 11517 3961 11529 3964
rect 11563 3961 11575 3995
rect 15838 3992 15844 4004
rect 11517 3955 11575 3961
rect 12406 3964 15844 3992
rect 9539 3896 9996 3924
rect 9539 3893 9551 3896
rect 9493 3887 9551 3893
rect 10042 3884 10048 3936
rect 10100 3924 10106 3936
rect 12406 3924 12434 3964
rect 15838 3952 15844 3964
rect 15896 3952 15902 4004
rect 17328 3992 17356 4023
rect 18506 4020 18512 4032
rect 18564 4020 18570 4072
rect 20990 3992 20996 4004
rect 17328 3964 20996 3992
rect 20990 3952 20996 3964
rect 21048 3952 21054 4004
rect 12618 3924 12624 3936
rect 10100 3896 12434 3924
rect 12579 3896 12624 3924
rect 10100 3884 10106 3896
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 12894 3924 12900 3936
rect 12855 3896 12900 3924
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 14553 3927 14611 3933
rect 14553 3893 14565 3927
rect 14599 3924 14611 3927
rect 14918 3924 14924 3936
rect 14599 3896 14924 3924
rect 14599 3893 14611 3896
rect 14553 3887 14611 3893
rect 14918 3884 14924 3896
rect 14976 3884 14982 3936
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 382 3680 388 3732
rect 440 3720 446 3732
rect 2314 3720 2320 3732
rect 440 3692 2320 3720
rect 440 3680 446 3692
rect 2314 3680 2320 3692
rect 2372 3720 2378 3732
rect 2685 3723 2743 3729
rect 2685 3720 2697 3723
rect 2372 3692 2697 3720
rect 2372 3680 2378 3692
rect 2685 3689 2697 3692
rect 2731 3689 2743 3723
rect 2685 3683 2743 3689
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 7006 3720 7012 3732
rect 5132 3692 7012 3720
rect 5132 3680 5138 3692
rect 1670 3652 1676 3664
rect 1631 3624 1676 3652
rect 1670 3612 1676 3624
rect 1728 3612 1734 3664
rect 2041 3655 2099 3661
rect 2041 3621 2053 3655
rect 2087 3652 2099 3655
rect 2406 3652 2412 3664
rect 2087 3624 2412 3652
rect 2087 3621 2099 3624
rect 2041 3615 2099 3621
rect 2406 3612 2412 3624
rect 2464 3612 2470 3664
rect 2590 3652 2596 3664
rect 2551 3624 2596 3652
rect 2590 3612 2596 3624
rect 2648 3612 2654 3664
rect 3970 3612 3976 3664
rect 4028 3652 4034 3664
rect 4801 3655 4859 3661
rect 4028 3624 4752 3652
rect 4028 3612 4034 3624
rect 2774 3584 2780 3596
rect 1504 3556 2780 3584
rect 1504 3528 1532 3556
rect 2774 3544 2780 3556
rect 2832 3544 2838 3596
rect 4246 3584 4252 3596
rect 4207 3556 4252 3584
rect 4246 3544 4252 3556
rect 4304 3544 4310 3596
rect 4724 3584 4752 3624
rect 4801 3621 4813 3655
rect 4847 3652 4859 3655
rect 4847 3624 5488 3652
rect 4847 3621 4859 3624
rect 4801 3615 4859 3621
rect 4724 3556 5304 3584
rect 1486 3516 1492 3528
rect 1399 3488 1492 3516
rect 1486 3476 1492 3488
rect 1544 3476 1550 3528
rect 2133 3519 2191 3525
rect 2133 3516 2145 3519
rect 1688 3488 2145 3516
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 1688 3448 1716 3488
rect 2133 3485 2145 3488
rect 2179 3485 2191 3519
rect 2133 3479 2191 3485
rect 2314 3476 2320 3528
rect 2372 3516 2378 3528
rect 2409 3519 2467 3525
rect 2409 3516 2421 3519
rect 2372 3488 2421 3516
rect 2372 3476 2378 3488
rect 2409 3485 2421 3488
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 1854 3448 1860 3460
rect 1360 3420 1716 3448
rect 1815 3420 1860 3448
rect 1360 3408 1366 3420
rect 1854 3408 1860 3420
rect 1912 3448 1918 3460
rect 5276 3457 5304 3556
rect 5460 3516 5488 3624
rect 5552 3593 5580 3692
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 7101 3723 7159 3729
rect 7101 3689 7113 3723
rect 7147 3720 7159 3723
rect 10505 3723 10563 3729
rect 7147 3692 9536 3720
rect 7147 3689 7159 3692
rect 7101 3683 7159 3689
rect 6380 3624 9260 3652
rect 5537 3587 5595 3593
rect 5537 3553 5549 3587
rect 5583 3553 5595 3587
rect 5537 3547 5595 3553
rect 6380 3516 6408 3624
rect 6546 3584 6552 3596
rect 6507 3556 6552 3584
rect 6546 3544 6552 3556
rect 6604 3544 6610 3596
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 8938 3584 8944 3596
rect 7708 3556 8944 3584
rect 7708 3544 7714 3556
rect 8938 3544 8944 3556
rect 8996 3544 9002 3596
rect 9122 3584 9128 3596
rect 9083 3556 9128 3584
rect 9122 3544 9128 3556
rect 9180 3544 9186 3596
rect 9232 3593 9260 3624
rect 9217 3587 9275 3593
rect 9217 3553 9229 3587
rect 9263 3553 9275 3587
rect 9217 3547 9275 3553
rect 6730 3516 6736 3528
rect 5460 3488 6408 3516
rect 6691 3488 6736 3516
rect 6730 3476 6736 3488
rect 6788 3476 6794 3528
rect 7377 3519 7435 3525
rect 7377 3516 7389 3519
rect 7300 3488 7389 3516
rect 3053 3451 3111 3457
rect 3053 3448 3065 3451
rect 1912 3420 3065 3448
rect 1912 3408 1918 3420
rect 3053 3417 3065 3420
rect 3099 3417 3111 3451
rect 3053 3411 3111 3417
rect 4433 3451 4491 3457
rect 4433 3417 4445 3451
rect 4479 3448 4491 3451
rect 5261 3451 5319 3457
rect 4479 3420 4936 3448
rect 4479 3417 4491 3420
rect 4433 3411 4491 3417
rect 2314 3380 2320 3392
rect 2275 3352 2320 3380
rect 2314 3340 2320 3352
rect 2372 3340 2378 3392
rect 2774 3340 2780 3392
rect 2832 3380 2838 3392
rect 2869 3383 2927 3389
rect 2869 3380 2881 3383
rect 2832 3352 2881 3380
rect 2832 3340 2838 3352
rect 2869 3349 2881 3352
rect 2915 3349 2927 3383
rect 2869 3343 2927 3349
rect 3142 3340 3148 3392
rect 3200 3380 3206 3392
rect 3237 3383 3295 3389
rect 3237 3380 3249 3383
rect 3200 3352 3249 3380
rect 3200 3340 3206 3352
rect 3237 3349 3249 3352
rect 3283 3349 3295 3383
rect 3418 3380 3424 3392
rect 3379 3352 3424 3380
rect 3237 3343 3295 3349
rect 3418 3340 3424 3352
rect 3476 3340 3482 3392
rect 4246 3340 4252 3392
rect 4304 3380 4310 3392
rect 4908 3389 4936 3420
rect 5261 3417 5273 3451
rect 5307 3417 5319 3451
rect 7190 3448 7196 3460
rect 5261 3411 5319 3417
rect 5368 3420 7196 3448
rect 5368 3392 5396 3420
rect 7190 3408 7196 3420
rect 7248 3408 7254 3460
rect 7300 3392 7328 3488
rect 7377 3485 7389 3488
rect 7423 3485 7435 3519
rect 7377 3479 7435 3485
rect 8297 3519 8355 3525
rect 8297 3485 8309 3519
rect 8343 3516 8355 3519
rect 8573 3519 8631 3525
rect 8573 3516 8585 3519
rect 8343 3488 8585 3516
rect 8343 3485 8355 3488
rect 8297 3479 8355 3485
rect 8573 3485 8585 3488
rect 8619 3516 8631 3519
rect 8662 3516 8668 3528
rect 8619 3488 8668 3516
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 8662 3476 8668 3488
rect 8720 3476 8726 3528
rect 9306 3516 9312 3528
rect 9267 3488 9312 3516
rect 9306 3476 9312 3488
rect 9364 3476 9370 3528
rect 9508 3516 9536 3692
rect 10505 3689 10517 3723
rect 10551 3720 10563 3723
rect 10870 3720 10876 3732
rect 10551 3692 10876 3720
rect 10551 3689 10563 3692
rect 10505 3683 10563 3689
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 12437 3723 12495 3729
rect 12437 3689 12449 3723
rect 12483 3720 12495 3723
rect 12483 3692 13768 3720
rect 12483 3689 12495 3692
rect 12437 3683 12495 3689
rect 9677 3655 9735 3661
rect 9677 3621 9689 3655
rect 9723 3652 9735 3655
rect 13740 3652 13768 3692
rect 13814 3680 13820 3732
rect 13872 3720 13878 3732
rect 14090 3720 14096 3732
rect 13872 3692 14096 3720
rect 13872 3680 13878 3692
rect 14090 3680 14096 3692
rect 14148 3680 14154 3732
rect 17218 3720 17224 3732
rect 17179 3692 17224 3720
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 17862 3680 17868 3732
rect 17920 3720 17926 3732
rect 18417 3723 18475 3729
rect 18417 3720 18429 3723
rect 17920 3692 18429 3720
rect 17920 3680 17926 3692
rect 18417 3689 18429 3692
rect 18463 3689 18475 3723
rect 18417 3683 18475 3689
rect 19518 3680 19524 3732
rect 19576 3720 19582 3732
rect 19981 3723 20039 3729
rect 19981 3720 19993 3723
rect 19576 3692 19993 3720
rect 19576 3680 19582 3692
rect 19981 3689 19993 3692
rect 20027 3720 20039 3723
rect 20346 3720 20352 3732
rect 20027 3692 20352 3720
rect 20027 3689 20039 3692
rect 19981 3683 20039 3689
rect 20346 3680 20352 3692
rect 20404 3680 20410 3732
rect 21358 3720 21364 3732
rect 21319 3692 21364 3720
rect 21358 3680 21364 3692
rect 21416 3680 21422 3732
rect 14550 3652 14556 3664
rect 9723 3624 13400 3652
rect 13740 3624 14556 3652
rect 9723 3621 9735 3624
rect 9677 3615 9735 3621
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 9861 3587 9919 3593
rect 9861 3584 9873 3587
rect 9640 3556 9873 3584
rect 9640 3544 9646 3556
rect 9861 3553 9873 3556
rect 9907 3553 9919 3587
rect 10042 3584 10048 3596
rect 10003 3556 10048 3584
rect 9861 3547 9919 3553
rect 10042 3544 10048 3556
rect 10100 3544 10106 3596
rect 10686 3584 10692 3596
rect 10647 3556 10692 3584
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 11514 3584 11520 3596
rect 11475 3556 11520 3584
rect 11514 3544 11520 3556
rect 11572 3544 11578 3596
rect 11606 3544 11612 3596
rect 11664 3584 11670 3596
rect 12529 3587 12587 3593
rect 12529 3584 12541 3587
rect 11664 3556 12541 3584
rect 11664 3544 11670 3556
rect 12268 3525 12296 3556
rect 12529 3553 12541 3556
rect 12575 3553 12587 3587
rect 12529 3547 12587 3553
rect 12805 3587 12863 3593
rect 12805 3553 12817 3587
rect 12851 3584 12863 3587
rect 13078 3584 13084 3596
rect 12851 3556 13084 3584
rect 12851 3553 12863 3556
rect 12805 3547 12863 3553
rect 13078 3544 13084 3556
rect 13136 3544 13142 3596
rect 13173 3587 13231 3593
rect 13173 3553 13185 3587
rect 13219 3584 13231 3587
rect 13262 3584 13268 3596
rect 13219 3556 13268 3584
rect 13219 3553 13231 3556
rect 13173 3547 13231 3553
rect 13262 3544 13268 3556
rect 13320 3544 13326 3596
rect 13372 3525 13400 3624
rect 14550 3612 14556 3624
rect 14608 3612 14614 3664
rect 16206 3612 16212 3664
rect 16264 3652 16270 3664
rect 17405 3655 17463 3661
rect 17405 3652 17417 3655
rect 16264 3624 17417 3652
rect 16264 3612 16270 3624
rect 17405 3621 17417 3624
rect 17451 3652 17463 3655
rect 17586 3652 17592 3664
rect 17451 3624 17592 3652
rect 17451 3621 17463 3624
rect 17405 3615 17463 3621
rect 17586 3612 17592 3624
rect 17644 3652 17650 3664
rect 18874 3652 18880 3664
rect 17644 3624 18880 3652
rect 17644 3612 17650 3624
rect 18874 3612 18880 3624
rect 18932 3612 18938 3664
rect 11793 3519 11851 3525
rect 11793 3516 11805 3519
rect 9508 3488 11805 3516
rect 11793 3485 11805 3488
rect 11839 3485 11851 3519
rect 11793 3479 11851 3485
rect 12253 3519 12311 3525
rect 12253 3485 12265 3519
rect 12299 3485 12311 3519
rect 12253 3479 12311 3485
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3485 13415 3519
rect 13817 3519 13875 3525
rect 13817 3516 13829 3519
rect 13357 3479 13415 3485
rect 13464 3488 13829 3516
rect 8205 3451 8263 3457
rect 8205 3417 8217 3451
rect 8251 3448 8263 3451
rect 8386 3448 8392 3460
rect 8251 3420 8392 3448
rect 8251 3417 8263 3420
rect 8205 3411 8263 3417
rect 8386 3408 8392 3420
rect 8444 3408 8450 3460
rect 8757 3451 8815 3457
rect 8757 3417 8769 3451
rect 8803 3448 8815 3451
rect 9490 3448 9496 3460
rect 8803 3420 9496 3448
rect 8803 3417 8815 3420
rect 8757 3411 8815 3417
rect 9490 3408 9496 3420
rect 9548 3408 9554 3460
rect 10873 3451 10931 3457
rect 10873 3417 10885 3451
rect 10919 3448 10931 3451
rect 11882 3448 11888 3460
rect 10919 3420 11888 3448
rect 10919 3417 10931 3420
rect 10873 3411 10931 3417
rect 11882 3408 11888 3420
rect 11940 3408 11946 3460
rect 13265 3451 13323 3457
rect 13265 3448 13277 3451
rect 12176 3420 13277 3448
rect 4341 3383 4399 3389
rect 4341 3380 4353 3383
rect 4304 3352 4353 3380
rect 4304 3340 4310 3352
rect 4341 3349 4353 3352
rect 4387 3349 4399 3383
rect 4341 3343 4399 3349
rect 4893 3383 4951 3389
rect 4893 3349 4905 3383
rect 4939 3349 4951 3383
rect 5350 3380 5356 3392
rect 5311 3352 5356 3380
rect 4893 3343 4951 3349
rect 5350 3340 5356 3352
rect 5408 3340 5414 3392
rect 5442 3340 5448 3392
rect 5500 3380 5506 3392
rect 5721 3383 5779 3389
rect 5721 3380 5733 3383
rect 5500 3352 5733 3380
rect 5500 3340 5506 3352
rect 5721 3349 5733 3352
rect 5767 3349 5779 3383
rect 6638 3380 6644 3392
rect 6599 3352 6644 3380
rect 5721 3343 5779 3349
rect 6638 3340 6644 3352
rect 6696 3340 6702 3392
rect 7282 3380 7288 3392
rect 7243 3352 7288 3380
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 7558 3380 7564 3392
rect 7519 3352 7564 3380
rect 7558 3340 7564 3352
rect 7616 3340 7622 3392
rect 7742 3380 7748 3392
rect 7703 3352 7748 3380
rect 7742 3340 7748 3352
rect 7800 3340 7806 3392
rect 8021 3383 8079 3389
rect 8021 3349 8033 3383
rect 8067 3380 8079 3383
rect 8294 3380 8300 3392
rect 8067 3352 8300 3380
rect 8067 3349 8079 3352
rect 8021 3343 8079 3349
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 9674 3340 9680 3392
rect 9732 3380 9738 3392
rect 10137 3383 10195 3389
rect 10137 3380 10149 3383
rect 9732 3352 10149 3380
rect 9732 3340 9738 3352
rect 10137 3349 10149 3352
rect 10183 3349 10195 3383
rect 10137 3343 10195 3349
rect 10226 3340 10232 3392
rect 10284 3380 10290 3392
rect 12176 3389 12204 3420
rect 13265 3417 13277 3420
rect 13311 3417 13323 3451
rect 13464 3448 13492 3488
rect 13817 3485 13829 3488
rect 13863 3485 13875 3519
rect 13817 3479 13875 3485
rect 21269 3519 21327 3525
rect 21269 3485 21281 3519
rect 21315 3516 21327 3519
rect 21545 3519 21603 3525
rect 21545 3516 21557 3519
rect 21315 3488 21557 3516
rect 21315 3485 21327 3488
rect 21269 3479 21327 3485
rect 21545 3485 21557 3488
rect 21591 3516 21603 3519
rect 22462 3516 22468 3528
rect 21591 3488 22468 3516
rect 21591 3485 21603 3488
rect 21545 3479 21603 3485
rect 22462 3476 22468 3488
rect 22520 3476 22526 3528
rect 13265 3411 13323 3417
rect 13372 3420 13492 3448
rect 10965 3383 11023 3389
rect 10965 3380 10977 3383
rect 10284 3352 10977 3380
rect 10284 3340 10290 3352
rect 10965 3349 10977 3352
rect 11011 3349 11023 3383
rect 10965 3343 11023 3349
rect 11333 3383 11391 3389
rect 11333 3349 11345 3383
rect 11379 3380 11391 3383
rect 11701 3383 11759 3389
rect 11701 3380 11713 3383
rect 11379 3352 11713 3380
rect 11379 3349 11391 3352
rect 11333 3343 11391 3349
rect 11701 3349 11713 3352
rect 11747 3349 11759 3383
rect 11701 3343 11759 3349
rect 12161 3383 12219 3389
rect 12161 3349 12173 3383
rect 12207 3349 12219 3383
rect 12161 3343 12219 3349
rect 12986 3340 12992 3392
rect 13044 3380 13050 3392
rect 13372 3380 13400 3420
rect 13630 3408 13636 3460
rect 13688 3448 13694 3460
rect 14277 3451 14335 3457
rect 14277 3448 14289 3451
rect 13688 3420 14289 3448
rect 13688 3408 13694 3420
rect 14277 3417 14289 3420
rect 14323 3417 14335 3451
rect 14277 3411 14335 3417
rect 13722 3380 13728 3392
rect 13044 3352 13400 3380
rect 13683 3352 13728 3380
rect 13044 3340 13050 3352
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 2130 3136 2136 3188
rect 2188 3176 2194 3188
rect 2774 3176 2780 3188
rect 2188 3148 2780 3176
rect 2188 3136 2194 3148
rect 2774 3136 2780 3148
rect 2832 3136 2838 3188
rect 2869 3179 2927 3185
rect 2869 3145 2881 3179
rect 2915 3176 2927 3179
rect 4062 3176 4068 3188
rect 2915 3148 4068 3176
rect 2915 3145 2927 3148
rect 2869 3139 2927 3145
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 4246 3176 4252 3188
rect 4207 3148 4252 3176
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 4338 3136 4344 3188
rect 4396 3176 4402 3188
rect 4614 3176 4620 3188
rect 4396 3148 4620 3176
rect 4396 3136 4402 3148
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 4908 3148 6592 3176
rect 2409 3111 2467 3117
rect 2409 3077 2421 3111
rect 2455 3108 2467 3111
rect 3789 3111 3847 3117
rect 3789 3108 3801 3111
rect 2455 3080 2820 3108
rect 2455 3077 2467 3080
rect 2409 3071 2467 3077
rect 2792 3052 2820 3080
rect 2884 3080 3801 3108
rect 1762 3000 1768 3052
rect 1820 3040 1826 3052
rect 2682 3040 2688 3052
rect 1820 3012 2688 3040
rect 1820 3000 1826 3012
rect 2682 3000 2688 3012
rect 2740 3000 2746 3052
rect 2774 3000 2780 3052
rect 2832 3000 2838 3052
rect 1949 2975 2007 2981
rect 1949 2941 1961 2975
rect 1995 2972 2007 2975
rect 2038 2972 2044 2984
rect 1995 2944 2044 2972
rect 1995 2941 2007 2944
rect 1949 2935 2007 2941
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 2130 2932 2136 2984
rect 2188 2972 2194 2984
rect 2225 2975 2283 2981
rect 2225 2972 2237 2975
rect 2188 2944 2237 2972
rect 2188 2932 2194 2944
rect 2225 2941 2237 2944
rect 2271 2941 2283 2975
rect 2225 2935 2283 2941
rect 2314 2932 2320 2984
rect 2372 2972 2378 2984
rect 2884 2972 2912 3080
rect 3789 3077 3801 3080
rect 3835 3077 3847 3111
rect 4908 3108 4936 3148
rect 5074 3108 5080 3120
rect 3789 3071 3847 3077
rect 4080 3080 4936 3108
rect 5000 3080 5080 3108
rect 2961 3043 3019 3049
rect 2961 3009 2973 3043
rect 3007 3040 3019 3043
rect 3237 3043 3295 3049
rect 3237 3040 3249 3043
rect 3007 3012 3249 3040
rect 3007 3009 3019 3012
rect 2961 3003 3019 3009
rect 3237 3009 3249 3012
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 2372 2944 2912 2972
rect 2372 2932 2378 2944
rect 842 2864 848 2916
rect 900 2904 906 2916
rect 2976 2904 3004 3003
rect 3421 2907 3479 2913
rect 3421 2904 3433 2907
rect 900 2876 3004 2904
rect 3068 2876 3433 2904
rect 900 2864 906 2876
rect 2498 2836 2504 2848
rect 2459 2808 2504 2836
rect 2498 2796 2504 2808
rect 2556 2796 2562 2848
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 3068 2836 3096 2876
rect 3421 2873 3433 2876
rect 3467 2873 3479 2907
rect 3421 2867 3479 2873
rect 3697 2907 3755 2913
rect 3697 2873 3709 2907
rect 3743 2904 3755 2907
rect 3878 2904 3884 2916
rect 3743 2876 3884 2904
rect 3743 2873 3755 2876
rect 3697 2867 3755 2873
rect 3878 2864 3884 2876
rect 3936 2864 3942 2916
rect 2832 2808 3096 2836
rect 3145 2839 3203 2845
rect 2832 2796 2838 2808
rect 3145 2805 3157 2839
rect 3191 2836 3203 2839
rect 4080 2836 4108 3080
rect 4706 2972 4712 2984
rect 4667 2944 4712 2972
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 4893 2975 4951 2981
rect 4893 2941 4905 2975
rect 4939 2972 4951 2975
rect 5000 2972 5028 3080
rect 5074 3068 5080 3080
rect 5132 3068 5138 3120
rect 6564 3040 6592 3148
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 7377 3179 7435 3185
rect 7377 3176 7389 3179
rect 6696 3148 7389 3176
rect 6696 3136 6702 3148
rect 7377 3145 7389 3148
rect 7423 3145 7435 3179
rect 7377 3139 7435 3145
rect 7650 3136 7656 3188
rect 7708 3176 7714 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7708 3148 7757 3176
rect 7708 3136 7714 3148
rect 7745 3145 7757 3148
rect 7791 3176 7803 3179
rect 8202 3176 8208 3188
rect 7791 3148 8208 3176
rect 7791 3145 7803 3148
rect 7745 3139 7803 3145
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 8478 3176 8484 3188
rect 8439 3148 8484 3176
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 8938 3176 8944 3188
rect 8899 3148 8944 3176
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 10045 3179 10103 3185
rect 9456 3148 9996 3176
rect 9456 3136 9462 3148
rect 7006 3068 7012 3120
rect 7064 3108 7070 3120
rect 8294 3108 8300 3120
rect 7064 3080 8064 3108
rect 8207 3080 8300 3108
rect 7064 3068 7070 3080
rect 7837 3043 7895 3049
rect 7837 3040 7849 3043
rect 6564 3012 7849 3040
rect 7837 3009 7849 3012
rect 7883 3009 7895 3043
rect 7837 3003 7895 3009
rect 4939 2944 5028 2972
rect 5077 2975 5135 2981
rect 4939 2941 4951 2944
rect 4893 2935 4951 2941
rect 5077 2941 5089 2975
rect 5123 2941 5135 2975
rect 5077 2935 5135 2941
rect 4157 2907 4215 2913
rect 4157 2873 4169 2907
rect 4203 2904 4215 2907
rect 4982 2904 4988 2916
rect 4203 2876 4988 2904
rect 4203 2873 4215 2876
rect 4157 2867 4215 2873
rect 4982 2864 4988 2876
rect 5040 2904 5046 2916
rect 5092 2904 5120 2935
rect 5258 2932 5264 2984
rect 5316 2972 5322 2984
rect 5353 2975 5411 2981
rect 5353 2972 5365 2975
rect 5316 2944 5365 2972
rect 5316 2932 5322 2944
rect 5353 2941 5365 2944
rect 5399 2941 5411 2975
rect 5353 2935 5411 2941
rect 6181 2975 6239 2981
rect 6181 2941 6193 2975
rect 6227 2972 6239 2975
rect 6457 2975 6515 2981
rect 6457 2972 6469 2975
rect 6227 2944 6469 2972
rect 6227 2941 6239 2944
rect 6181 2935 6239 2941
rect 6457 2941 6469 2944
rect 6503 2972 6515 2975
rect 6546 2972 6552 2984
rect 6503 2944 6552 2972
rect 6503 2941 6515 2944
rect 6457 2935 6515 2941
rect 6546 2932 6552 2944
rect 6604 2932 6610 2984
rect 6733 2975 6791 2981
rect 6733 2941 6745 2975
rect 6779 2972 6791 2975
rect 7466 2972 7472 2984
rect 6779 2944 7472 2972
rect 6779 2941 6791 2944
rect 6733 2935 6791 2941
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 5040 2876 5120 2904
rect 5040 2864 5046 2876
rect 3191 2808 4108 2836
rect 3191 2805 3203 2808
rect 3145 2799 3203 2805
rect 4246 2796 4252 2848
rect 4304 2836 4310 2848
rect 5350 2836 5356 2848
rect 4304 2808 5356 2836
rect 4304 2796 4310 2808
rect 5350 2796 5356 2808
rect 5408 2796 5414 2848
rect 7852 2836 7880 3003
rect 8036 2981 8064 3080
rect 8220 3049 8248 3080
rect 8294 3068 8300 3080
rect 8352 3108 8358 3120
rect 9122 3108 9128 3120
rect 8352 3080 9128 3108
rect 8352 3068 8358 3080
rect 9122 3068 9128 3080
rect 9180 3068 9186 3120
rect 9582 3068 9588 3120
rect 9640 3068 9646 3120
rect 9968 3108 9996 3148
rect 10045 3145 10057 3179
rect 10091 3176 10103 3179
rect 10226 3176 10232 3188
rect 10091 3148 10232 3176
rect 10091 3145 10103 3148
rect 10045 3139 10103 3145
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 11882 3136 11888 3188
rect 11940 3176 11946 3188
rect 12437 3179 12495 3185
rect 12437 3176 12449 3179
rect 11940 3148 12449 3176
rect 11940 3136 11946 3148
rect 12437 3145 12449 3148
rect 12483 3145 12495 3179
rect 12437 3139 12495 3145
rect 12618 3136 12624 3188
rect 12676 3176 12682 3188
rect 12897 3179 12955 3185
rect 12897 3176 12909 3179
rect 12676 3148 12909 3176
rect 12676 3136 12682 3148
rect 12897 3145 12909 3148
rect 12943 3176 12955 3179
rect 14829 3179 14887 3185
rect 12943 3148 13584 3176
rect 12943 3145 12955 3148
rect 12897 3139 12955 3145
rect 11241 3111 11299 3117
rect 11241 3108 11253 3111
rect 9968 3080 11253 3108
rect 11241 3077 11253 3080
rect 11287 3077 11299 3111
rect 11241 3071 11299 3077
rect 12805 3111 12863 3117
rect 12805 3077 12817 3111
rect 12851 3108 12863 3111
rect 13078 3108 13084 3120
rect 12851 3080 13084 3108
rect 12851 3077 12863 3080
rect 12805 3071 12863 3077
rect 8205 3043 8263 3049
rect 8205 3009 8217 3043
rect 8251 3009 8263 3043
rect 8205 3003 8263 3009
rect 8570 3000 8576 3052
rect 8628 3040 8634 3052
rect 8849 3043 8907 3049
rect 8849 3040 8861 3043
rect 8628 3012 8861 3040
rect 8628 3000 8634 3012
rect 8849 3009 8861 3012
rect 8895 3009 8907 3043
rect 9600 3040 9628 3068
rect 8849 3003 8907 3009
rect 9140 3012 9628 3040
rect 9677 3043 9735 3049
rect 9140 2981 9168 3012
rect 9677 3009 9689 3043
rect 9723 3040 9735 3043
rect 9766 3040 9772 3052
rect 9723 3012 9772 3040
rect 9723 3009 9735 3012
rect 9677 3003 9735 3009
rect 9766 3000 9772 3012
rect 9824 3000 9830 3052
rect 9950 3000 9956 3052
rect 10008 3040 10014 3052
rect 10137 3043 10195 3049
rect 10137 3040 10149 3043
rect 10008 3012 10149 3040
rect 10008 3000 10014 3012
rect 10137 3009 10149 3012
rect 10183 3009 10195 3043
rect 10410 3040 10416 3052
rect 10371 3012 10416 3040
rect 10137 3003 10195 3009
rect 10410 3000 10416 3012
rect 10468 3000 10474 3052
rect 8021 2975 8079 2981
rect 8021 2941 8033 2975
rect 8067 2972 8079 2975
rect 9125 2975 9183 2981
rect 8067 2944 8892 2972
rect 8067 2941 8079 2944
rect 8021 2935 8079 2941
rect 8389 2907 8447 2913
rect 8389 2873 8401 2907
rect 8435 2904 8447 2907
rect 8754 2904 8760 2916
rect 8435 2876 8760 2904
rect 8435 2873 8447 2876
rect 8389 2867 8447 2873
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 8864 2904 8892 2944
rect 9125 2941 9137 2975
rect 9171 2941 9183 2975
rect 9398 2972 9404 2984
rect 9359 2944 9404 2972
rect 9125 2935 9183 2941
rect 9398 2932 9404 2944
rect 9456 2932 9462 2984
rect 9585 2975 9643 2981
rect 9585 2941 9597 2975
rect 9631 2972 9643 2975
rect 10042 2972 10048 2984
rect 9631 2944 10048 2972
rect 9631 2941 9643 2944
rect 9585 2935 9643 2941
rect 10042 2932 10048 2944
rect 10100 2932 10106 2984
rect 11256 2972 11284 3071
rect 13078 3068 13084 3080
rect 13136 3068 13142 3120
rect 13556 3108 13584 3148
rect 14829 3145 14841 3179
rect 14875 3176 14887 3179
rect 16114 3176 16120 3188
rect 14875 3148 16120 3176
rect 14875 3145 14887 3148
rect 14829 3139 14887 3145
rect 16114 3136 16120 3148
rect 16172 3136 16178 3188
rect 17310 3136 17316 3188
rect 17368 3176 17374 3188
rect 17681 3179 17739 3185
rect 17681 3176 17693 3179
rect 17368 3148 17693 3176
rect 17368 3136 17374 3148
rect 17681 3145 17693 3148
rect 17727 3145 17739 3179
rect 17954 3176 17960 3188
rect 17915 3148 17960 3176
rect 17681 3139 17739 3145
rect 15197 3111 15255 3117
rect 15197 3108 15209 3111
rect 13556 3080 15209 3108
rect 11517 3043 11575 3049
rect 11517 3009 11529 3043
rect 11563 3040 11575 3043
rect 11698 3040 11704 3052
rect 11563 3012 11704 3040
rect 11563 3009 11575 3012
rect 11517 3003 11575 3009
rect 11698 3000 11704 3012
rect 11756 3000 11762 3052
rect 11790 3000 11796 3052
rect 11848 3040 11854 3052
rect 13446 3040 13452 3052
rect 11848 3012 11893 3040
rect 13407 3012 13452 3040
rect 11848 3000 11854 3012
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 13538 3000 13544 3052
rect 13596 3040 13602 3052
rect 13596 3012 13641 3040
rect 13596 3000 13602 3012
rect 13722 3000 13728 3052
rect 13780 3040 13786 3052
rect 13817 3043 13875 3049
rect 13817 3040 13829 3043
rect 13780 3012 13829 3040
rect 13780 3000 13786 3012
rect 13817 3009 13829 3012
rect 13863 3009 13875 3043
rect 14090 3040 14096 3052
rect 14051 3012 14096 3040
rect 13817 3003 13875 3009
rect 14090 3000 14096 3012
rect 14148 3000 14154 3052
rect 14660 3049 14688 3080
rect 15197 3077 15209 3080
rect 15243 3077 15255 3111
rect 15930 3108 15936 3120
rect 15891 3080 15936 3108
rect 15197 3071 15255 3077
rect 15930 3068 15936 3080
rect 15988 3068 15994 3120
rect 17126 3108 17132 3120
rect 16684 3080 17132 3108
rect 14369 3043 14427 3049
rect 14369 3009 14381 3043
rect 14415 3009 14427 3043
rect 14369 3003 14427 3009
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3009 14703 3043
rect 14918 3040 14924 3052
rect 14879 3012 14924 3040
rect 14645 3003 14703 3009
rect 12986 2972 12992 2984
rect 11256 2944 12992 2972
rect 12986 2932 12992 2944
rect 13044 2932 13050 2984
rect 14384 2972 14412 3003
rect 14918 3000 14924 3012
rect 14976 3000 14982 3052
rect 15102 3000 15108 3052
rect 15160 3040 15166 3052
rect 15473 3043 15531 3049
rect 15473 3040 15485 3043
rect 15160 3012 15485 3040
rect 15160 3000 15166 3012
rect 15473 3009 15485 3012
rect 15519 3040 15531 3043
rect 15657 3043 15715 3049
rect 15657 3040 15669 3043
rect 15519 3012 15669 3040
rect 15519 3009 15531 3012
rect 15473 3003 15531 3009
rect 15657 3009 15669 3012
rect 15703 3009 15715 3043
rect 15948 3040 15976 3068
rect 16684 3049 16712 3080
rect 17126 3068 17132 3080
rect 17184 3108 17190 3120
rect 17221 3111 17279 3117
rect 17221 3108 17233 3111
rect 17184 3080 17233 3108
rect 17184 3068 17190 3080
rect 17221 3077 17233 3080
rect 17267 3077 17279 3111
rect 17221 3071 17279 3077
rect 16117 3043 16175 3049
rect 16117 3040 16129 3043
rect 15948 3012 16129 3040
rect 15657 3003 15715 3009
rect 16117 3009 16129 3012
rect 16163 3009 16175 3043
rect 16117 3003 16175 3009
rect 16669 3043 16727 3049
rect 16669 3009 16681 3043
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 16945 3043 17003 3049
rect 16945 3009 16957 3043
rect 16991 3040 17003 3043
rect 17034 3040 17040 3052
rect 16991 3012 17040 3040
rect 16991 3009 17003 3012
rect 16945 3003 17003 3009
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 14016 2944 14412 2972
rect 17696 2972 17724 3139
rect 17954 3136 17960 3148
rect 18012 3136 18018 3188
rect 18233 3179 18291 3185
rect 18233 3145 18245 3179
rect 18279 3145 18291 3179
rect 18233 3139 18291 3145
rect 19061 3179 19119 3185
rect 19061 3145 19073 3179
rect 19107 3176 19119 3179
rect 19150 3176 19156 3188
rect 19107 3148 19156 3176
rect 19107 3145 19119 3148
rect 19061 3139 19119 3145
rect 17972 3040 18000 3136
rect 18248 3108 18276 3139
rect 19150 3136 19156 3148
rect 19208 3136 19214 3188
rect 19426 3136 19432 3188
rect 19484 3136 19490 3188
rect 19702 3136 19708 3188
rect 19760 3176 19766 3188
rect 19760 3148 21312 3176
rect 19760 3136 19766 3148
rect 19444 3108 19472 3136
rect 18248 3080 19196 3108
rect 19444 3080 20944 3108
rect 18049 3043 18107 3049
rect 18049 3040 18061 3043
rect 17972 3012 18061 3040
rect 18049 3009 18061 3012
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 18509 3043 18567 3049
rect 18509 3009 18521 3043
rect 18555 3009 18567 3043
rect 18509 3003 18567 3009
rect 18601 3043 18659 3049
rect 18601 3009 18613 3043
rect 18647 3009 18659 3043
rect 18874 3040 18880 3052
rect 18835 3012 18880 3040
rect 18601 3003 18659 3009
rect 18524 2972 18552 3003
rect 17696 2944 18552 2972
rect 14016 2913 14044 2944
rect 11057 2907 11115 2913
rect 11057 2904 11069 2907
rect 8864 2876 11069 2904
rect 11057 2873 11069 2876
rect 11103 2873 11115 2907
rect 11057 2867 11115 2873
rect 14001 2907 14059 2913
rect 14001 2873 14013 2907
rect 14047 2873 14059 2907
rect 14001 2867 14059 2873
rect 14277 2907 14335 2913
rect 14277 2873 14289 2907
rect 14323 2904 14335 2907
rect 14734 2904 14740 2916
rect 14323 2876 14740 2904
rect 14323 2873 14335 2876
rect 14277 2867 14335 2873
rect 14734 2864 14740 2876
rect 14792 2864 14798 2916
rect 15105 2907 15163 2913
rect 15105 2873 15117 2907
rect 15151 2904 15163 2907
rect 15286 2904 15292 2916
rect 15151 2876 15292 2904
rect 15151 2873 15163 2876
rect 15105 2867 15163 2873
rect 15286 2864 15292 2876
rect 15344 2864 15350 2916
rect 15841 2907 15899 2913
rect 15841 2873 15853 2907
rect 15887 2904 15899 2907
rect 16758 2904 16764 2916
rect 15887 2876 16764 2904
rect 15887 2873 15899 2876
rect 15841 2867 15899 2873
rect 16758 2864 16764 2876
rect 16816 2864 16822 2916
rect 16853 2907 16911 2913
rect 16853 2873 16865 2907
rect 16899 2904 16911 2907
rect 17494 2904 17500 2916
rect 16899 2876 17500 2904
rect 16899 2873 16911 2876
rect 16853 2867 16911 2873
rect 17494 2864 17500 2876
rect 17552 2864 17558 2916
rect 17862 2864 17868 2916
rect 17920 2904 17926 2916
rect 18616 2904 18644 3003
rect 18874 3000 18880 3012
rect 18932 3000 18938 3052
rect 19168 2972 19196 3080
rect 19334 3040 19340 3052
rect 19295 3012 19340 3040
rect 19334 3000 19340 3012
rect 19392 3040 19398 3052
rect 19613 3043 19671 3049
rect 19613 3040 19625 3043
rect 19392 3012 19625 3040
rect 19392 3000 19398 3012
rect 19613 3009 19625 3012
rect 19659 3009 19671 3043
rect 19886 3040 19892 3052
rect 19847 3012 19892 3040
rect 19613 3003 19671 3009
rect 19886 3000 19892 3012
rect 19944 3000 19950 3052
rect 20346 3040 20352 3052
rect 20307 3012 20352 3040
rect 20346 3000 20352 3012
rect 20404 3000 20410 3052
rect 20714 3040 20720 3052
rect 20675 3012 20720 3040
rect 20714 3000 20720 3012
rect 20772 3000 20778 3052
rect 20916 3049 20944 3080
rect 21284 3049 21312 3148
rect 20901 3043 20959 3049
rect 20901 3009 20913 3043
rect 20947 3009 20959 3043
rect 20901 3003 20959 3009
rect 21269 3043 21327 3049
rect 21269 3009 21281 3043
rect 21315 3009 21327 3043
rect 21269 3003 21327 3009
rect 19702 2972 19708 2984
rect 19168 2944 19708 2972
rect 19702 2932 19708 2944
rect 19760 2932 19766 2984
rect 21174 2972 21180 2984
rect 19812 2944 21180 2972
rect 17920 2876 18644 2904
rect 17920 2864 17926 2876
rect 18690 2864 18696 2916
rect 18748 2904 18754 2916
rect 19153 2907 19211 2913
rect 19153 2904 19165 2907
rect 18748 2876 19165 2904
rect 18748 2864 18754 2876
rect 19153 2873 19165 2876
rect 19199 2873 19211 2907
rect 19153 2867 19211 2873
rect 19242 2864 19248 2916
rect 19300 2904 19306 2916
rect 19429 2907 19487 2913
rect 19429 2904 19441 2907
rect 19300 2876 19441 2904
rect 19300 2864 19306 2876
rect 19429 2873 19441 2876
rect 19475 2873 19487 2907
rect 19429 2867 19487 2873
rect 9674 2836 9680 2848
rect 7852 2808 9680 2836
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 13265 2839 13323 2845
rect 13265 2805 13277 2839
rect 13311 2836 13323 2839
rect 13354 2836 13360 2848
rect 13311 2808 13360 2836
rect 13311 2805 13323 2808
rect 13265 2799 13323 2805
rect 13354 2796 13360 2808
rect 13412 2796 13418 2848
rect 13725 2839 13783 2845
rect 13725 2805 13737 2839
rect 13771 2836 13783 2839
rect 13814 2836 13820 2848
rect 13771 2808 13820 2836
rect 13771 2805 13783 2808
rect 13725 2799 13783 2805
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 14458 2796 14464 2848
rect 14516 2836 14522 2848
rect 14553 2839 14611 2845
rect 14553 2836 14565 2839
rect 14516 2808 14565 2836
rect 14516 2796 14522 2808
rect 14553 2805 14565 2808
rect 14599 2805 14611 2839
rect 14553 2799 14611 2805
rect 16301 2839 16359 2845
rect 16301 2805 16313 2839
rect 16347 2836 16359 2839
rect 16666 2836 16672 2848
rect 16347 2808 16672 2836
rect 16347 2805 16359 2808
rect 16301 2799 16359 2805
rect 16666 2796 16672 2808
rect 16724 2796 16730 2848
rect 17126 2836 17132 2848
rect 17087 2808 17132 2836
rect 17126 2796 17132 2808
rect 17184 2796 17190 2848
rect 18322 2796 18328 2848
rect 18380 2836 18386 2848
rect 18785 2839 18843 2845
rect 18380 2808 18425 2836
rect 18380 2796 18386 2808
rect 18785 2805 18797 2839
rect 18831 2836 18843 2839
rect 19812 2836 19840 2944
rect 21174 2932 21180 2944
rect 21232 2932 21238 2984
rect 19886 2864 19892 2916
rect 19944 2904 19950 2916
rect 20165 2907 20223 2913
rect 20165 2904 20177 2907
rect 19944 2876 20177 2904
rect 19944 2864 19950 2876
rect 20165 2873 20177 2876
rect 20211 2873 20223 2907
rect 20714 2904 20720 2916
rect 20165 2867 20223 2873
rect 20364 2876 20720 2904
rect 18831 2808 19840 2836
rect 20073 2839 20131 2845
rect 18831 2805 18843 2808
rect 18785 2799 18843 2805
rect 20073 2805 20085 2839
rect 20119 2836 20131 2839
rect 20364 2836 20392 2876
rect 20714 2864 20720 2876
rect 20772 2864 20778 2916
rect 21085 2907 21143 2913
rect 21085 2873 21097 2907
rect 21131 2904 21143 2907
rect 22094 2904 22100 2916
rect 21131 2876 22100 2904
rect 21131 2873 21143 2876
rect 21085 2867 21143 2873
rect 22094 2864 22100 2876
rect 22152 2864 22158 2916
rect 20119 2808 20392 2836
rect 20119 2805 20131 2808
rect 20073 2799 20131 2805
rect 20438 2796 20444 2848
rect 20496 2836 20502 2848
rect 20533 2839 20591 2845
rect 20533 2836 20545 2839
rect 20496 2808 20545 2836
rect 20496 2796 20502 2808
rect 20533 2805 20545 2808
rect 20579 2805 20591 2839
rect 20533 2799 20591 2805
rect 21453 2839 21511 2845
rect 21453 2805 21465 2839
rect 21499 2836 21511 2839
rect 21542 2836 21548 2848
rect 21499 2808 21548 2836
rect 21499 2805 21511 2808
rect 21453 2799 21511 2805
rect 21542 2796 21548 2808
rect 21600 2796 21606 2848
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 2222 2632 2228 2644
rect 1964 2604 2228 2632
rect 1964 2505 1992 2604
rect 2222 2592 2228 2604
rect 2280 2592 2286 2644
rect 2961 2635 3019 2641
rect 2961 2601 2973 2635
rect 3007 2632 3019 2635
rect 3973 2635 4031 2641
rect 3007 2604 3924 2632
rect 3007 2601 3019 2604
rect 2961 2595 3019 2601
rect 3418 2564 3424 2576
rect 2240 2536 3424 2564
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2465 2007 2499
rect 1949 2459 2007 2465
rect 2240 2440 2268 2536
rect 3418 2524 3424 2536
rect 3476 2524 3482 2576
rect 3896 2564 3924 2604
rect 3973 2601 3985 2635
rect 4019 2632 4031 2635
rect 4246 2632 4252 2644
rect 4019 2604 4252 2632
rect 4019 2601 4031 2604
rect 3973 2595 4031 2601
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 4798 2632 4804 2644
rect 4759 2604 4804 2632
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 4890 2592 4896 2644
rect 4948 2632 4954 2644
rect 5261 2635 5319 2641
rect 5261 2632 5273 2635
rect 4948 2604 5273 2632
rect 4948 2592 4954 2604
rect 5261 2601 5273 2604
rect 5307 2601 5319 2635
rect 5261 2595 5319 2601
rect 5350 2592 5356 2644
rect 5408 2632 5414 2644
rect 8570 2632 8576 2644
rect 5408 2604 8576 2632
rect 5408 2592 5414 2604
rect 8570 2592 8576 2604
rect 8628 2632 8634 2644
rect 9490 2632 9496 2644
rect 8628 2604 9496 2632
rect 8628 2592 8634 2604
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 10137 2635 10195 2641
rect 10137 2601 10149 2635
rect 10183 2632 10195 2635
rect 10413 2635 10471 2641
rect 10183 2604 10364 2632
rect 10183 2601 10195 2604
rect 10137 2595 10195 2601
rect 4341 2567 4399 2573
rect 3896 2536 4292 2564
rect 3053 2499 3111 2505
rect 3053 2465 3065 2499
rect 3099 2496 3111 2499
rect 4264 2496 4292 2536
rect 4341 2533 4353 2567
rect 4387 2564 4399 2567
rect 5534 2564 5540 2576
rect 4387 2536 5540 2564
rect 4387 2533 4399 2536
rect 4341 2527 4399 2533
rect 5534 2524 5540 2536
rect 5592 2524 5598 2576
rect 10336 2564 10364 2604
rect 10413 2601 10425 2635
rect 10459 2632 10471 2635
rect 11146 2632 11152 2644
rect 10459 2604 11152 2632
rect 10459 2601 10471 2604
rect 10413 2595 10471 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 12115 2635 12173 2641
rect 12115 2601 12127 2635
rect 12161 2632 12173 2635
rect 12434 2632 12440 2644
rect 12161 2604 12440 2632
rect 12161 2601 12173 2604
rect 12115 2595 12173 2601
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 13722 2592 13728 2644
rect 13780 2632 13786 2644
rect 14277 2635 14335 2641
rect 14277 2632 14289 2635
rect 13780 2604 14289 2632
rect 13780 2592 13786 2604
rect 14277 2601 14289 2604
rect 14323 2601 14335 2635
rect 14277 2595 14335 2601
rect 16666 2592 16672 2644
rect 16724 2632 16730 2644
rect 16724 2604 20392 2632
rect 16724 2592 16730 2604
rect 9508 2536 10180 2564
rect 10336 2536 13400 2564
rect 4706 2496 4712 2508
rect 3099 2468 4108 2496
rect 4264 2468 4712 2496
rect 3099 2465 3111 2468
rect 3053 2459 3111 2465
rect 4080 2440 4108 2468
rect 4706 2456 4712 2468
rect 4764 2496 4770 2508
rect 5350 2496 5356 2508
rect 4764 2468 5356 2496
rect 4764 2456 4770 2468
rect 5350 2456 5356 2468
rect 5408 2456 5414 2508
rect 5626 2456 5632 2508
rect 5684 2496 5690 2508
rect 5905 2499 5963 2505
rect 5905 2496 5917 2499
rect 5684 2468 5917 2496
rect 5684 2456 5690 2468
rect 5905 2465 5917 2468
rect 5951 2465 5963 2499
rect 5905 2459 5963 2465
rect 7193 2499 7251 2505
rect 7193 2465 7205 2499
rect 7239 2496 7251 2499
rect 9214 2496 9220 2508
rect 7239 2468 9220 2496
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 9214 2456 9220 2468
rect 9272 2456 9278 2508
rect 9508 2505 9536 2536
rect 10152 2508 10180 2536
rect 9493 2499 9551 2505
rect 9493 2465 9505 2499
rect 9539 2465 9551 2499
rect 9674 2496 9680 2508
rect 9635 2468 9680 2496
rect 9493 2459 9551 2465
rect 9674 2456 9680 2468
rect 9732 2456 9738 2508
rect 10134 2456 10140 2508
rect 10192 2456 10198 2508
rect 10778 2456 10784 2508
rect 10836 2496 10842 2508
rect 11333 2499 11391 2505
rect 11333 2496 11345 2499
rect 10836 2468 11345 2496
rect 10836 2456 10842 2468
rect 11333 2465 11345 2468
rect 11379 2465 11391 2499
rect 12434 2496 12440 2508
rect 12347 2468 12440 2496
rect 11333 2459 11391 2465
rect 12434 2456 12440 2468
rect 12492 2496 12498 2508
rect 12894 2496 12900 2508
rect 12492 2468 12900 2496
rect 12492 2456 12498 2468
rect 12894 2456 12900 2468
rect 12952 2456 12958 2508
rect 13372 2496 13400 2536
rect 14182 2524 14188 2576
rect 14240 2564 14246 2576
rect 14645 2567 14703 2573
rect 14645 2564 14657 2567
rect 14240 2536 14657 2564
rect 14240 2524 14246 2536
rect 14645 2533 14657 2536
rect 14691 2533 14703 2567
rect 14645 2527 14703 2533
rect 19242 2524 19248 2576
rect 19300 2564 19306 2576
rect 19705 2567 19763 2573
rect 19705 2564 19717 2567
rect 19300 2536 19717 2564
rect 19300 2524 19306 2536
rect 19705 2533 19717 2536
rect 19751 2533 19763 2567
rect 19705 2527 19763 2533
rect 17678 2496 17684 2508
rect 13372 2468 17684 2496
rect 17678 2456 17684 2468
rect 17736 2456 17742 2508
rect 20254 2496 20260 2508
rect 19536 2468 20260 2496
rect 2222 2428 2228 2440
rect 2183 2400 2228 2428
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 2314 2388 2320 2440
rect 2372 2428 2378 2440
rect 2777 2431 2835 2437
rect 2372 2400 2417 2428
rect 2372 2388 2378 2400
rect 2777 2397 2789 2431
rect 2823 2428 2835 2431
rect 2866 2428 2872 2440
rect 2823 2400 2872 2428
rect 2823 2397 2835 2400
rect 2777 2391 2835 2397
rect 2866 2388 2872 2400
rect 2924 2388 2930 2440
rect 3142 2388 3148 2440
rect 3200 2428 3206 2440
rect 3237 2431 3295 2437
rect 3237 2428 3249 2431
rect 3200 2400 3249 2428
rect 3200 2388 3206 2400
rect 3237 2397 3249 2400
rect 3283 2397 3295 2431
rect 3237 2391 3295 2397
rect 3789 2431 3847 2437
rect 3789 2397 3801 2431
rect 3835 2428 3847 2431
rect 3878 2428 3884 2440
rect 3835 2400 3884 2428
rect 3835 2397 3847 2400
rect 3789 2391 3847 2397
rect 3878 2388 3884 2400
rect 3936 2388 3942 2440
rect 4062 2388 4068 2440
rect 4120 2428 4126 2440
rect 4157 2431 4215 2437
rect 4157 2428 4169 2431
rect 4120 2400 4169 2428
rect 4120 2388 4126 2400
rect 4157 2397 4169 2400
rect 4203 2397 4215 2431
rect 4157 2391 4215 2397
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4580 2400 4629 2428
rect 4580 2388 4586 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 5077 2431 5135 2437
rect 5077 2397 5089 2431
rect 5123 2428 5135 2431
rect 5442 2428 5448 2440
rect 5123 2400 5448 2428
rect 5123 2397 5135 2400
rect 5077 2391 5135 2397
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 6181 2431 6239 2437
rect 6181 2428 6193 2431
rect 5920 2400 6193 2428
rect 2685 2363 2743 2369
rect 2685 2329 2697 2363
rect 2731 2360 2743 2363
rect 3160 2360 3188 2388
rect 2731 2332 3188 2360
rect 3605 2363 3663 2369
rect 2731 2329 2743 2332
rect 2685 2323 2743 2329
rect 3605 2329 3617 2363
rect 3651 2360 3663 2363
rect 4540 2360 4568 2388
rect 5920 2372 5948 2400
rect 6181 2397 6193 2400
rect 6227 2397 6239 2431
rect 6822 2428 6828 2440
rect 6181 2391 6239 2397
rect 6288 2400 6828 2428
rect 5902 2360 5908 2372
rect 3651 2332 4568 2360
rect 4816 2332 5908 2360
rect 3651 2329 3663 2332
rect 3605 2323 3663 2329
rect 2498 2292 2504 2304
rect 2459 2264 2504 2292
rect 2498 2252 2504 2264
rect 2556 2252 2562 2304
rect 3421 2295 3479 2301
rect 3421 2261 3433 2295
rect 3467 2292 3479 2295
rect 4246 2292 4252 2304
rect 3467 2264 4252 2292
rect 3467 2261 3479 2264
rect 3421 2255 3479 2261
rect 4246 2252 4252 2264
rect 4304 2252 4310 2304
rect 4525 2295 4583 2301
rect 4525 2261 4537 2295
rect 4571 2292 4583 2295
rect 4816 2292 4844 2332
rect 5902 2320 5908 2332
rect 5960 2320 5966 2372
rect 4571 2264 4844 2292
rect 4985 2295 5043 2301
rect 4571 2261 4583 2264
rect 4525 2255 4583 2261
rect 4985 2261 4997 2295
rect 5031 2292 5043 2295
rect 6288 2292 6316 2400
rect 6822 2388 6828 2400
rect 6880 2428 6886 2440
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6880 2400 6929 2428
rect 6880 2388 6886 2400
rect 6917 2397 6929 2400
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7800 2400 7849 2428
rect 7800 2388 7806 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 8113 2431 8171 2437
rect 8113 2397 8125 2431
rect 8159 2428 8171 2431
rect 9858 2428 9864 2440
rect 8159 2400 9864 2428
rect 8159 2397 8171 2400
rect 8113 2391 8171 2397
rect 9858 2388 9864 2400
rect 9916 2388 9922 2440
rect 10229 2431 10287 2437
rect 10229 2397 10241 2431
rect 10275 2428 10287 2431
rect 10870 2428 10876 2440
rect 10275 2400 10876 2428
rect 10275 2397 10287 2400
rect 10229 2391 10287 2397
rect 10870 2388 10876 2400
rect 10928 2388 10934 2440
rect 11054 2428 11060 2440
rect 11015 2400 11060 2428
rect 11054 2388 11060 2400
rect 11112 2388 11118 2440
rect 12342 2428 12348 2440
rect 12303 2400 12348 2428
rect 12342 2388 12348 2400
rect 12400 2388 12406 2440
rect 12713 2431 12771 2437
rect 12713 2397 12725 2431
rect 12759 2397 12771 2431
rect 13354 2428 13360 2440
rect 13315 2400 13360 2428
rect 12713 2391 12771 2397
rect 6457 2363 6515 2369
rect 6457 2329 6469 2363
rect 6503 2360 6515 2363
rect 6641 2363 6699 2369
rect 6641 2360 6653 2363
rect 6503 2332 6653 2360
rect 6503 2329 6515 2332
rect 6457 2323 6515 2329
rect 6641 2329 6653 2332
rect 6687 2360 6699 2363
rect 8202 2360 8208 2372
rect 6687 2332 8208 2360
rect 6687 2329 6699 2332
rect 6641 2323 6699 2329
rect 8202 2320 8208 2332
rect 8260 2320 8266 2372
rect 8386 2320 8392 2372
rect 8444 2360 8450 2372
rect 9125 2363 9183 2369
rect 9125 2360 9137 2363
rect 8444 2332 9137 2360
rect 8444 2320 8450 2332
rect 9125 2329 9137 2332
rect 9171 2360 9183 2363
rect 9582 2360 9588 2372
rect 9171 2332 9588 2360
rect 9171 2329 9183 2332
rect 9125 2323 9183 2329
rect 9582 2320 9588 2332
rect 9640 2320 9646 2372
rect 12158 2320 12164 2372
rect 12216 2360 12222 2372
rect 12728 2360 12756 2391
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 13725 2431 13783 2437
rect 13725 2397 13737 2431
rect 13771 2397 13783 2431
rect 13725 2391 13783 2397
rect 12216 2332 12756 2360
rect 12216 2320 12222 2332
rect 12802 2320 12808 2372
rect 12860 2360 12866 2372
rect 13630 2360 13636 2372
rect 12860 2332 13636 2360
rect 12860 2320 12866 2332
rect 13630 2320 13636 2332
rect 13688 2360 13694 2372
rect 13740 2360 13768 2391
rect 13814 2388 13820 2440
rect 13872 2428 13878 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 13872 2400 14105 2428
rect 13872 2388 13878 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14458 2428 14464 2440
rect 14419 2400 14464 2428
rect 14093 2391 14151 2397
rect 14458 2388 14464 2400
rect 14516 2388 14522 2440
rect 14734 2388 14740 2440
rect 14792 2428 14798 2440
rect 14829 2431 14887 2437
rect 14829 2428 14841 2431
rect 14792 2400 14841 2428
rect 14792 2388 14798 2400
rect 14829 2397 14841 2400
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 15197 2431 15255 2437
rect 15197 2397 15209 2431
rect 15243 2428 15255 2431
rect 15286 2428 15292 2440
rect 15243 2400 15292 2428
rect 15243 2397 15255 2400
rect 15197 2391 15255 2397
rect 15286 2388 15292 2400
rect 15344 2388 15350 2440
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2397 15715 2431
rect 16114 2428 16120 2440
rect 16075 2400 16120 2428
rect 15657 2391 15715 2397
rect 13688 2332 13768 2360
rect 13688 2320 13694 2332
rect 14550 2320 14556 2372
rect 14608 2360 14614 2372
rect 15672 2360 15700 2391
rect 16114 2388 16120 2400
rect 16172 2388 16178 2440
rect 16669 2431 16727 2437
rect 16669 2397 16681 2431
rect 16715 2428 16727 2431
rect 16942 2428 16948 2440
rect 16715 2400 16948 2428
rect 16715 2397 16727 2400
rect 16669 2391 16727 2397
rect 16942 2388 16948 2400
rect 17000 2388 17006 2440
rect 17126 2388 17132 2440
rect 17184 2428 17190 2440
rect 17313 2431 17371 2437
rect 17313 2428 17325 2431
rect 17184 2400 17325 2428
rect 17184 2388 17190 2400
rect 17313 2397 17325 2400
rect 17359 2397 17371 2431
rect 17494 2428 17500 2440
rect 17455 2400 17500 2428
rect 17313 2391 17371 2397
rect 17494 2388 17500 2400
rect 17552 2388 17558 2440
rect 18233 2431 18291 2437
rect 18233 2397 18245 2431
rect 18279 2428 18291 2431
rect 18322 2428 18328 2440
rect 18279 2400 18328 2428
rect 18279 2397 18291 2400
rect 18233 2391 18291 2397
rect 18322 2388 18328 2400
rect 18380 2388 18386 2440
rect 18690 2428 18696 2440
rect 18651 2400 18696 2428
rect 18690 2388 18696 2400
rect 18748 2388 18754 2440
rect 19536 2437 19564 2468
rect 20254 2456 20260 2468
rect 20312 2456 20318 2508
rect 19521 2431 19579 2437
rect 19521 2397 19533 2431
rect 19567 2397 19579 2431
rect 19886 2428 19892 2440
rect 19847 2400 19892 2428
rect 19521 2391 19579 2397
rect 19886 2388 19892 2400
rect 19944 2388 19950 2440
rect 20364 2437 20392 2604
rect 19981 2431 20039 2437
rect 19981 2397 19993 2431
rect 20027 2397 20039 2431
rect 19981 2391 20039 2397
rect 20349 2431 20407 2437
rect 20349 2397 20361 2431
rect 20395 2397 20407 2431
rect 20714 2428 20720 2440
rect 20675 2400 20720 2428
rect 20349 2391 20407 2397
rect 14608 2332 15700 2360
rect 14608 2320 14614 2332
rect 16758 2320 16764 2372
rect 16816 2360 16822 2372
rect 19996 2360 20024 2391
rect 20714 2388 20720 2400
rect 20772 2388 20778 2440
rect 21174 2428 21180 2440
rect 21135 2400 21180 2428
rect 21174 2388 21180 2400
rect 21232 2388 21238 2440
rect 16816 2332 20024 2360
rect 16816 2320 16822 2332
rect 6730 2292 6736 2304
rect 5031 2264 6316 2292
rect 6691 2264 6736 2292
rect 5031 2261 5043 2264
rect 4985 2255 5043 2261
rect 6730 2252 6736 2264
rect 6788 2252 6794 2304
rect 9214 2292 9220 2304
rect 9175 2264 9220 2292
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 9490 2252 9496 2304
rect 9548 2292 9554 2304
rect 9769 2295 9827 2301
rect 9769 2292 9781 2295
rect 9548 2264 9781 2292
rect 9548 2252 9554 2264
rect 9769 2261 9781 2264
rect 9815 2261 9827 2295
rect 9769 2255 9827 2261
rect 13262 2252 13268 2304
rect 13320 2292 13326 2304
rect 13541 2295 13599 2301
rect 13541 2292 13553 2295
rect 13320 2264 13553 2292
rect 13320 2252 13326 2264
rect 13541 2261 13553 2264
rect 13587 2261 13599 2295
rect 13541 2255 13599 2261
rect 13909 2295 13967 2301
rect 13909 2261 13921 2295
rect 13955 2292 13967 2295
rect 14274 2292 14280 2304
rect 13955 2264 14280 2292
rect 13955 2261 13967 2264
rect 13909 2255 13967 2261
rect 14274 2252 14280 2264
rect 14332 2252 14338 2304
rect 14734 2252 14740 2304
rect 14792 2292 14798 2304
rect 15013 2295 15071 2301
rect 15013 2292 15025 2295
rect 14792 2264 15025 2292
rect 14792 2252 14798 2264
rect 15013 2261 15025 2264
rect 15059 2261 15071 2295
rect 15013 2255 15071 2261
rect 15102 2252 15108 2304
rect 15160 2292 15166 2304
rect 15381 2295 15439 2301
rect 15381 2292 15393 2295
rect 15160 2264 15393 2292
rect 15160 2252 15166 2264
rect 15381 2261 15393 2264
rect 15427 2261 15439 2295
rect 15381 2255 15439 2261
rect 15562 2252 15568 2304
rect 15620 2292 15626 2304
rect 15841 2295 15899 2301
rect 15841 2292 15853 2295
rect 15620 2264 15853 2292
rect 15620 2252 15626 2264
rect 15841 2261 15853 2264
rect 15887 2261 15899 2295
rect 15841 2255 15899 2261
rect 16022 2252 16028 2304
rect 16080 2292 16086 2304
rect 16301 2295 16359 2301
rect 16301 2292 16313 2295
rect 16080 2264 16313 2292
rect 16080 2252 16086 2264
rect 16301 2261 16313 2264
rect 16347 2261 16359 2295
rect 16301 2255 16359 2261
rect 16390 2252 16396 2304
rect 16448 2292 16454 2304
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 16448 2264 16865 2292
rect 16448 2252 16454 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 16942 2252 16948 2304
rect 17000 2292 17006 2304
rect 17129 2295 17187 2301
rect 17129 2292 17141 2295
rect 17000 2264 17141 2292
rect 17000 2252 17006 2264
rect 17129 2261 17141 2264
rect 17175 2261 17187 2295
rect 17129 2255 17187 2261
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 17681 2255 17739 2261
rect 17862 2252 17868 2304
rect 17920 2292 17926 2304
rect 18049 2295 18107 2301
rect 18049 2292 18061 2295
rect 17920 2264 18061 2292
rect 17920 2252 17926 2264
rect 18049 2261 18061 2264
rect 18095 2261 18107 2295
rect 18049 2255 18107 2261
rect 18322 2252 18328 2304
rect 18380 2292 18386 2304
rect 18509 2295 18567 2301
rect 18509 2292 18521 2295
rect 18380 2264 18521 2292
rect 18380 2252 18386 2264
rect 18509 2261 18521 2264
rect 18555 2261 18567 2295
rect 18509 2255 18567 2261
rect 18782 2252 18788 2304
rect 18840 2292 18846 2304
rect 19337 2295 19395 2301
rect 19337 2292 19349 2295
rect 18840 2264 19349 2292
rect 18840 2252 18846 2264
rect 19337 2261 19349 2264
rect 19383 2261 19395 2295
rect 19337 2255 19395 2261
rect 19702 2252 19708 2304
rect 19760 2292 19766 2304
rect 20165 2295 20223 2301
rect 20165 2292 20177 2295
rect 19760 2264 20177 2292
rect 19760 2252 19766 2264
rect 20165 2261 20177 2264
rect 20211 2261 20223 2295
rect 20165 2255 20223 2261
rect 20254 2252 20260 2304
rect 20312 2292 20318 2304
rect 20533 2295 20591 2301
rect 20533 2292 20545 2295
rect 20312 2264 20545 2292
rect 20312 2252 20318 2264
rect 20533 2261 20545 2264
rect 20579 2261 20591 2295
rect 20533 2255 20591 2261
rect 20622 2252 20628 2304
rect 20680 2292 20686 2304
rect 20901 2295 20959 2301
rect 20901 2292 20913 2295
rect 20680 2264 20913 2292
rect 20680 2252 20686 2264
rect 20901 2261 20913 2264
rect 20947 2261 20959 2295
rect 20901 2255 20959 2261
rect 21082 2252 21088 2304
rect 21140 2292 21146 2304
rect 21361 2295 21419 2301
rect 21361 2292 21373 2295
rect 21140 2264 21373 2292
rect 21140 2252 21146 2264
rect 21361 2261 21373 2264
rect 21407 2261 21419 2295
rect 21361 2255 21419 2261
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
rect 2498 2048 2504 2100
rect 2556 2088 2562 2100
rect 6638 2088 6644 2100
rect 2556 2060 6644 2088
rect 2556 2048 2562 2060
rect 6638 2048 6644 2060
rect 6696 2048 6702 2100
rect 11054 2048 11060 2100
rect 11112 2088 11118 2100
rect 14366 2088 14372 2100
rect 11112 2060 14372 2088
rect 11112 2048 11118 2060
rect 14366 2048 14372 2060
rect 14424 2048 14430 2100
rect 9214 1980 9220 2032
rect 9272 2020 9278 2032
rect 17770 2020 17776 2032
rect 9272 1992 17776 2020
rect 9272 1980 9278 1992
rect 17770 1980 17776 1992
rect 17828 1980 17834 2032
rect 6730 1912 6736 1964
rect 6788 1952 6794 1964
rect 15010 1952 15016 1964
rect 6788 1924 15016 1952
rect 6788 1912 6794 1924
rect 15010 1912 15016 1924
rect 15068 1912 15074 1964
<< via1 >>
rect 10508 20952 10560 21004
rect 15200 20952 15252 21004
rect 11796 20884 11848 20936
rect 14096 20884 14148 20936
rect 11888 20816 11940 20868
rect 12808 20816 12860 20868
rect 12164 20748 12216 20800
rect 13912 20748 13964 20800
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 1860 20587 1912 20596
rect 1860 20553 1869 20587
rect 1869 20553 1903 20587
rect 1903 20553 1912 20587
rect 1860 20544 1912 20553
rect 2228 20587 2280 20596
rect 2228 20553 2237 20587
rect 2237 20553 2271 20587
rect 2271 20553 2280 20587
rect 2228 20544 2280 20553
rect 2964 20587 3016 20596
rect 2964 20553 2973 20587
rect 2973 20553 3007 20587
rect 3007 20553 3016 20587
rect 2964 20544 3016 20553
rect 4160 20544 4212 20596
rect 6828 20544 6880 20596
rect 9128 20544 9180 20596
rect 9496 20544 9548 20596
rect 1768 20408 1820 20460
rect 2044 20451 2096 20460
rect 2044 20417 2053 20451
rect 2053 20417 2087 20451
rect 2087 20417 2096 20451
rect 2044 20408 2096 20417
rect 2412 20451 2464 20460
rect 2412 20417 2421 20451
rect 2421 20417 2455 20451
rect 2455 20417 2464 20451
rect 2412 20408 2464 20417
rect 2504 20408 2556 20460
rect 3424 20451 3476 20460
rect 3424 20417 3433 20451
rect 3433 20417 3467 20451
rect 3467 20417 3476 20451
rect 3424 20408 3476 20417
rect 3884 20451 3936 20460
rect 3884 20417 3893 20451
rect 3893 20417 3927 20451
rect 3927 20417 3936 20451
rect 3884 20408 3936 20417
rect 4344 20408 4396 20460
rect 4804 20408 4856 20460
rect 5724 20408 5776 20460
rect 7104 20408 7156 20460
rect 7564 20408 7616 20460
rect 8300 20408 8352 20460
rect 8944 20451 8996 20460
rect 8944 20417 8953 20451
rect 8953 20417 8987 20451
rect 8987 20417 8996 20451
rect 8944 20408 8996 20417
rect 9404 20408 9456 20460
rect 4436 20272 4488 20324
rect 4988 20383 5040 20392
rect 4988 20349 4997 20383
rect 4997 20349 5031 20383
rect 5031 20349 5040 20383
rect 4988 20340 5040 20349
rect 5816 20272 5868 20324
rect 6644 20340 6696 20392
rect 7012 20383 7064 20392
rect 7012 20349 7021 20383
rect 7021 20349 7055 20383
rect 7055 20349 7064 20383
rect 7012 20340 7064 20349
rect 7748 20340 7800 20392
rect 10140 20383 10192 20392
rect 7380 20272 7432 20324
rect 10140 20349 10149 20383
rect 10149 20349 10183 20383
rect 10183 20349 10192 20383
rect 10140 20340 10192 20349
rect 9956 20272 10008 20324
rect 10324 20408 10376 20460
rect 12624 20519 12676 20528
rect 12624 20485 12642 20519
rect 12642 20485 12676 20519
rect 12624 20476 12676 20485
rect 12808 20476 12860 20528
rect 11704 20408 11756 20460
rect 12072 20408 12124 20460
rect 14096 20451 14148 20460
rect 14096 20417 14105 20451
rect 14105 20417 14139 20451
rect 14139 20417 14148 20451
rect 14096 20408 14148 20417
rect 12900 20383 12952 20392
rect 12900 20349 12909 20383
rect 12909 20349 12943 20383
rect 12943 20349 12952 20383
rect 12900 20340 12952 20349
rect 13452 20340 13504 20392
rect 11888 20272 11940 20324
rect 13912 20340 13964 20392
rect 14556 20544 14608 20596
rect 15384 20544 15436 20596
rect 15844 20544 15896 20596
rect 16304 20544 16356 20596
rect 17224 20544 17276 20596
rect 17960 20587 18012 20596
rect 17960 20553 17969 20587
rect 17969 20553 18003 20587
rect 18003 20553 18012 20587
rect 17960 20544 18012 20553
rect 18144 20544 18196 20596
rect 18604 20544 18656 20596
rect 14648 20476 14700 20528
rect 14556 20408 14608 20460
rect 15200 20451 15252 20460
rect 15200 20417 15209 20451
rect 15209 20417 15243 20451
rect 15243 20417 15252 20451
rect 15200 20408 15252 20417
rect 16028 20408 16080 20460
rect 17040 20451 17092 20460
rect 17040 20417 17049 20451
rect 17049 20417 17083 20451
rect 17083 20417 17092 20451
rect 17040 20408 17092 20417
rect 17132 20408 17184 20460
rect 17776 20451 17828 20460
rect 17776 20417 17785 20451
rect 17785 20417 17819 20451
rect 17819 20417 17828 20451
rect 17776 20408 17828 20417
rect 18236 20451 18288 20460
rect 18236 20417 18245 20451
rect 18245 20417 18279 20451
rect 18279 20417 18288 20451
rect 18236 20408 18288 20417
rect 18696 20451 18748 20460
rect 18696 20417 18705 20451
rect 18705 20417 18739 20451
rect 18739 20417 18748 20451
rect 18696 20408 18748 20417
rect 22744 20476 22796 20528
rect 19616 20408 19668 20460
rect 22284 20408 22336 20460
rect 18328 20340 18380 20392
rect 20812 20383 20864 20392
rect 20812 20349 20821 20383
rect 20821 20349 20855 20383
rect 20855 20349 20864 20383
rect 20812 20340 20864 20349
rect 14004 20272 14056 20324
rect 14924 20272 14976 20324
rect 16948 20272 17000 20324
rect 1492 20247 1544 20256
rect 1492 20213 1501 20247
rect 1501 20213 1535 20247
rect 1535 20213 1544 20247
rect 1492 20204 1544 20213
rect 3976 20204 4028 20256
rect 5908 20204 5960 20256
rect 6736 20204 6788 20256
rect 11060 20204 11112 20256
rect 13728 20204 13780 20256
rect 13820 20204 13872 20256
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 2412 20000 2464 20052
rect 3424 20000 3476 20052
rect 3884 20000 3936 20052
rect 4344 20000 4396 20052
rect 4804 20000 4856 20052
rect 5264 20043 5316 20052
rect 5264 20009 5273 20043
rect 5273 20009 5307 20043
rect 5307 20009 5316 20043
rect 5264 20000 5316 20009
rect 6000 20043 6052 20052
rect 6000 20009 6009 20043
rect 6009 20009 6043 20043
rect 6043 20009 6052 20043
rect 6000 20000 6052 20009
rect 7104 20000 7156 20052
rect 7472 20043 7524 20052
rect 7472 20009 7481 20043
rect 7481 20009 7515 20043
rect 7515 20009 7524 20043
rect 7472 20000 7524 20009
rect 9220 20000 9272 20052
rect 11796 20000 11848 20052
rect 11888 20000 11940 20052
rect 12900 20000 12952 20052
rect 13084 20000 13136 20052
rect 13728 20000 13780 20052
rect 2136 19932 2188 19984
rect 1676 19839 1728 19848
rect 1676 19805 1685 19839
rect 1685 19805 1719 19839
rect 1719 19805 1728 19839
rect 1676 19796 1728 19805
rect 2596 19864 2648 19916
rect 2136 19839 2188 19848
rect 2136 19805 2145 19839
rect 2145 19805 2179 19839
rect 2179 19805 2188 19839
rect 2136 19796 2188 19805
rect 9864 19864 9916 19916
rect 10692 19864 10744 19916
rect 11244 19864 11296 19916
rect 1584 19728 1636 19780
rect 5264 19796 5316 19848
rect 6552 19839 6604 19848
rect 6552 19805 6561 19839
rect 6561 19805 6595 19839
rect 6595 19805 6604 19839
rect 6552 19796 6604 19805
rect 7104 19796 7156 19848
rect 7656 19796 7708 19848
rect 8024 19839 8076 19848
rect 8024 19805 8033 19839
rect 8033 19805 8067 19839
rect 8067 19805 8076 19839
rect 8024 19796 8076 19805
rect 8116 19796 8168 19848
rect 8668 19796 8720 19848
rect 9404 19839 9456 19848
rect 9404 19805 9413 19839
rect 9413 19805 9447 19839
rect 9447 19805 9456 19839
rect 9404 19796 9456 19805
rect 10232 19839 10284 19848
rect 10232 19805 10241 19839
rect 10241 19805 10275 19839
rect 10275 19805 10284 19839
rect 10232 19796 10284 19805
rect 11152 19839 11204 19848
rect 11152 19805 11161 19839
rect 11161 19805 11195 19839
rect 11195 19805 11204 19839
rect 11152 19796 11204 19805
rect 13452 19932 13504 19984
rect 17776 20000 17828 20052
rect 19616 20000 19668 20052
rect 12992 19864 13044 19916
rect 13544 19864 13596 19916
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 1860 19703 1912 19712
rect 1860 19669 1869 19703
rect 1869 19669 1903 19703
rect 1903 19669 1912 19703
rect 1860 19660 1912 19669
rect 2320 19703 2372 19712
rect 2320 19669 2329 19703
rect 2329 19669 2363 19703
rect 2363 19669 2372 19703
rect 2320 19660 2372 19669
rect 2688 19660 2740 19712
rect 5540 19703 5592 19712
rect 5540 19669 5549 19703
rect 5549 19669 5583 19703
rect 5583 19669 5592 19703
rect 5540 19660 5592 19669
rect 6644 19728 6696 19780
rect 8484 19728 8536 19780
rect 9220 19771 9272 19780
rect 9220 19737 9229 19771
rect 9229 19737 9263 19771
rect 9263 19737 9272 19771
rect 9220 19728 9272 19737
rect 10048 19728 10100 19780
rect 10600 19660 10652 19712
rect 11796 19660 11848 19712
rect 12624 19771 12676 19780
rect 12624 19737 12642 19771
rect 12642 19737 12676 19771
rect 12900 19839 12952 19848
rect 12900 19805 12909 19839
rect 12909 19805 12943 19839
rect 12943 19805 12952 19839
rect 13176 19839 13228 19848
rect 12900 19796 12952 19805
rect 13176 19805 13185 19839
rect 13185 19805 13219 19839
rect 13219 19805 13228 19839
rect 13176 19796 13228 19805
rect 14096 19839 14148 19848
rect 14096 19805 14105 19839
rect 14105 19805 14139 19839
rect 14139 19805 14148 19839
rect 14096 19796 14148 19805
rect 14464 19796 14516 19848
rect 19064 19932 19116 19984
rect 19524 19932 19576 19984
rect 21364 20000 21416 20052
rect 12624 19728 12676 19737
rect 14556 19728 14608 19780
rect 19524 19796 19576 19848
rect 20812 19728 20864 19780
rect 21272 19771 21324 19780
rect 21272 19737 21290 19771
rect 21290 19737 21324 19771
rect 21272 19728 21324 19737
rect 13452 19660 13504 19712
rect 13636 19660 13688 19712
rect 14096 19660 14148 19712
rect 14832 19660 14884 19712
rect 16304 19660 16356 19712
rect 19616 19660 19668 19712
rect 19984 19703 20036 19712
rect 19984 19669 19993 19703
rect 19993 19669 20027 19703
rect 20027 19669 20036 19703
rect 19984 19660 20036 19669
rect 20168 19703 20220 19712
rect 20168 19669 20177 19703
rect 20177 19669 20211 19703
rect 20211 19669 20220 19703
rect 20168 19660 20220 19669
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 2504 19456 2556 19508
rect 5724 19456 5776 19508
rect 8116 19456 8168 19508
rect 9588 19456 9640 19508
rect 9772 19499 9824 19508
rect 9772 19465 9781 19499
rect 9781 19465 9815 19499
rect 9815 19465 9824 19499
rect 9772 19456 9824 19465
rect 10048 19499 10100 19508
rect 10048 19465 10057 19499
rect 10057 19465 10091 19499
rect 10091 19465 10100 19499
rect 10048 19456 10100 19465
rect 11244 19499 11296 19508
rect 1860 19320 1912 19372
rect 204 19252 256 19304
rect 2688 19320 2740 19372
rect 6000 19320 6052 19372
rect 1124 19184 1176 19236
rect 1860 19184 1912 19236
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 5540 19184 5592 19236
rect 7196 19184 7248 19236
rect 8392 19363 8444 19372
rect 8392 19329 8401 19363
rect 8401 19329 8435 19363
rect 8435 19329 8444 19363
rect 8392 19320 8444 19329
rect 8944 19320 8996 19372
rect 9680 19388 9732 19440
rect 9588 19363 9640 19372
rect 9588 19329 9597 19363
rect 9597 19329 9631 19363
rect 9631 19329 9640 19363
rect 9588 19320 9640 19329
rect 10416 19388 10468 19440
rect 11244 19465 11253 19499
rect 11253 19465 11287 19499
rect 11287 19465 11296 19499
rect 11244 19456 11296 19465
rect 12440 19456 12492 19508
rect 20076 19456 20128 19508
rect 8300 19252 8352 19304
rect 10140 19320 10192 19372
rect 18236 19388 18288 19440
rect 10784 19252 10836 19304
rect 9312 19184 9364 19236
rect 9496 19227 9548 19236
rect 9496 19193 9505 19227
rect 9505 19193 9539 19227
rect 9539 19193 9548 19227
rect 9496 19184 9548 19193
rect 9864 19184 9916 19236
rect 11704 19363 11756 19372
rect 11704 19329 11713 19363
rect 11713 19329 11747 19363
rect 11747 19329 11756 19363
rect 11704 19320 11756 19329
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 12164 19363 12216 19372
rect 11888 19320 11940 19329
rect 12164 19329 12198 19363
rect 12198 19329 12216 19363
rect 12164 19320 12216 19329
rect 12440 19320 12492 19372
rect 13176 19320 13228 19372
rect 17040 19320 17092 19372
rect 13544 19295 13596 19304
rect 13544 19261 13553 19295
rect 13553 19261 13587 19295
rect 13587 19261 13596 19295
rect 13544 19252 13596 19261
rect 19984 19388 20036 19440
rect 20444 19388 20496 19440
rect 19892 19320 19944 19372
rect 20720 19320 20772 19372
rect 21180 19363 21232 19372
rect 21180 19329 21189 19363
rect 21189 19329 21223 19363
rect 21223 19329 21232 19363
rect 21180 19320 21232 19329
rect 11244 19184 11296 19236
rect 13268 19227 13320 19236
rect 7104 19116 7156 19168
rect 7380 19159 7432 19168
rect 7380 19125 7389 19159
rect 7389 19125 7423 19159
rect 7423 19125 7432 19159
rect 7380 19116 7432 19125
rect 8576 19159 8628 19168
rect 8576 19125 8585 19159
rect 8585 19125 8619 19159
rect 8619 19125 8628 19159
rect 8576 19116 8628 19125
rect 8944 19116 8996 19168
rect 9128 19116 9180 19168
rect 9772 19116 9824 19168
rect 10876 19159 10928 19168
rect 10876 19125 10885 19159
rect 10885 19125 10919 19159
rect 10919 19125 10928 19159
rect 10876 19116 10928 19125
rect 10968 19116 11020 19168
rect 13268 19193 13277 19227
rect 13277 19193 13311 19227
rect 13311 19193 13320 19227
rect 13268 19184 13320 19193
rect 13452 19227 13504 19236
rect 13452 19193 13461 19227
rect 13461 19193 13495 19227
rect 13495 19193 13504 19227
rect 13452 19184 13504 19193
rect 14648 19184 14700 19236
rect 16948 19116 17000 19168
rect 17684 19116 17736 19168
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 7564 18955 7616 18964
rect 7564 18921 7573 18955
rect 7573 18921 7607 18955
rect 7607 18921 7616 18955
rect 7564 18912 7616 18921
rect 8484 18912 8536 18964
rect 9128 18912 9180 18964
rect 9588 18912 9640 18964
rect 6920 18844 6972 18896
rect 9312 18844 9364 18896
rect 664 18776 716 18828
rect 1676 18751 1728 18760
rect 1676 18717 1685 18751
rect 1685 18717 1719 18751
rect 1719 18717 1728 18751
rect 1676 18708 1728 18717
rect 8576 18776 8628 18828
rect 8300 18751 8352 18760
rect 8300 18717 8309 18751
rect 8309 18717 8343 18751
rect 8343 18717 8352 18751
rect 8300 18708 8352 18717
rect 8760 18708 8812 18760
rect 10048 18844 10100 18896
rect 17132 18912 17184 18964
rect 20904 18912 20956 18964
rect 13452 18776 13504 18828
rect 9772 18751 9824 18760
rect 9772 18717 9781 18751
rect 9781 18717 9815 18751
rect 9815 18717 9824 18751
rect 9772 18708 9824 18717
rect 12900 18708 12952 18760
rect 14648 18708 14700 18760
rect 16948 18708 17000 18760
rect 17684 18708 17736 18760
rect 20352 18708 20404 18760
rect 20812 18708 20864 18760
rect 7656 18640 7708 18692
rect 8208 18640 8260 18692
rect 1492 18615 1544 18624
rect 1492 18581 1501 18615
rect 1501 18581 1535 18615
rect 1535 18581 1544 18615
rect 1492 18572 1544 18581
rect 5448 18572 5500 18624
rect 8484 18615 8536 18624
rect 8484 18581 8493 18615
rect 8493 18581 8527 18615
rect 8527 18581 8536 18615
rect 8484 18572 8536 18581
rect 9220 18572 9272 18624
rect 9496 18572 9548 18624
rect 9956 18615 10008 18624
rect 9956 18581 9965 18615
rect 9965 18581 9999 18615
rect 9999 18581 10008 18615
rect 9956 18572 10008 18581
rect 11060 18640 11112 18692
rect 11244 18572 11296 18624
rect 11888 18640 11940 18692
rect 11980 18572 12032 18624
rect 13084 18572 13136 18624
rect 16120 18615 16172 18624
rect 16120 18581 16129 18615
rect 16129 18581 16163 18615
rect 16163 18581 16172 18615
rect 16120 18572 16172 18581
rect 16396 18572 16448 18624
rect 18144 18640 18196 18692
rect 20444 18640 20496 18692
rect 20996 18751 21048 18760
rect 20996 18717 21005 18751
rect 21005 18717 21039 18751
rect 21039 18717 21048 18751
rect 20996 18708 21048 18717
rect 20076 18572 20128 18624
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 2044 18368 2096 18420
rect 5816 18368 5868 18420
rect 5908 18368 5960 18420
rect 9680 18368 9732 18420
rect 10324 18368 10376 18420
rect 5264 18300 5316 18352
rect 5724 18300 5776 18352
rect 6920 18300 6972 18352
rect 19524 18368 19576 18420
rect 19892 18368 19944 18420
rect 20812 18368 20864 18420
rect 10784 18343 10836 18352
rect 1952 18232 2004 18284
rect 2228 18232 2280 18284
rect 2872 18232 2924 18284
rect 7656 18232 7708 18284
rect 4988 18164 5040 18216
rect 7932 18207 7984 18216
rect 7932 18173 7941 18207
rect 7941 18173 7975 18207
rect 7975 18173 7984 18207
rect 7932 18164 7984 18173
rect 10784 18309 10793 18343
rect 10793 18309 10827 18343
rect 10827 18309 10836 18343
rect 10784 18300 10836 18309
rect 12532 18300 12584 18352
rect 14648 18343 14700 18352
rect 9220 18259 9272 18268
rect 9220 18225 9229 18259
rect 9229 18225 9263 18259
rect 9263 18225 9272 18259
rect 9220 18216 9272 18225
rect 10692 18232 10744 18284
rect 11704 18232 11756 18284
rect 12900 18275 12952 18284
rect 12900 18241 12920 18275
rect 12920 18241 12952 18275
rect 12900 18232 12952 18241
rect 13452 18232 13504 18284
rect 13820 18232 13872 18284
rect 14648 18309 14657 18343
rect 14657 18309 14691 18343
rect 14691 18309 14700 18343
rect 14648 18300 14700 18309
rect 16212 18275 16264 18284
rect 16212 18241 16230 18275
rect 16230 18241 16264 18275
rect 16212 18232 16264 18241
rect 16580 18232 16632 18284
rect 16948 18232 17000 18284
rect 17408 18232 17460 18284
rect 18144 18232 18196 18284
rect 19616 18300 19668 18352
rect 20444 18232 20496 18284
rect 21640 18368 21692 18420
rect 1860 18139 1912 18148
rect 1860 18105 1869 18139
rect 1869 18105 1903 18139
rect 1903 18105 1912 18139
rect 1860 18096 1912 18105
rect 8484 18096 8536 18148
rect 9128 18096 9180 18148
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 5356 18028 5408 18080
rect 7656 18028 7708 18080
rect 7840 18028 7892 18080
rect 8300 18028 8352 18080
rect 9496 18096 9548 18148
rect 9864 18096 9916 18148
rect 9404 18071 9456 18080
rect 9404 18037 9413 18071
rect 9413 18037 9447 18071
rect 9447 18037 9456 18071
rect 9404 18028 9456 18037
rect 10232 18028 10284 18080
rect 10416 18028 10468 18080
rect 10692 18028 10744 18080
rect 11520 18071 11572 18080
rect 11520 18037 11529 18071
rect 11529 18037 11563 18071
rect 11563 18037 11572 18071
rect 11520 18028 11572 18037
rect 12992 18028 13044 18080
rect 14648 18028 14700 18080
rect 16212 18028 16264 18080
rect 17868 18028 17920 18080
rect 19524 18096 19576 18148
rect 18144 18071 18196 18080
rect 18144 18037 18153 18071
rect 18153 18037 18187 18071
rect 18187 18037 18196 18071
rect 18144 18028 18196 18037
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 6920 17824 6972 17876
rect 9496 17824 9548 17876
rect 9680 17824 9732 17876
rect 10232 17824 10284 17876
rect 10416 17824 10468 17876
rect 12808 17824 12860 17876
rect 12900 17824 12952 17876
rect 5172 17731 5224 17740
rect 5172 17697 5181 17731
rect 5181 17697 5215 17731
rect 5215 17697 5224 17731
rect 5172 17688 5224 17697
rect 5356 17731 5408 17740
rect 5356 17697 5365 17731
rect 5365 17697 5399 17731
rect 5399 17697 5408 17731
rect 5356 17688 5408 17697
rect 6000 17688 6052 17740
rect 7748 17756 7800 17808
rect 9864 17756 9916 17808
rect 2504 17620 2556 17672
rect 4804 17620 4856 17672
rect 5448 17620 5500 17672
rect 7288 17688 7340 17740
rect 9680 17688 9732 17740
rect 13728 17824 13780 17876
rect 18328 17824 18380 17876
rect 13176 17688 13228 17740
rect 16396 17756 16448 17808
rect 17776 17756 17828 17808
rect 6552 17620 6604 17672
rect 9404 17620 9456 17672
rect 16212 17620 16264 17672
rect 16580 17620 16632 17672
rect 17868 17620 17920 17672
rect 21272 17663 21324 17672
rect 21272 17629 21281 17663
rect 21281 17629 21315 17663
rect 21315 17629 21324 17663
rect 21272 17620 21324 17629
rect 7472 17552 7524 17604
rect 12164 17552 12216 17604
rect 12992 17552 13044 17604
rect 16396 17552 16448 17604
rect 17040 17552 17092 17604
rect 20076 17595 20128 17604
rect 20076 17561 20110 17595
rect 20110 17561 20128 17595
rect 20076 17552 20128 17561
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 4896 17484 4948 17536
rect 5724 17484 5776 17536
rect 5908 17527 5960 17536
rect 5908 17493 5917 17527
rect 5917 17493 5951 17527
rect 5951 17493 5960 17527
rect 5908 17484 5960 17493
rect 7380 17484 7432 17536
rect 9128 17484 9180 17536
rect 9956 17484 10008 17536
rect 11704 17527 11756 17536
rect 11704 17493 11713 17527
rect 11713 17493 11747 17527
rect 11747 17493 11756 17527
rect 11704 17484 11756 17493
rect 16212 17484 16264 17536
rect 21180 17527 21232 17536
rect 21180 17493 21189 17527
rect 21189 17493 21223 17527
rect 21223 17493 21232 17527
rect 21180 17484 21232 17493
rect 21456 17527 21508 17536
rect 21456 17493 21465 17527
rect 21465 17493 21499 17527
rect 21499 17493 21508 17527
rect 21456 17484 21508 17493
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 1768 17280 1820 17332
rect 2596 17323 2648 17332
rect 2596 17289 2605 17323
rect 2605 17289 2639 17323
rect 2639 17289 2648 17323
rect 2596 17280 2648 17289
rect 2688 17280 2740 17332
rect 4436 17323 4488 17332
rect 4436 17289 4445 17323
rect 4445 17289 4479 17323
rect 4479 17289 4488 17323
rect 4436 17280 4488 17289
rect 4896 17323 4948 17332
rect 4896 17289 4905 17323
rect 4905 17289 4939 17323
rect 4939 17289 4948 17323
rect 4896 17280 4948 17289
rect 5816 17280 5868 17332
rect 7380 17323 7432 17332
rect 7380 17289 7389 17323
rect 7389 17289 7423 17323
rect 7423 17289 7432 17323
rect 7380 17280 7432 17289
rect 7932 17323 7984 17332
rect 7932 17289 7941 17323
rect 7941 17289 7975 17323
rect 7975 17289 7984 17323
rect 7932 17280 7984 17289
rect 8024 17280 8076 17332
rect 8484 17280 8536 17332
rect 9128 17323 9180 17332
rect 9128 17289 9137 17323
rect 9137 17289 9171 17323
rect 9171 17289 9180 17323
rect 9128 17280 9180 17289
rect 10048 17323 10100 17332
rect 10048 17289 10057 17323
rect 10057 17289 10091 17323
rect 10091 17289 10100 17323
rect 10048 17280 10100 17289
rect 1676 17187 1728 17196
rect 1676 17153 1685 17187
rect 1685 17153 1719 17187
rect 1719 17153 1728 17187
rect 1676 17144 1728 17153
rect 4160 17212 4212 17264
rect 4620 17212 4672 17264
rect 5724 17212 5776 17264
rect 7840 17255 7892 17264
rect 7840 17221 7849 17255
rect 7849 17221 7883 17255
rect 7883 17221 7892 17255
rect 7840 17212 7892 17221
rect 8116 17212 8168 17264
rect 12808 17280 12860 17332
rect 13176 17280 13228 17332
rect 3056 17187 3108 17196
rect 3056 17153 3065 17187
rect 3065 17153 3099 17187
rect 3099 17153 3108 17187
rect 3056 17144 3108 17153
rect 2964 17076 3016 17128
rect 3516 17144 3568 17196
rect 4712 17144 4764 17196
rect 8484 17187 8536 17196
rect 8484 17153 8493 17187
rect 8493 17153 8527 17187
rect 8527 17153 8536 17187
rect 8484 17144 8536 17153
rect 9956 17187 10008 17196
rect 9956 17153 9965 17187
rect 9965 17153 9999 17187
rect 9999 17153 10008 17187
rect 9956 17144 10008 17153
rect 1492 16983 1544 16992
rect 1492 16949 1501 16983
rect 1501 16949 1535 16983
rect 1535 16949 1544 16983
rect 1492 16940 1544 16949
rect 1584 16940 1636 16992
rect 4436 17076 4488 17128
rect 5172 17076 5224 17128
rect 5724 17076 5776 17128
rect 6920 17076 6972 17128
rect 7748 17119 7800 17128
rect 7748 17085 7757 17119
rect 7757 17085 7791 17119
rect 7791 17085 7800 17119
rect 7748 17076 7800 17085
rect 9404 17119 9456 17128
rect 9404 17085 9413 17119
rect 9413 17085 9447 17119
rect 9447 17085 9456 17119
rect 9404 17076 9456 17085
rect 12440 17212 12492 17264
rect 13268 17255 13320 17264
rect 13268 17221 13302 17255
rect 13302 17221 13320 17255
rect 13268 17212 13320 17221
rect 9680 16940 9732 16992
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 13728 17212 13780 17264
rect 14648 17280 14700 17332
rect 16212 17255 16264 17264
rect 16212 17221 16230 17255
rect 16230 17221 16264 17255
rect 16212 17212 16264 17221
rect 14372 17144 14424 17196
rect 14648 17144 14700 17196
rect 16948 17144 17000 17196
rect 17868 17280 17920 17332
rect 16488 17119 16540 17128
rect 11796 17008 11848 17060
rect 11612 16940 11664 16992
rect 16488 17085 16497 17119
rect 16497 17085 16531 17119
rect 16531 17085 16540 17119
rect 16488 17076 16540 17085
rect 13176 16940 13228 16992
rect 14372 16983 14424 16992
rect 14372 16949 14381 16983
rect 14381 16949 14415 16983
rect 14415 16949 14424 16983
rect 14372 16940 14424 16949
rect 17408 16940 17460 16992
rect 18144 17076 18196 17128
rect 20168 16940 20220 16992
rect 20352 16983 20404 16992
rect 20352 16949 20361 16983
rect 20361 16949 20395 16983
rect 20395 16949 20404 16983
rect 20352 16940 20404 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 2964 16779 3016 16788
rect 2964 16745 2973 16779
rect 2973 16745 3007 16779
rect 3007 16745 3016 16779
rect 2964 16736 3016 16745
rect 3424 16779 3476 16788
rect 3424 16745 3433 16779
rect 3433 16745 3467 16779
rect 3467 16745 3476 16779
rect 3424 16736 3476 16745
rect 4712 16779 4764 16788
rect 4712 16745 4721 16779
rect 4721 16745 4755 16779
rect 4755 16745 4764 16779
rect 4712 16736 4764 16745
rect 5356 16736 5408 16788
rect 8116 16736 8168 16788
rect 12348 16736 12400 16788
rect 12532 16736 12584 16788
rect 12992 16736 13044 16788
rect 4436 16668 4488 16720
rect 4988 16668 5040 16720
rect 4252 16643 4304 16652
rect 4252 16609 4261 16643
rect 4261 16609 4295 16643
rect 4295 16609 4304 16643
rect 6184 16643 6236 16652
rect 4252 16600 4304 16609
rect 6184 16609 6193 16643
rect 6193 16609 6227 16643
rect 6227 16609 6236 16643
rect 6184 16600 6236 16609
rect 7564 16643 7616 16652
rect 7564 16609 7573 16643
rect 7573 16609 7607 16643
rect 7607 16609 7616 16643
rect 7564 16600 7616 16609
rect 8116 16643 8168 16652
rect 8116 16609 8125 16643
rect 8125 16609 8159 16643
rect 8159 16609 8168 16643
rect 8116 16600 8168 16609
rect 8392 16600 8444 16652
rect 9680 16643 9732 16652
rect 1584 16532 1636 16584
rect 2044 16575 2096 16584
rect 2044 16541 2053 16575
rect 2053 16541 2087 16575
rect 2087 16541 2096 16575
rect 2044 16532 2096 16541
rect 4160 16532 4212 16584
rect 4344 16575 4396 16584
rect 4344 16541 4353 16575
rect 4353 16541 4387 16575
rect 4387 16541 4396 16575
rect 4344 16532 4396 16541
rect 4620 16532 4672 16584
rect 8208 16532 8260 16584
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 1860 16439 1912 16448
rect 1860 16405 1869 16439
rect 1869 16405 1903 16439
rect 1903 16405 1912 16439
rect 1860 16396 1912 16405
rect 3148 16396 3200 16448
rect 5908 16439 5960 16448
rect 5908 16405 5917 16439
rect 5917 16405 5951 16439
rect 5951 16405 5960 16439
rect 5908 16396 5960 16405
rect 6000 16439 6052 16448
rect 6000 16405 6009 16439
rect 6009 16405 6043 16439
rect 6043 16405 6052 16439
rect 6000 16396 6052 16405
rect 8116 16396 8168 16448
rect 8668 16439 8720 16448
rect 8668 16405 8677 16439
rect 8677 16405 8711 16439
rect 8711 16405 8720 16439
rect 8668 16396 8720 16405
rect 9680 16609 9689 16643
rect 9689 16609 9723 16643
rect 9723 16609 9732 16643
rect 9680 16600 9732 16609
rect 9220 16575 9272 16584
rect 9220 16541 9229 16575
rect 9229 16541 9263 16575
rect 9263 16541 9272 16575
rect 9220 16532 9272 16541
rect 9588 16532 9640 16584
rect 9128 16464 9180 16516
rect 10416 16600 10468 16652
rect 11612 16600 11664 16652
rect 15476 16736 15528 16788
rect 16212 16736 16264 16788
rect 17960 16736 18012 16788
rect 13636 16600 13688 16652
rect 19340 16600 19392 16652
rect 10232 16532 10284 16584
rect 11888 16532 11940 16584
rect 15752 16575 15804 16584
rect 10048 16464 10100 16516
rect 9312 16439 9364 16448
rect 9312 16405 9321 16439
rect 9321 16405 9355 16439
rect 9355 16405 9364 16439
rect 9312 16396 9364 16405
rect 9404 16396 9456 16448
rect 10324 16439 10376 16448
rect 10324 16405 10333 16439
rect 10333 16405 10367 16439
rect 10367 16405 10376 16439
rect 10324 16396 10376 16405
rect 12900 16464 12952 16516
rect 15476 16507 15528 16516
rect 15476 16473 15494 16507
rect 15494 16473 15528 16507
rect 15476 16464 15528 16473
rect 15752 16541 15761 16575
rect 15761 16541 15795 16575
rect 15795 16541 15804 16575
rect 15752 16532 15804 16541
rect 16488 16532 16540 16584
rect 21456 16575 21508 16584
rect 21456 16541 21465 16575
rect 21465 16541 21499 16575
rect 21499 16541 21508 16575
rect 21456 16532 21508 16541
rect 10784 16439 10836 16448
rect 10784 16405 10793 16439
rect 10793 16405 10827 16439
rect 10827 16405 10836 16439
rect 10784 16396 10836 16405
rect 11060 16396 11112 16448
rect 12532 16396 12584 16448
rect 13636 16396 13688 16448
rect 14280 16396 14332 16448
rect 15200 16396 15252 16448
rect 15752 16396 15804 16448
rect 17960 16464 18012 16516
rect 18236 16464 18288 16516
rect 19064 16396 19116 16448
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 2872 16192 2924 16244
rect 3056 16192 3108 16244
rect 5908 16192 5960 16244
rect 8392 16235 8444 16244
rect 8392 16201 8401 16235
rect 8401 16201 8435 16235
rect 8435 16201 8444 16235
rect 8392 16192 8444 16201
rect 8760 16192 8812 16244
rect 9312 16192 9364 16244
rect 9772 16235 9824 16244
rect 9772 16201 9781 16235
rect 9781 16201 9815 16235
rect 9815 16201 9824 16235
rect 9772 16192 9824 16201
rect 2136 16056 2188 16108
rect 3148 16099 3200 16108
rect 3148 16065 3157 16099
rect 3157 16065 3191 16099
rect 3191 16065 3200 16099
rect 3148 16056 3200 16065
rect 5080 16056 5132 16108
rect 6368 16124 6420 16176
rect 6552 16124 6604 16176
rect 8116 16124 8168 16176
rect 9128 16124 9180 16176
rect 5172 15920 5224 15972
rect 5908 16056 5960 16108
rect 7840 16099 7892 16108
rect 7840 16065 7849 16099
rect 7849 16065 7883 16099
rect 7883 16065 7892 16099
rect 7840 16056 7892 16065
rect 8576 16056 8628 16108
rect 6000 15920 6052 15972
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 4896 15852 4948 15904
rect 5356 15852 5408 15904
rect 5908 15852 5960 15904
rect 6368 15895 6420 15904
rect 6368 15861 6377 15895
rect 6377 15861 6411 15895
rect 6411 15861 6420 15895
rect 6368 15852 6420 15861
rect 6920 15920 6972 15972
rect 7748 15988 7800 16040
rect 8576 15920 8628 15972
rect 7932 15852 7984 15904
rect 8392 15852 8444 15904
rect 9404 16056 9456 16108
rect 9864 16056 9916 16108
rect 10876 16192 10928 16244
rect 11060 16235 11112 16244
rect 11060 16201 11069 16235
rect 11069 16201 11103 16235
rect 11103 16201 11112 16235
rect 11060 16192 11112 16201
rect 11244 16192 11296 16244
rect 10784 16124 10836 16176
rect 13084 16124 13136 16176
rect 9956 16031 10008 16040
rect 9956 15997 9965 16031
rect 9965 15997 9999 16031
rect 9999 15997 10008 16031
rect 9956 15988 10008 15997
rect 9404 15895 9456 15904
rect 9404 15861 9413 15895
rect 9413 15861 9447 15895
rect 9447 15861 9456 15895
rect 9404 15852 9456 15861
rect 9772 15852 9824 15904
rect 12900 16056 12952 16108
rect 10508 16031 10560 16040
rect 10508 15997 10517 16031
rect 10517 15997 10551 16031
rect 10551 15997 10560 16031
rect 10508 15988 10560 15997
rect 11152 16031 11204 16040
rect 11152 15997 11161 16031
rect 11161 15997 11195 16031
rect 11195 15997 11204 16031
rect 11152 15988 11204 15997
rect 14924 16192 14976 16244
rect 15200 16124 15252 16176
rect 13636 16099 13688 16108
rect 13636 16065 13645 16099
rect 13645 16065 13679 16099
rect 13679 16065 13688 16099
rect 13636 16056 13688 16065
rect 15568 16056 15620 16108
rect 15200 16031 15252 16040
rect 12164 15963 12216 15972
rect 12164 15929 12173 15963
rect 12173 15929 12207 15963
rect 12207 15929 12216 15963
rect 12164 15920 12216 15929
rect 12440 15852 12492 15904
rect 15200 15997 15209 16031
rect 15209 15997 15243 16031
rect 15243 15997 15252 16031
rect 15200 15988 15252 15997
rect 20076 16124 20128 16176
rect 19064 16099 19116 16108
rect 19064 16065 19082 16099
rect 19082 16065 19116 16099
rect 19340 16099 19392 16108
rect 19064 16056 19116 16065
rect 19340 16065 19349 16099
rect 19349 16065 19383 16099
rect 19383 16065 19392 16099
rect 19340 16056 19392 16065
rect 21180 16099 21232 16108
rect 21180 16065 21198 16099
rect 21198 16065 21232 16099
rect 21180 16056 21232 16065
rect 21456 16099 21508 16108
rect 21456 16065 21465 16099
rect 21465 16065 21499 16099
rect 21499 16065 21508 16099
rect 21456 16056 21508 16065
rect 15568 15895 15620 15904
rect 15568 15861 15577 15895
rect 15577 15861 15611 15895
rect 15611 15861 15620 15895
rect 15568 15852 15620 15861
rect 16028 15852 16080 15904
rect 16396 15852 16448 15904
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 1676 15648 1728 15700
rect 1952 15648 2004 15700
rect 2504 15691 2556 15700
rect 2504 15657 2513 15691
rect 2513 15657 2547 15691
rect 2547 15657 2556 15691
rect 2504 15648 2556 15657
rect 5172 15691 5224 15700
rect 5172 15657 5181 15691
rect 5181 15657 5215 15691
rect 5215 15657 5224 15691
rect 5172 15648 5224 15657
rect 6000 15691 6052 15700
rect 6000 15657 6009 15691
rect 6009 15657 6043 15691
rect 6043 15657 6052 15691
rect 6000 15648 6052 15657
rect 6092 15691 6144 15700
rect 6092 15657 6101 15691
rect 6101 15657 6135 15691
rect 6135 15657 6144 15691
rect 6092 15648 6144 15657
rect 7840 15648 7892 15700
rect 1400 15444 1452 15496
rect 4068 15512 4120 15564
rect 4896 15580 4948 15632
rect 5448 15580 5500 15632
rect 5724 15580 5776 15632
rect 6368 15580 6420 15632
rect 5264 15512 5316 15564
rect 5356 15555 5408 15564
rect 5356 15521 5365 15555
rect 5365 15521 5399 15555
rect 5399 15521 5408 15555
rect 5356 15512 5408 15521
rect 5632 15512 5684 15564
rect 6736 15555 6788 15564
rect 6736 15521 6745 15555
rect 6745 15521 6779 15555
rect 6779 15521 6788 15555
rect 6736 15512 6788 15521
rect 7748 15555 7800 15564
rect 7748 15521 7757 15555
rect 7757 15521 7791 15555
rect 7791 15521 7800 15555
rect 7748 15512 7800 15521
rect 7932 15555 7984 15564
rect 7932 15521 7941 15555
rect 7941 15521 7975 15555
rect 7975 15521 7984 15555
rect 7932 15512 7984 15521
rect 8300 15580 8352 15632
rect 9772 15648 9824 15700
rect 10416 15648 10468 15700
rect 11336 15648 11388 15700
rect 11796 15648 11848 15700
rect 4436 15444 4488 15496
rect 4620 15444 4672 15496
rect 9312 15487 9364 15496
rect 4252 15376 4304 15428
rect 4528 15376 4580 15428
rect 9312 15453 9321 15487
rect 9321 15453 9355 15487
rect 9355 15453 9364 15487
rect 9312 15444 9364 15453
rect 9404 15444 9456 15496
rect 10600 15580 10652 15632
rect 16212 15648 16264 15700
rect 18236 15648 18288 15700
rect 11244 15512 11296 15564
rect 11152 15444 11204 15496
rect 13636 15512 13688 15564
rect 15384 15444 15436 15496
rect 17592 15444 17644 15496
rect 21456 15444 21508 15496
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 2872 15308 2924 15360
rect 3884 15308 3936 15360
rect 6552 15376 6604 15428
rect 7748 15376 7800 15428
rect 10968 15376 11020 15428
rect 13728 15376 13780 15428
rect 14556 15376 14608 15428
rect 14924 15376 14976 15428
rect 16396 15376 16448 15428
rect 21272 15419 21324 15428
rect 21272 15385 21290 15419
rect 21290 15385 21324 15419
rect 21272 15376 21324 15385
rect 6000 15308 6052 15360
rect 7012 15308 7064 15360
rect 8668 15308 8720 15360
rect 9680 15308 9732 15360
rect 10692 15351 10744 15360
rect 10692 15317 10701 15351
rect 10701 15317 10735 15351
rect 10735 15317 10744 15351
rect 10692 15308 10744 15317
rect 12808 15308 12860 15360
rect 13636 15308 13688 15360
rect 13820 15308 13872 15360
rect 19800 15351 19852 15360
rect 19800 15317 19809 15351
rect 19809 15317 19843 15351
rect 19843 15317 19852 15351
rect 19800 15308 19852 15317
rect 20628 15308 20680 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 2044 15104 2096 15156
rect 2228 15104 2280 15156
rect 3884 15104 3936 15156
rect 1768 14968 1820 15020
rect 2044 15011 2096 15020
rect 2044 14977 2053 15011
rect 2053 14977 2087 15011
rect 2087 14977 2096 15011
rect 2044 14968 2096 14977
rect 4344 15036 4396 15088
rect 5816 15104 5868 15156
rect 7472 15147 7524 15156
rect 7472 15113 7481 15147
rect 7481 15113 7515 15147
rect 7515 15113 7524 15147
rect 7472 15104 7524 15113
rect 7564 15104 7616 15156
rect 7932 15104 7984 15156
rect 4804 15036 4856 15088
rect 6828 15036 6880 15088
rect 2964 14900 3016 14952
rect 1860 14875 1912 14884
rect 1860 14841 1869 14875
rect 1869 14841 1903 14875
rect 1903 14841 1912 14875
rect 1860 14832 1912 14841
rect 2872 14832 2924 14884
rect 3424 14900 3476 14952
rect 4528 14900 4580 14952
rect 4896 14943 4948 14952
rect 4896 14909 4905 14943
rect 4905 14909 4939 14943
rect 4939 14909 4948 14943
rect 4896 14900 4948 14909
rect 5356 14900 5408 14952
rect 5724 14968 5776 15020
rect 8208 15011 8260 15020
rect 8208 14977 8217 15011
rect 8217 14977 8251 15011
rect 8251 14977 8260 15011
rect 8208 14968 8260 14977
rect 8576 15104 8628 15156
rect 9036 15147 9088 15156
rect 9036 15113 9045 15147
rect 9045 15113 9079 15147
rect 9079 15113 9088 15147
rect 9496 15147 9548 15156
rect 9036 15104 9088 15113
rect 9496 15113 9505 15147
rect 9505 15113 9539 15147
rect 9539 15113 9548 15147
rect 9496 15104 9548 15113
rect 10692 15104 10744 15156
rect 13452 15104 13504 15156
rect 13084 15036 13136 15088
rect 16948 15079 17000 15088
rect 16948 15045 16982 15079
rect 16982 15045 17000 15079
rect 16948 15036 17000 15045
rect 9772 14968 9824 15020
rect 10416 14968 10468 15020
rect 6736 14900 6788 14952
rect 6920 14943 6972 14952
rect 6920 14909 6929 14943
rect 6929 14909 6963 14943
rect 6963 14909 6972 14943
rect 6920 14900 6972 14909
rect 7288 14900 7340 14952
rect 8116 14900 8168 14952
rect 4620 14832 4672 14884
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 3976 14764 4028 14816
rect 6828 14832 6880 14884
rect 5816 14764 5868 14816
rect 6000 14807 6052 14816
rect 6000 14773 6009 14807
rect 6009 14773 6043 14807
rect 6043 14773 6052 14807
rect 6000 14764 6052 14773
rect 6736 14764 6788 14816
rect 7932 14832 7984 14884
rect 8024 14832 8076 14884
rect 9128 14900 9180 14952
rect 11704 14968 11756 15020
rect 11244 14943 11296 14952
rect 11244 14909 11253 14943
rect 11253 14909 11287 14943
rect 11287 14909 11296 14943
rect 11244 14900 11296 14909
rect 9680 14832 9732 14884
rect 12716 14968 12768 15020
rect 12900 14968 12952 15020
rect 15016 15011 15068 15020
rect 15016 14977 15034 15011
rect 15034 14977 15068 15011
rect 15016 14968 15068 14977
rect 15200 14968 15252 15020
rect 17684 14968 17736 15020
rect 19800 15036 19852 15088
rect 20720 14968 20772 15020
rect 19800 14900 19852 14952
rect 13636 14875 13688 14884
rect 13636 14841 13645 14875
rect 13645 14841 13679 14875
rect 13679 14841 13688 14875
rect 13636 14832 13688 14841
rect 7380 14764 7432 14816
rect 8116 14764 8168 14816
rect 9404 14807 9456 14816
rect 9404 14773 9413 14807
rect 9413 14773 9447 14807
rect 9447 14773 9456 14807
rect 9404 14764 9456 14773
rect 10416 14807 10468 14816
rect 10416 14773 10425 14807
rect 10425 14773 10459 14807
rect 10459 14773 10468 14807
rect 10416 14764 10468 14773
rect 12716 14764 12768 14816
rect 14280 14832 14332 14884
rect 14372 14764 14424 14816
rect 15752 14764 15804 14816
rect 18052 14807 18104 14816
rect 18052 14773 18061 14807
rect 18061 14773 18095 14807
rect 18095 14773 18104 14807
rect 18052 14764 18104 14773
rect 18328 14807 18380 14816
rect 18328 14773 18337 14807
rect 18337 14773 18371 14807
rect 18371 14773 18380 14807
rect 18328 14764 18380 14773
rect 21088 14764 21140 14816
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 4896 14560 4948 14612
rect 9128 14560 9180 14612
rect 9864 14603 9916 14612
rect 9864 14569 9873 14603
rect 9873 14569 9907 14603
rect 9907 14569 9916 14603
rect 9864 14560 9916 14569
rect 11244 14560 11296 14612
rect 4712 14492 4764 14544
rect 4620 14424 4672 14476
rect 5080 14467 5132 14476
rect 5080 14433 5089 14467
rect 5089 14433 5123 14467
rect 5123 14433 5132 14467
rect 5080 14424 5132 14433
rect 5816 14492 5868 14544
rect 1860 14356 1912 14408
rect 4160 14356 4212 14408
rect 5264 14399 5316 14408
rect 5264 14365 5273 14399
rect 5273 14365 5307 14399
rect 5307 14365 5316 14399
rect 7104 14424 7156 14476
rect 7472 14467 7524 14476
rect 7472 14433 7481 14467
rect 7481 14433 7515 14467
rect 7515 14433 7524 14467
rect 7472 14424 7524 14433
rect 7932 14424 7984 14476
rect 8300 14492 8352 14544
rect 8760 14492 8812 14544
rect 12164 14492 12216 14544
rect 8116 14467 8168 14476
rect 8116 14433 8125 14467
rect 8125 14433 8159 14467
rect 8159 14433 8168 14467
rect 9312 14467 9364 14476
rect 8116 14424 8168 14433
rect 9312 14433 9321 14467
rect 9321 14433 9355 14467
rect 9355 14433 9364 14467
rect 9312 14424 9364 14433
rect 9404 14424 9456 14476
rect 10508 14467 10560 14476
rect 10508 14433 10517 14467
rect 10517 14433 10551 14467
rect 10551 14433 10560 14467
rect 10508 14424 10560 14433
rect 11152 14424 11204 14476
rect 13636 14424 13688 14476
rect 13912 14424 13964 14476
rect 5264 14356 5316 14365
rect 6276 14356 6328 14408
rect 8852 14356 8904 14408
rect 10324 14399 10376 14408
rect 10324 14365 10333 14399
rect 10333 14365 10367 14399
rect 10367 14365 10376 14399
rect 10324 14356 10376 14365
rect 3424 14288 3476 14340
rect 7932 14331 7984 14340
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 4528 14220 4580 14272
rect 5632 14263 5684 14272
rect 5632 14229 5641 14263
rect 5641 14229 5675 14263
rect 5675 14229 5684 14263
rect 5632 14220 5684 14229
rect 6552 14220 6604 14272
rect 7564 14263 7616 14272
rect 7564 14229 7573 14263
rect 7573 14229 7607 14263
rect 7607 14229 7616 14263
rect 7564 14220 7616 14229
rect 7932 14297 7941 14331
rect 7941 14297 7975 14331
rect 7975 14297 7984 14331
rect 7932 14288 7984 14297
rect 9864 14220 9916 14272
rect 10968 14288 11020 14340
rect 13820 14356 13872 14408
rect 12164 14263 12216 14272
rect 12164 14229 12173 14263
rect 12173 14229 12207 14263
rect 12207 14229 12216 14263
rect 12164 14220 12216 14229
rect 13544 14220 13596 14272
rect 14464 14263 14516 14272
rect 14464 14229 14473 14263
rect 14473 14229 14507 14263
rect 14507 14229 14516 14263
rect 14464 14220 14516 14229
rect 15200 14560 15252 14612
rect 16212 14603 16264 14612
rect 16212 14569 16221 14603
rect 16221 14569 16255 14603
rect 16255 14569 16264 14603
rect 16212 14560 16264 14569
rect 18144 14560 18196 14612
rect 14832 14356 14884 14408
rect 15752 14356 15804 14408
rect 17592 14399 17644 14408
rect 17592 14365 17601 14399
rect 17601 14365 17635 14399
rect 17635 14365 17644 14399
rect 17592 14356 17644 14365
rect 21088 14399 21140 14408
rect 21088 14365 21097 14399
rect 21097 14365 21131 14399
rect 21131 14365 21140 14399
rect 21088 14356 21140 14365
rect 17500 14288 17552 14340
rect 20352 14288 20404 14340
rect 20904 14288 20956 14340
rect 19800 14220 19852 14272
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 5356 14059 5408 14068
rect 5356 14025 5365 14059
rect 5365 14025 5399 14059
rect 5399 14025 5408 14059
rect 5356 14016 5408 14025
rect 5724 14059 5776 14068
rect 5724 14025 5733 14059
rect 5733 14025 5767 14059
rect 5767 14025 5776 14059
rect 5724 14016 5776 14025
rect 6552 14016 6604 14068
rect 6736 14016 6788 14068
rect 7288 14059 7340 14068
rect 5264 13948 5316 14000
rect 1952 13880 2004 13932
rect 5448 13880 5500 13932
rect 5172 13812 5224 13864
rect 5540 13812 5592 13864
rect 7288 14025 7297 14059
rect 7297 14025 7331 14059
rect 7331 14025 7340 14059
rect 7288 14016 7340 14025
rect 7104 13948 7156 14000
rect 7564 13948 7616 14000
rect 7840 13948 7892 14000
rect 8484 14016 8536 14068
rect 10324 14016 10376 14068
rect 11244 14059 11296 14068
rect 11244 14025 11253 14059
rect 11253 14025 11287 14059
rect 11287 14025 11296 14059
rect 11244 14016 11296 14025
rect 8852 13948 8904 14000
rect 10140 13948 10192 14000
rect 10692 13948 10744 14000
rect 8392 13880 8444 13932
rect 9496 13880 9548 13932
rect 9680 13923 9732 13932
rect 9680 13889 9689 13923
rect 9689 13889 9723 13923
rect 9723 13889 9732 13923
rect 9680 13880 9732 13889
rect 9864 13880 9916 13932
rect 6920 13855 6972 13864
rect 6920 13821 6929 13855
rect 6929 13821 6963 13855
rect 6963 13821 6972 13855
rect 6920 13812 6972 13821
rect 7932 13812 7984 13864
rect 12164 13948 12216 14000
rect 14464 14016 14516 14068
rect 12532 13923 12584 13932
rect 12532 13889 12566 13923
rect 12566 13889 12584 13923
rect 12532 13880 12584 13889
rect 12900 13880 12952 13932
rect 10692 13812 10744 13864
rect 14924 13948 14976 14000
rect 17500 14016 17552 14068
rect 21272 14016 21324 14068
rect 21548 14059 21600 14068
rect 21548 14025 21557 14059
rect 21557 14025 21591 14059
rect 21591 14025 21600 14059
rect 21548 14016 21600 14025
rect 13820 13880 13872 13932
rect 17316 13880 17368 13932
rect 18328 13880 18380 13932
rect 20260 13880 20312 13932
rect 10784 13744 10836 13796
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 7656 13676 7708 13728
rect 10600 13676 10652 13728
rect 10876 13719 10928 13728
rect 10876 13685 10885 13719
rect 10885 13685 10919 13719
rect 10919 13685 10928 13719
rect 10876 13676 10928 13685
rect 17960 13812 18012 13864
rect 19524 13855 19576 13864
rect 13820 13787 13872 13796
rect 13820 13753 13829 13787
rect 13829 13753 13863 13787
rect 13863 13753 13872 13787
rect 13820 13744 13872 13753
rect 16028 13744 16080 13796
rect 19524 13821 19533 13855
rect 19533 13821 19567 13855
rect 19567 13821 19576 13855
rect 19524 13812 19576 13821
rect 12624 13676 12676 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 4436 13472 4488 13524
rect 5632 13472 5684 13524
rect 7932 13515 7984 13524
rect 5356 13404 5408 13456
rect 7104 13447 7156 13456
rect 6184 13379 6236 13388
rect 6184 13345 6193 13379
rect 6193 13345 6227 13379
rect 6227 13345 6236 13379
rect 6184 13336 6236 13345
rect 6460 13379 6512 13388
rect 6460 13345 6469 13379
rect 6469 13345 6503 13379
rect 6503 13345 6512 13379
rect 6460 13336 6512 13345
rect 7104 13413 7113 13447
rect 7113 13413 7147 13447
rect 7147 13413 7156 13447
rect 7104 13404 7156 13413
rect 7380 13379 7432 13388
rect 7380 13345 7389 13379
rect 7389 13345 7423 13379
rect 7423 13345 7432 13379
rect 7380 13336 7432 13345
rect 7932 13481 7941 13515
rect 7941 13481 7975 13515
rect 7975 13481 7984 13515
rect 7932 13472 7984 13481
rect 9220 13472 9272 13524
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 3148 13268 3200 13320
rect 8760 13404 8812 13456
rect 11888 13472 11940 13524
rect 8668 13379 8720 13388
rect 8668 13345 8677 13379
rect 8677 13345 8711 13379
rect 8711 13345 8720 13379
rect 8668 13336 8720 13345
rect 5724 13200 5776 13252
rect 6828 13200 6880 13252
rect 9404 13268 9456 13320
rect 10968 13336 11020 13388
rect 11980 13336 12032 13388
rect 12440 13336 12492 13388
rect 10876 13268 10928 13320
rect 11612 13268 11664 13320
rect 12624 13268 12676 13320
rect 12808 13311 12860 13320
rect 12808 13277 12842 13311
rect 12842 13277 12860 13311
rect 12808 13268 12860 13277
rect 17316 13472 17368 13524
rect 15200 13404 15252 13456
rect 17592 13472 17644 13524
rect 19524 13472 19576 13524
rect 18972 13447 19024 13456
rect 18972 13413 18981 13447
rect 18981 13413 19015 13447
rect 19015 13413 19024 13447
rect 20904 13472 20956 13524
rect 18972 13404 19024 13413
rect 17684 13268 17736 13320
rect 21180 13268 21232 13320
rect 9956 13200 10008 13252
rect 11796 13200 11848 13252
rect 18052 13200 18104 13252
rect 20168 13200 20220 13252
rect 7564 13175 7616 13184
rect 7564 13141 7573 13175
rect 7573 13141 7607 13175
rect 7607 13141 7616 13175
rect 8392 13175 8444 13184
rect 7564 13132 7616 13141
rect 8392 13141 8401 13175
rect 8401 13141 8435 13175
rect 8435 13141 8444 13175
rect 8392 13132 8444 13141
rect 9864 13175 9916 13184
rect 9864 13141 9873 13175
rect 9873 13141 9907 13175
rect 9907 13141 9916 13175
rect 9864 13132 9916 13141
rect 10416 13132 10468 13184
rect 10876 13132 10928 13184
rect 11244 13132 11296 13184
rect 13268 13132 13320 13184
rect 14096 13175 14148 13184
rect 14096 13141 14105 13175
rect 14105 13141 14139 13175
rect 14139 13141 14148 13175
rect 14096 13132 14148 13141
rect 15936 13175 15988 13184
rect 15936 13141 15945 13175
rect 15945 13141 15979 13175
rect 15979 13141 15988 13175
rect 15936 13132 15988 13141
rect 19892 13175 19944 13184
rect 19892 13141 19901 13175
rect 19901 13141 19935 13175
rect 19935 13141 19944 13175
rect 19892 13132 19944 13141
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 3148 12971 3200 12980
rect 3148 12937 3157 12971
rect 3157 12937 3191 12971
rect 3191 12937 3200 12971
rect 3148 12928 3200 12937
rect 4252 12971 4304 12980
rect 4252 12937 4261 12971
rect 4261 12937 4295 12971
rect 4295 12937 4304 12971
rect 4252 12928 4304 12937
rect 4160 12860 4212 12912
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 3884 12792 3936 12844
rect 6460 12928 6512 12980
rect 6736 12971 6788 12980
rect 6736 12937 6745 12971
rect 6745 12937 6779 12971
rect 6779 12937 6788 12971
rect 6736 12928 6788 12937
rect 4988 12835 5040 12844
rect 4528 12656 4580 12708
rect 4988 12801 4997 12835
rect 4997 12801 5031 12835
rect 5031 12801 5040 12835
rect 4988 12792 5040 12801
rect 5816 12835 5868 12844
rect 5816 12801 5825 12835
rect 5825 12801 5859 12835
rect 5859 12801 5868 12835
rect 5816 12792 5868 12801
rect 7656 12860 7708 12912
rect 8392 12928 8444 12980
rect 9588 12928 9640 12980
rect 10416 12971 10468 12980
rect 10416 12937 10425 12971
rect 10425 12937 10459 12971
rect 10459 12937 10468 12971
rect 10416 12928 10468 12937
rect 10876 12928 10928 12980
rect 13268 12928 13320 12980
rect 8392 12792 8444 12844
rect 8760 12792 8812 12844
rect 9312 12792 9364 12844
rect 9864 12792 9916 12844
rect 10600 12860 10652 12912
rect 13544 12860 13596 12912
rect 14188 12928 14240 12980
rect 17592 12928 17644 12980
rect 17868 12928 17920 12980
rect 5264 12767 5316 12776
rect 5264 12733 5273 12767
rect 5273 12733 5307 12767
rect 5307 12733 5316 12767
rect 5264 12724 5316 12733
rect 6276 12724 6328 12776
rect 6552 12724 6604 12776
rect 7288 12724 7340 12776
rect 7380 12724 7432 12776
rect 4160 12588 4212 12640
rect 4896 12588 4948 12640
rect 6920 12588 6972 12640
rect 8024 12588 8076 12640
rect 8576 12724 8628 12776
rect 9680 12656 9732 12708
rect 12164 12724 12216 12776
rect 14096 12835 14148 12844
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 14280 12792 14332 12844
rect 14832 12792 14884 12844
rect 15292 12835 15344 12844
rect 15936 12860 15988 12912
rect 16396 12860 16448 12912
rect 19892 12860 19944 12912
rect 20076 12860 20128 12912
rect 15292 12801 15310 12835
rect 15310 12801 15344 12835
rect 15292 12792 15344 12801
rect 16672 12835 16724 12844
rect 16672 12801 16681 12835
rect 16681 12801 16715 12835
rect 16715 12801 16724 12835
rect 16672 12792 16724 12801
rect 21088 12928 21140 12980
rect 21272 12928 21324 12980
rect 10968 12656 11020 12708
rect 11796 12656 11848 12708
rect 17684 12656 17736 12708
rect 8668 12588 8720 12640
rect 10232 12588 10284 12640
rect 10600 12588 10652 12640
rect 12624 12631 12676 12640
rect 12624 12597 12633 12631
rect 12633 12597 12667 12631
rect 12667 12597 12676 12631
rect 12624 12588 12676 12597
rect 12716 12631 12768 12640
rect 12716 12597 12725 12631
rect 12725 12597 12759 12631
rect 12759 12597 12768 12631
rect 12716 12588 12768 12597
rect 12992 12588 13044 12640
rect 13452 12588 13504 12640
rect 19524 12588 19576 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 1584 12384 1636 12436
rect 4068 12384 4120 12436
rect 4988 12384 5040 12436
rect 6828 12384 6880 12436
rect 7104 12384 7156 12436
rect 7840 12384 7892 12436
rect 8024 12384 8076 12436
rect 8208 12384 8260 12436
rect 6000 12316 6052 12368
rect 8576 12384 8628 12436
rect 8668 12384 8720 12436
rect 9956 12384 10008 12436
rect 10784 12384 10836 12436
rect 9312 12316 9364 12368
rect 5632 12248 5684 12300
rect 6276 12291 6328 12300
rect 6276 12257 6285 12291
rect 6285 12257 6319 12291
rect 6319 12257 6328 12291
rect 6276 12248 6328 12257
rect 6644 12248 6696 12300
rect 7380 12248 7432 12300
rect 8116 12291 8168 12300
rect 8116 12257 8125 12291
rect 8125 12257 8159 12291
rect 8159 12257 8168 12291
rect 8116 12248 8168 12257
rect 8208 12248 8260 12300
rect 9588 12291 9640 12300
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 3240 12180 3292 12232
rect 9312 12180 9364 12232
rect 9588 12257 9597 12291
rect 9597 12257 9631 12291
rect 9631 12257 9640 12291
rect 9588 12248 9640 12257
rect 11152 12316 11204 12368
rect 13728 12316 13780 12368
rect 17868 12384 17920 12436
rect 10968 12248 11020 12300
rect 16672 12291 16724 12300
rect 16672 12257 16681 12291
rect 16681 12257 16715 12291
rect 16715 12257 16724 12291
rect 16672 12248 16724 12257
rect 11060 12180 11112 12232
rect 2688 12044 2740 12096
rect 5080 12044 5132 12096
rect 6000 12087 6052 12096
rect 6000 12053 6009 12087
rect 6009 12053 6043 12087
rect 6043 12053 6052 12087
rect 6000 12044 6052 12053
rect 6552 12044 6604 12096
rect 7196 12112 7248 12164
rect 10416 12112 10468 12164
rect 10784 12112 10836 12164
rect 12348 12180 12400 12232
rect 12532 12223 12584 12232
rect 12532 12189 12541 12223
rect 12541 12189 12575 12223
rect 12575 12189 12584 12223
rect 12532 12180 12584 12189
rect 17040 12223 17092 12232
rect 17040 12189 17074 12223
rect 17074 12189 17092 12223
rect 18236 12248 18288 12300
rect 17040 12180 17092 12189
rect 11704 12112 11756 12164
rect 12072 12112 12124 12164
rect 12992 12112 13044 12164
rect 9128 12044 9180 12096
rect 10048 12044 10100 12096
rect 10600 12087 10652 12096
rect 10600 12053 10609 12087
rect 10609 12053 10643 12087
rect 10643 12053 10652 12087
rect 10600 12044 10652 12053
rect 10968 12044 11020 12096
rect 11152 12044 11204 12096
rect 13452 12044 13504 12096
rect 13544 12044 13596 12096
rect 15292 12112 15344 12164
rect 19524 12112 19576 12164
rect 14188 12087 14240 12096
rect 14188 12053 14197 12087
rect 14197 12053 14231 12087
rect 14231 12053 14240 12087
rect 14188 12044 14240 12053
rect 15016 12044 15068 12096
rect 20260 12112 20312 12164
rect 20996 12044 21048 12096
rect 21272 12180 21324 12232
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 2964 11840 3016 11892
rect 6552 11840 6604 11892
rect 7288 11883 7340 11892
rect 7288 11849 7297 11883
rect 7297 11849 7331 11883
rect 7331 11849 7340 11883
rect 7288 11840 7340 11849
rect 9680 11840 9732 11892
rect 10324 11840 10376 11892
rect 11244 11840 11296 11892
rect 12348 11840 12400 11892
rect 16304 11840 16356 11892
rect 5448 11772 5500 11824
rect 6920 11772 6972 11824
rect 7932 11772 7984 11824
rect 8116 11772 8168 11824
rect 10784 11772 10836 11824
rect 1400 11747 1452 11756
rect 1400 11713 1409 11747
rect 1409 11713 1443 11747
rect 1443 11713 1452 11747
rect 1400 11704 1452 11713
rect 1676 11747 1728 11756
rect 1676 11713 1685 11747
rect 1685 11713 1719 11747
rect 1719 11713 1728 11747
rect 1676 11704 1728 11713
rect 4160 11747 4212 11756
rect 4160 11713 4169 11747
rect 4169 11713 4203 11747
rect 4203 11713 4212 11747
rect 4160 11704 4212 11713
rect 6092 11704 6144 11756
rect 4988 11636 5040 11688
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 4528 11500 4580 11552
rect 6092 11500 6144 11552
rect 7288 11636 7340 11688
rect 8668 11704 8720 11756
rect 9220 11704 9272 11756
rect 9496 11704 9548 11756
rect 9680 11747 9732 11756
rect 9680 11713 9689 11747
rect 9689 11713 9723 11747
rect 9723 11713 9732 11747
rect 9680 11704 9732 11713
rect 11704 11704 11756 11756
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 13636 11747 13688 11756
rect 13636 11713 13654 11747
rect 13654 11713 13688 11747
rect 13636 11704 13688 11713
rect 16396 11704 16448 11756
rect 16488 11747 16540 11756
rect 16488 11713 16497 11747
rect 16497 11713 16531 11747
rect 16531 11713 16540 11747
rect 16488 11704 16540 11713
rect 7932 11679 7984 11688
rect 7932 11645 7941 11679
rect 7941 11645 7975 11679
rect 7975 11645 7984 11679
rect 7932 11636 7984 11645
rect 9956 11679 10008 11688
rect 9956 11645 9965 11679
rect 9965 11645 9999 11679
rect 9999 11645 10008 11679
rect 9956 11636 10008 11645
rect 10784 11679 10836 11688
rect 10784 11645 10793 11679
rect 10793 11645 10827 11679
rect 10827 11645 10836 11679
rect 10784 11636 10836 11645
rect 10968 11636 11020 11688
rect 11796 11636 11848 11688
rect 11980 11679 12032 11688
rect 11980 11645 11989 11679
rect 11989 11645 12023 11679
rect 12023 11645 12032 11679
rect 11980 11636 12032 11645
rect 9312 11611 9364 11620
rect 9312 11577 9321 11611
rect 9321 11577 9355 11611
rect 9355 11577 9364 11611
rect 9312 11568 9364 11577
rect 11060 11568 11112 11620
rect 12624 11568 12676 11620
rect 7104 11500 7156 11552
rect 7840 11500 7892 11552
rect 11152 11500 11204 11552
rect 11704 11500 11756 11552
rect 12532 11500 12584 11552
rect 13268 11500 13320 11552
rect 14188 11636 14240 11688
rect 20996 11772 21048 11824
rect 19892 11704 19944 11756
rect 16488 11568 16540 11620
rect 15016 11500 15068 11552
rect 15476 11500 15528 11552
rect 18236 11500 18288 11552
rect 18420 11500 18472 11552
rect 19616 11500 19668 11552
rect 20904 11500 20956 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 1768 11296 1820 11348
rect 2136 11339 2188 11348
rect 2136 11305 2145 11339
rect 2145 11305 2179 11339
rect 2179 11305 2188 11339
rect 2136 11296 2188 11305
rect 5264 11296 5316 11348
rect 5724 11296 5776 11348
rect 6000 11296 6052 11348
rect 7012 11339 7064 11348
rect 7012 11305 7021 11339
rect 7021 11305 7055 11339
rect 7055 11305 7064 11339
rect 7012 11296 7064 11305
rect 7288 11296 7340 11348
rect 4160 11228 4212 11280
rect 5448 11160 5500 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 3884 11092 3936 11144
rect 4988 11135 5040 11144
rect 4988 11101 4997 11135
rect 4997 11101 5031 11135
rect 5031 11101 5040 11135
rect 4988 11092 5040 11101
rect 5908 11160 5960 11212
rect 6920 11160 6972 11212
rect 7288 11160 7340 11212
rect 12808 11296 12860 11348
rect 10048 11271 10100 11280
rect 10048 11237 10057 11271
rect 10057 11237 10091 11271
rect 10091 11237 10100 11271
rect 10048 11228 10100 11237
rect 10324 11228 10376 11280
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 10416 11135 10468 11144
rect 10416 11101 10425 11135
rect 10425 11101 10459 11135
rect 10459 11101 10468 11135
rect 10416 11092 10468 11101
rect 3056 11024 3108 11076
rect 4252 11024 4304 11076
rect 4620 11024 4672 11076
rect 4896 11067 4948 11076
rect 4896 11033 4905 11067
rect 4905 11033 4939 11067
rect 4939 11033 4948 11067
rect 4896 11024 4948 11033
rect 5632 11024 5684 11076
rect 9312 11067 9364 11076
rect 9312 11033 9321 11067
rect 9321 11033 9355 11067
rect 9355 11033 9364 11067
rect 9312 11024 9364 11033
rect 10600 11203 10652 11212
rect 10600 11169 10609 11203
rect 10609 11169 10643 11203
rect 10643 11169 10652 11203
rect 10600 11160 10652 11169
rect 10876 11160 10928 11212
rect 11520 11228 11572 11280
rect 12624 11228 12676 11280
rect 15936 11296 15988 11348
rect 16120 11296 16172 11348
rect 16488 11296 16540 11348
rect 16948 11228 17000 11280
rect 11244 11092 11296 11144
rect 14280 11160 14332 11212
rect 15200 11203 15252 11212
rect 15200 11169 15209 11203
rect 15209 11169 15243 11203
rect 15243 11169 15252 11203
rect 15200 11160 15252 11169
rect 16396 11160 16448 11212
rect 12256 11092 12308 11144
rect 15292 11092 15344 11144
rect 20996 11203 21048 11212
rect 20996 11169 21005 11203
rect 21005 11169 21039 11203
rect 21039 11169 21048 11203
rect 20996 11160 21048 11169
rect 11428 11067 11480 11076
rect 6552 10999 6604 11008
rect 6552 10965 6561 10999
rect 6561 10965 6595 10999
rect 6595 10965 6604 10999
rect 6552 10956 6604 10965
rect 6644 10999 6696 11008
rect 6644 10965 6653 10999
rect 6653 10965 6687 10999
rect 6687 10965 6696 10999
rect 6644 10956 6696 10965
rect 8760 10956 8812 11008
rect 9404 10999 9456 11008
rect 9404 10965 9413 10999
rect 9413 10965 9447 10999
rect 9447 10965 9456 10999
rect 11428 11033 11437 11067
rect 11437 11033 11471 11067
rect 11471 11033 11480 11067
rect 11428 11024 11480 11033
rect 11612 11024 11664 11076
rect 12164 11024 12216 11076
rect 9404 10956 9456 10965
rect 12532 10956 12584 11008
rect 15568 11024 15620 11076
rect 17960 11024 18012 11076
rect 13268 10999 13320 11008
rect 13268 10965 13277 10999
rect 13277 10965 13311 10999
rect 13311 10965 13320 10999
rect 13268 10956 13320 10965
rect 13360 10956 13412 11008
rect 14648 10956 14700 11008
rect 19800 11024 19852 11076
rect 18420 10956 18472 11008
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 5172 10752 5224 10804
rect 5264 10752 5316 10804
rect 6644 10752 6696 10804
rect 7932 10752 7984 10804
rect 8760 10752 8812 10804
rect 9036 10795 9088 10804
rect 9036 10761 9045 10795
rect 9045 10761 9079 10795
rect 9079 10761 9088 10795
rect 9036 10752 9088 10761
rect 9404 10752 9456 10804
rect 9496 10795 9548 10804
rect 9496 10761 9505 10795
rect 9505 10761 9539 10795
rect 9539 10761 9548 10795
rect 9496 10752 9548 10761
rect 9680 10752 9732 10804
rect 11704 10752 11756 10804
rect 12440 10752 12492 10804
rect 12808 10752 12860 10804
rect 13360 10752 13412 10804
rect 3148 10684 3200 10736
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 4160 10616 4212 10668
rect 4436 10616 4488 10668
rect 8576 10727 8628 10736
rect 8576 10693 8585 10727
rect 8585 10693 8619 10727
rect 8619 10693 8628 10727
rect 8576 10684 8628 10693
rect 1584 10548 1636 10600
rect 2320 10548 2372 10600
rect 4068 10548 4120 10600
rect 4896 10548 4948 10600
rect 5724 10548 5776 10600
rect 7104 10616 7156 10668
rect 10600 10684 10652 10736
rect 10968 10684 11020 10736
rect 11244 10684 11296 10736
rect 6460 10591 6512 10600
rect 6460 10557 6469 10591
rect 6469 10557 6503 10591
rect 6503 10557 6512 10591
rect 6460 10548 6512 10557
rect 4804 10480 4856 10532
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 2964 10412 3016 10464
rect 6828 10548 6880 10600
rect 7932 10548 7984 10600
rect 9772 10616 9824 10668
rect 12808 10616 12860 10668
rect 15200 10684 15252 10736
rect 9496 10548 9548 10600
rect 9956 10591 10008 10600
rect 9956 10557 9965 10591
rect 9965 10557 9999 10591
rect 9999 10557 10008 10591
rect 9956 10548 10008 10557
rect 10876 10591 10928 10600
rect 10876 10557 10885 10591
rect 10885 10557 10919 10591
rect 10919 10557 10928 10591
rect 15108 10616 15160 10668
rect 15384 10659 15436 10668
rect 17500 10684 17552 10736
rect 15384 10625 15402 10659
rect 15402 10625 15436 10659
rect 15384 10616 15436 10625
rect 10876 10548 10928 10557
rect 13268 10548 13320 10600
rect 17868 10616 17920 10668
rect 18420 10591 18472 10600
rect 7288 10480 7340 10532
rect 11060 10480 11112 10532
rect 12992 10523 13044 10532
rect 12992 10489 13001 10523
rect 13001 10489 13035 10523
rect 13035 10489 13044 10523
rect 12992 10480 13044 10489
rect 9772 10412 9824 10464
rect 9864 10412 9916 10464
rect 13084 10412 13136 10464
rect 13820 10412 13872 10464
rect 18420 10557 18429 10591
rect 18429 10557 18463 10591
rect 18463 10557 18472 10591
rect 18420 10548 18472 10557
rect 21364 10591 21416 10600
rect 21364 10557 21373 10591
rect 21373 10557 21407 10591
rect 21407 10557 21416 10591
rect 21364 10548 21416 10557
rect 16488 10412 16540 10464
rect 17776 10412 17828 10464
rect 19708 10480 19760 10532
rect 19800 10455 19852 10464
rect 19800 10421 19809 10455
rect 19809 10421 19843 10455
rect 19843 10421 19852 10455
rect 19800 10412 19852 10421
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 2044 10208 2096 10260
rect 3148 10251 3200 10260
rect 3148 10217 3157 10251
rect 3157 10217 3191 10251
rect 3191 10217 3200 10251
rect 3148 10208 3200 10217
rect 3424 10208 3476 10260
rect 4344 10208 4396 10260
rect 5816 10208 5868 10260
rect 6828 10208 6880 10260
rect 7196 10251 7248 10260
rect 4896 10140 4948 10192
rect 3332 10072 3384 10124
rect 3792 10072 3844 10124
rect 4068 10115 4120 10124
rect 4068 10081 4077 10115
rect 4077 10081 4111 10115
rect 4111 10081 4120 10115
rect 4068 10072 4120 10081
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 3424 10004 3476 10056
rect 3976 10004 4028 10056
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 4988 10047 5040 10056
rect 4988 10013 4997 10047
rect 4997 10013 5031 10047
rect 5031 10013 5040 10047
rect 4988 10004 5040 10013
rect 5632 10072 5684 10124
rect 6092 10115 6144 10124
rect 6092 10081 6101 10115
rect 6101 10081 6135 10115
rect 6135 10081 6144 10115
rect 6092 10072 6144 10081
rect 6920 10140 6972 10192
rect 7196 10217 7205 10251
rect 7205 10217 7239 10251
rect 7239 10217 7248 10251
rect 7196 10208 7248 10217
rect 7564 10208 7616 10260
rect 7932 10208 7984 10260
rect 8668 10208 8720 10260
rect 14464 10208 14516 10260
rect 6644 10115 6696 10124
rect 6644 10081 6653 10115
rect 6653 10081 6687 10115
rect 6687 10081 6696 10115
rect 6644 10072 6696 10081
rect 6828 10072 6880 10124
rect 7012 10072 7064 10124
rect 13268 10115 13320 10124
rect 13268 10081 13277 10115
rect 13277 10081 13311 10115
rect 13311 10081 13320 10115
rect 13268 10072 13320 10081
rect 13452 10072 13504 10124
rect 8024 10004 8076 10056
rect 8576 10004 8628 10056
rect 9956 10004 10008 10056
rect 11244 10004 11296 10056
rect 17040 10047 17092 10056
rect 17040 10013 17049 10047
rect 17049 10013 17083 10047
rect 17083 10013 17092 10047
rect 17040 10004 17092 10013
rect 17776 10004 17828 10056
rect 2688 9911 2740 9920
rect 2688 9877 2697 9911
rect 2697 9877 2731 9911
rect 2731 9877 2740 9911
rect 2688 9868 2740 9877
rect 2780 9911 2832 9920
rect 2780 9877 2789 9911
rect 2789 9877 2823 9911
rect 2823 9877 2832 9911
rect 2780 9868 2832 9877
rect 4436 9868 4488 9920
rect 5908 9868 5960 9920
rect 6460 9868 6512 9920
rect 8484 9868 8536 9920
rect 9036 9868 9088 9920
rect 9404 9911 9456 9920
rect 9404 9877 9413 9911
rect 9413 9877 9447 9911
rect 9447 9877 9456 9911
rect 9404 9868 9456 9877
rect 9772 9911 9824 9920
rect 9772 9877 9781 9911
rect 9781 9877 9815 9911
rect 9815 9877 9824 9911
rect 9772 9868 9824 9877
rect 10048 9936 10100 9988
rect 14280 9936 14332 9988
rect 15936 9936 15988 9988
rect 16488 9936 16540 9988
rect 10508 9868 10560 9920
rect 10692 9868 10744 9920
rect 13728 9868 13780 9920
rect 15568 9911 15620 9920
rect 15568 9877 15577 9911
rect 15577 9877 15611 9911
rect 15611 9877 15620 9911
rect 15568 9868 15620 9877
rect 15660 9911 15712 9920
rect 15660 9877 15669 9911
rect 15669 9877 15703 9911
rect 15703 9877 15712 9911
rect 15660 9868 15712 9877
rect 16396 9868 16448 9920
rect 18052 9936 18104 9988
rect 18420 9936 18472 9988
rect 18512 9911 18564 9920
rect 18512 9877 18521 9911
rect 18521 9877 18555 9911
rect 18555 9877 18564 9911
rect 18512 9868 18564 9877
rect 19892 9868 19944 9920
rect 20536 9868 20588 9920
rect 20812 9911 20864 9920
rect 20812 9877 20821 9911
rect 20821 9877 20855 9911
rect 20855 9877 20864 9911
rect 20812 9868 20864 9877
rect 21364 9868 21416 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 1400 9707 1452 9716
rect 1400 9673 1409 9707
rect 1409 9673 1443 9707
rect 1443 9673 1452 9707
rect 1400 9664 1452 9673
rect 2780 9664 2832 9716
rect 10416 9664 10468 9716
rect 4436 9596 4488 9648
rect 5448 9639 5500 9648
rect 5448 9605 5457 9639
rect 5457 9605 5491 9639
rect 5491 9605 5500 9639
rect 5448 9596 5500 9605
rect 5540 9596 5592 9648
rect 1768 9571 1820 9580
rect 1768 9537 1777 9571
rect 1777 9537 1811 9571
rect 1811 9537 1820 9571
rect 1768 9528 1820 9537
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 2136 9528 2188 9580
rect 6092 9596 6144 9648
rect 6920 9596 6972 9648
rect 9772 9596 9824 9648
rect 12532 9664 12584 9716
rect 13176 9664 13228 9716
rect 10968 9596 11020 9648
rect 13820 9664 13872 9716
rect 20812 9664 20864 9716
rect 2228 9460 2280 9512
rect 5816 9528 5868 9580
rect 4804 9503 4856 9512
rect 4804 9469 4813 9503
rect 4813 9469 4847 9503
rect 4847 9469 4856 9503
rect 4804 9460 4856 9469
rect 1492 9392 1544 9444
rect 1860 9435 1912 9444
rect 1860 9401 1869 9435
rect 1869 9401 1903 9435
rect 1903 9401 1912 9435
rect 1860 9392 1912 9401
rect 1952 9392 2004 9444
rect 2412 9435 2464 9444
rect 2412 9401 2421 9435
rect 2421 9401 2455 9435
rect 2455 9401 2464 9435
rect 2412 9392 2464 9401
rect 2504 9392 2556 9444
rect 5172 9392 5224 9444
rect 5356 9460 5408 9512
rect 5448 9460 5500 9512
rect 9496 9528 9548 9580
rect 2780 9367 2832 9376
rect 2780 9333 2789 9367
rect 2789 9333 2823 9367
rect 2823 9333 2832 9367
rect 2780 9324 2832 9333
rect 4528 9324 4580 9376
rect 7012 9392 7064 9444
rect 7656 9392 7708 9444
rect 9772 9460 9824 9512
rect 12532 9528 12584 9580
rect 12624 9528 12676 9580
rect 13912 9596 13964 9648
rect 15660 9596 15712 9648
rect 5540 9324 5592 9376
rect 6736 9324 6788 9376
rect 8484 9324 8536 9376
rect 9312 9392 9364 9444
rect 10876 9460 10928 9512
rect 11888 9503 11940 9512
rect 11888 9469 11897 9503
rect 11897 9469 11931 9503
rect 11931 9469 11940 9503
rect 11888 9460 11940 9469
rect 12348 9460 12400 9512
rect 13820 9460 13872 9512
rect 15108 9528 15160 9580
rect 15200 9571 15252 9580
rect 15200 9537 15209 9571
rect 15209 9537 15243 9571
rect 15243 9537 15252 9571
rect 15200 9528 15252 9537
rect 17040 9528 17092 9580
rect 18236 9528 18288 9580
rect 20996 9528 21048 9580
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 16672 9435 16724 9444
rect 9036 9324 9088 9376
rect 9496 9324 9548 9376
rect 9772 9367 9824 9376
rect 9772 9333 9781 9367
rect 9781 9333 9815 9367
rect 9815 9333 9824 9367
rect 9772 9324 9824 9333
rect 10140 9324 10192 9376
rect 10508 9324 10560 9376
rect 10784 9324 10836 9376
rect 11704 9367 11756 9376
rect 11704 9333 11713 9367
rect 11713 9333 11747 9367
rect 11747 9333 11756 9367
rect 11704 9324 11756 9333
rect 12164 9324 12216 9376
rect 13452 9324 13504 9376
rect 16672 9401 16681 9435
rect 16681 9401 16715 9435
rect 16715 9401 16724 9435
rect 16672 9392 16724 9401
rect 13912 9324 13964 9376
rect 14280 9324 14332 9376
rect 17868 9324 17920 9376
rect 20720 9324 20772 9376
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 2136 9163 2188 9172
rect 2136 9129 2145 9163
rect 2145 9129 2179 9163
rect 2179 9129 2188 9163
rect 2136 9120 2188 9129
rect 2596 9120 2648 9172
rect 3056 9163 3108 9172
rect 3056 9129 3065 9163
rect 3065 9129 3099 9163
rect 3099 9129 3108 9163
rect 3056 9120 3108 9129
rect 3332 9163 3384 9172
rect 2964 9095 3016 9104
rect 2964 9061 2973 9095
rect 2973 9061 3007 9095
rect 3007 9061 3016 9095
rect 2964 9052 3016 9061
rect 3332 9129 3341 9163
rect 3341 9129 3375 9163
rect 3375 9129 3384 9163
rect 3332 9120 3384 9129
rect 3424 9120 3476 9172
rect 4344 8984 4396 9036
rect 5448 9120 5500 9172
rect 6552 9120 6604 9172
rect 7748 9120 7800 9172
rect 8024 9120 8076 9172
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 1676 8959 1728 8968
rect 1676 8925 1685 8959
rect 1685 8925 1719 8959
rect 1719 8925 1728 8959
rect 1676 8916 1728 8925
rect 2504 8916 2556 8968
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 2596 8916 2648 8925
rect 4068 8959 4120 8968
rect 2780 8848 2832 8900
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 8116 9052 8168 9104
rect 9588 9120 9640 9172
rect 9772 9120 9824 9172
rect 13636 9120 13688 9172
rect 10508 9052 10560 9104
rect 13452 9095 13504 9104
rect 13452 9061 13461 9095
rect 13461 9061 13495 9095
rect 13495 9061 13504 9095
rect 13452 9052 13504 9061
rect 13544 9052 13596 9104
rect 16120 9120 16172 9172
rect 5080 8984 5132 9036
rect 5724 8984 5776 9036
rect 5908 8984 5960 9036
rect 6828 9027 6880 9036
rect 6828 8993 6837 9027
rect 6837 8993 6871 9027
rect 6871 8993 6880 9027
rect 6828 8984 6880 8993
rect 8208 8984 8260 9036
rect 8484 9027 8536 9036
rect 8484 8993 8493 9027
rect 8493 8993 8527 9027
rect 8527 8993 8536 9027
rect 8484 8984 8536 8993
rect 8576 8984 8628 9036
rect 8760 8984 8812 9036
rect 10140 9027 10192 9036
rect 10140 8993 10149 9027
rect 10149 8993 10183 9027
rect 10183 8993 10192 9027
rect 10140 8984 10192 8993
rect 10324 9027 10376 9036
rect 10324 8993 10333 9027
rect 10333 8993 10367 9027
rect 10367 8993 10376 9027
rect 10324 8984 10376 8993
rect 10784 8984 10836 9036
rect 11704 8984 11756 9036
rect 4896 8959 4948 8968
rect 4896 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4948 8959
rect 4896 8916 4948 8925
rect 1952 8780 2004 8832
rect 2504 8823 2556 8832
rect 2504 8789 2513 8823
rect 2513 8789 2547 8823
rect 2547 8789 2556 8823
rect 2504 8780 2556 8789
rect 9956 8916 10008 8968
rect 10508 8916 10560 8968
rect 13820 8959 13872 8968
rect 13820 8925 13829 8959
rect 13829 8925 13863 8959
rect 13863 8925 13872 8959
rect 13820 8916 13872 8925
rect 15200 8916 15252 8968
rect 15752 8916 15804 8968
rect 18052 8916 18104 8968
rect 20628 8959 20680 8968
rect 20628 8925 20646 8959
rect 20646 8925 20680 8959
rect 20628 8916 20680 8925
rect 20812 8916 20864 8968
rect 5172 8848 5224 8900
rect 5356 8780 5408 8832
rect 5724 8823 5776 8832
rect 5724 8789 5733 8823
rect 5733 8789 5767 8823
rect 5767 8789 5776 8823
rect 7012 8848 7064 8900
rect 7288 8848 7340 8900
rect 5724 8780 5776 8789
rect 6552 8823 6604 8832
rect 6552 8789 6561 8823
rect 6561 8789 6595 8823
rect 6595 8789 6604 8823
rect 6552 8780 6604 8789
rect 6644 8823 6696 8832
rect 6644 8789 6653 8823
rect 6653 8789 6687 8823
rect 6687 8789 6696 8823
rect 6644 8780 6696 8789
rect 7748 8780 7800 8832
rect 7932 8848 7984 8900
rect 9772 8848 9824 8900
rect 12532 8848 12584 8900
rect 14464 8848 14516 8900
rect 16948 8848 17000 8900
rect 8208 8823 8260 8832
rect 8208 8789 8217 8823
rect 8217 8789 8251 8823
rect 8251 8789 8260 8823
rect 8208 8780 8260 8789
rect 8576 8780 8628 8832
rect 8760 8823 8812 8832
rect 8760 8789 8769 8823
rect 8769 8789 8803 8823
rect 8803 8789 8812 8823
rect 8760 8780 8812 8789
rect 10048 8823 10100 8832
rect 10048 8789 10057 8823
rect 10057 8789 10091 8823
rect 10091 8789 10100 8823
rect 10048 8780 10100 8789
rect 10508 8823 10560 8832
rect 10508 8789 10517 8823
rect 10517 8789 10551 8823
rect 10551 8789 10560 8823
rect 10508 8780 10560 8789
rect 13636 8823 13688 8832
rect 13636 8789 13645 8823
rect 13645 8789 13679 8823
rect 13679 8789 13688 8823
rect 13636 8780 13688 8789
rect 15200 8780 15252 8832
rect 16396 8780 16448 8832
rect 17500 8780 17552 8832
rect 19524 8823 19576 8832
rect 19524 8789 19533 8823
rect 19533 8789 19567 8823
rect 19567 8789 19576 8823
rect 19524 8780 19576 8789
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 1676 8619 1728 8628
rect 1676 8585 1685 8619
rect 1685 8585 1719 8619
rect 1719 8585 1728 8619
rect 1676 8576 1728 8585
rect 2044 8576 2096 8628
rect 2780 8576 2832 8628
rect 3976 8576 4028 8628
rect 4160 8576 4212 8628
rect 6000 8576 6052 8628
rect 6552 8576 6604 8628
rect 6920 8576 6972 8628
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 8576 8619 8628 8628
rect 8576 8585 8585 8619
rect 8585 8585 8619 8619
rect 8619 8585 8628 8619
rect 8576 8576 8628 8585
rect 9956 8619 10008 8628
rect 9956 8585 9965 8619
rect 9965 8585 9999 8619
rect 9999 8585 10008 8619
rect 9956 8576 10008 8585
rect 10048 8576 10100 8628
rect 10784 8576 10836 8628
rect 13544 8576 13596 8628
rect 13820 8619 13872 8628
rect 13820 8585 13829 8619
rect 13829 8585 13863 8619
rect 13863 8585 13872 8619
rect 13820 8576 13872 8585
rect 15108 8576 15160 8628
rect 15752 8619 15804 8628
rect 15752 8585 15761 8619
rect 15761 8585 15795 8619
rect 15795 8585 15804 8619
rect 15752 8576 15804 8585
rect 16120 8576 16172 8628
rect 17960 8576 18012 8628
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 2044 8440 2096 8492
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 3148 8440 3200 8492
rect 2136 8415 2188 8424
rect 2136 8381 2145 8415
rect 2145 8381 2179 8415
rect 2179 8381 2188 8415
rect 2136 8372 2188 8381
rect 2780 8304 2832 8356
rect 4344 8372 4396 8424
rect 6000 8440 6052 8492
rect 6092 8440 6144 8492
rect 6736 8440 6788 8492
rect 7472 8508 7524 8560
rect 9680 8508 9732 8560
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 5540 8372 5592 8381
rect 5724 8415 5776 8424
rect 5724 8381 5733 8415
rect 5733 8381 5767 8415
rect 5767 8381 5776 8415
rect 5724 8372 5776 8381
rect 5908 8372 5960 8424
rect 7380 8415 7432 8424
rect 7380 8381 7389 8415
rect 7389 8381 7423 8415
rect 7423 8381 7432 8415
rect 7380 8372 7432 8381
rect 7932 8415 7984 8424
rect 5172 8304 5224 8356
rect 7932 8381 7941 8415
rect 7941 8381 7975 8415
rect 7975 8381 7984 8415
rect 7932 8372 7984 8381
rect 8300 8372 8352 8424
rect 8208 8304 8260 8356
rect 8668 8372 8720 8424
rect 9128 8372 9180 8424
rect 9772 8440 9824 8492
rect 9864 8415 9916 8424
rect 9864 8381 9873 8415
rect 9873 8381 9907 8415
rect 9907 8381 9916 8415
rect 9864 8372 9916 8381
rect 10140 8508 10192 8560
rect 10048 8483 10100 8492
rect 10048 8449 10057 8483
rect 10057 8449 10091 8483
rect 10091 8449 10100 8483
rect 10048 8440 10100 8449
rect 10048 8304 10100 8356
rect 10416 8347 10468 8356
rect 10416 8313 10425 8347
rect 10425 8313 10459 8347
rect 10459 8313 10468 8347
rect 10416 8304 10468 8313
rect 10876 8304 10928 8356
rect 12164 8440 12216 8492
rect 14924 8508 14976 8560
rect 20628 8576 20680 8628
rect 13728 8372 13780 8424
rect 18052 8440 18104 8492
rect 20812 8508 20864 8560
rect 19432 8483 19484 8492
rect 19432 8449 19466 8483
rect 19466 8449 19484 8483
rect 19432 8440 19484 8449
rect 13636 8304 13688 8356
rect 5448 8236 5500 8288
rect 7656 8236 7708 8288
rect 8116 8236 8168 8288
rect 12716 8236 12768 8288
rect 18512 8304 18564 8356
rect 20444 8236 20496 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 1768 8032 1820 8084
rect 3884 8032 3936 8084
rect 5724 8032 5776 8084
rect 6920 8032 6972 8084
rect 7748 8032 7800 8084
rect 8024 8032 8076 8084
rect 9128 8032 9180 8084
rect 2412 7964 2464 8016
rect 4896 7964 4948 8016
rect 4988 7964 5040 8016
rect 6092 8007 6144 8016
rect 5448 7896 5500 7948
rect 6092 7973 6101 8007
rect 6101 7973 6135 8007
rect 6135 7973 6144 8007
rect 6092 7964 6144 7973
rect 5724 7939 5776 7948
rect 5724 7905 5733 7939
rect 5733 7905 5767 7939
rect 5767 7905 5776 7939
rect 5724 7896 5776 7905
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 2596 7828 2648 7880
rect 7196 7896 7248 7948
rect 8208 7896 8260 7948
rect 8484 7939 8536 7948
rect 8484 7905 8493 7939
rect 8493 7905 8527 7939
rect 8527 7905 8536 7939
rect 8484 7896 8536 7905
rect 10048 7896 10100 7948
rect 10324 7896 10376 7948
rect 10968 7896 11020 7948
rect 12808 8032 12860 8084
rect 14556 8032 14608 8084
rect 15108 8032 15160 8084
rect 17592 8032 17644 8084
rect 20168 8032 20220 8084
rect 20812 8032 20864 8084
rect 2688 7760 2740 7812
rect 5172 7760 5224 7812
rect 6552 7828 6604 7880
rect 6368 7760 6420 7812
rect 8668 7828 8720 7880
rect 9128 7828 9180 7880
rect 1952 7692 2004 7744
rect 4988 7692 5040 7744
rect 5908 7735 5960 7744
rect 5908 7701 5917 7735
rect 5917 7701 5951 7735
rect 5951 7701 5960 7735
rect 8024 7760 8076 7812
rect 9312 7760 9364 7812
rect 10508 7828 10560 7880
rect 11060 7828 11112 7880
rect 11336 7871 11388 7880
rect 11336 7837 11345 7871
rect 11345 7837 11379 7871
rect 11379 7837 11388 7871
rect 11336 7828 11388 7837
rect 14740 7964 14792 8016
rect 12348 7896 12400 7948
rect 12808 7939 12860 7948
rect 12808 7905 12817 7939
rect 12817 7905 12851 7939
rect 12851 7905 12860 7939
rect 19800 7964 19852 8016
rect 12808 7896 12860 7905
rect 5908 7692 5960 7701
rect 7288 7735 7340 7744
rect 7288 7701 7297 7735
rect 7297 7701 7331 7735
rect 7331 7701 7340 7735
rect 7288 7692 7340 7701
rect 8392 7692 8444 7744
rect 9772 7735 9824 7744
rect 9772 7701 9781 7735
rect 9781 7701 9815 7735
rect 9815 7701 9824 7735
rect 9772 7692 9824 7701
rect 10232 7735 10284 7744
rect 10232 7701 10241 7735
rect 10241 7701 10275 7735
rect 10275 7701 10284 7735
rect 11152 7760 11204 7812
rect 12532 7828 12584 7880
rect 12716 7828 12768 7880
rect 15292 7828 15344 7880
rect 13728 7760 13780 7812
rect 11796 7735 11848 7744
rect 10232 7692 10284 7701
rect 11796 7701 11805 7735
rect 11805 7701 11839 7735
rect 11839 7701 11848 7735
rect 11796 7692 11848 7701
rect 12072 7692 12124 7744
rect 12532 7692 12584 7744
rect 14280 7735 14332 7744
rect 14280 7701 14289 7735
rect 14289 7701 14323 7735
rect 14323 7701 14332 7735
rect 14280 7692 14332 7701
rect 15752 7692 15804 7744
rect 16028 7735 16080 7744
rect 16028 7701 16037 7735
rect 16037 7701 16071 7735
rect 16071 7701 16080 7735
rect 16028 7692 16080 7701
rect 17316 7692 17368 7744
rect 17408 7692 17460 7744
rect 21548 7828 21600 7880
rect 18512 7760 18564 7812
rect 20536 7803 20588 7812
rect 20536 7769 20554 7803
rect 20554 7769 20588 7803
rect 20536 7760 20588 7769
rect 17684 7735 17736 7744
rect 17684 7701 17693 7735
rect 17693 7701 17727 7735
rect 17727 7701 17736 7735
rect 17684 7692 17736 7701
rect 17868 7735 17920 7744
rect 17868 7701 17877 7735
rect 17877 7701 17911 7735
rect 17911 7701 17920 7735
rect 17868 7692 17920 7701
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 1492 7488 1544 7540
rect 2412 7488 2464 7540
rect 5632 7488 5684 7540
rect 6644 7488 6696 7540
rect 7288 7488 7340 7540
rect 7472 7531 7524 7540
rect 7472 7497 7481 7531
rect 7481 7497 7515 7531
rect 7515 7497 7524 7531
rect 7472 7488 7524 7497
rect 1584 7420 1636 7472
rect 5264 7420 5316 7472
rect 5448 7420 5500 7472
rect 8208 7420 8260 7472
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 4896 7352 4948 7404
rect 5632 7352 5684 7404
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 4988 7284 5040 7336
rect 5540 7327 5592 7336
rect 5540 7293 5549 7327
rect 5549 7293 5583 7327
rect 5583 7293 5592 7327
rect 5540 7284 5592 7293
rect 5908 7284 5960 7336
rect 6276 7284 6328 7336
rect 6920 7327 6972 7336
rect 6920 7293 6929 7327
rect 6929 7293 6963 7327
rect 6963 7293 6972 7327
rect 6920 7284 6972 7293
rect 7196 7352 7248 7404
rect 7840 7395 7892 7404
rect 7840 7361 7849 7395
rect 7849 7361 7883 7395
rect 7883 7361 7892 7395
rect 7840 7352 7892 7361
rect 8300 7352 8352 7404
rect 8116 7327 8168 7336
rect 8116 7293 8125 7327
rect 8125 7293 8159 7327
rect 8159 7293 8168 7327
rect 8116 7284 8168 7293
rect 8668 7395 8720 7404
rect 8668 7361 8677 7395
rect 8677 7361 8711 7395
rect 8711 7361 8720 7395
rect 8668 7352 8720 7361
rect 12072 7531 12124 7540
rect 12072 7497 12081 7531
rect 12081 7497 12115 7531
rect 12115 7497 12124 7531
rect 12072 7488 12124 7497
rect 13452 7531 13504 7540
rect 13452 7497 13461 7531
rect 13461 7497 13495 7531
rect 13495 7497 13504 7531
rect 13452 7488 13504 7497
rect 14280 7488 14332 7540
rect 14740 7531 14792 7540
rect 14740 7497 14749 7531
rect 14749 7497 14783 7531
rect 14783 7497 14792 7531
rect 14740 7488 14792 7497
rect 15108 7488 15160 7540
rect 17224 7488 17276 7540
rect 20812 7531 20864 7540
rect 10968 7463 11020 7472
rect 10968 7429 10977 7463
rect 10977 7429 11011 7463
rect 11011 7429 11020 7463
rect 10968 7420 11020 7429
rect 1584 7259 1636 7268
rect 1584 7225 1593 7259
rect 1593 7225 1627 7259
rect 1627 7225 1636 7259
rect 1584 7216 1636 7225
rect 5080 7216 5132 7268
rect 5172 7216 5224 7268
rect 5448 7148 5500 7200
rect 6000 7216 6052 7268
rect 9404 7284 9456 7336
rect 18236 7420 18288 7472
rect 20812 7497 20821 7531
rect 20821 7497 20855 7531
rect 20855 7497 20864 7531
rect 20812 7488 20864 7497
rect 11704 7284 11756 7336
rect 12716 7327 12768 7336
rect 12716 7293 12725 7327
rect 12725 7293 12759 7327
rect 12759 7293 12768 7327
rect 12716 7284 12768 7293
rect 9864 7148 9916 7200
rect 10600 7148 10652 7200
rect 11704 7148 11756 7200
rect 12164 7148 12216 7200
rect 12440 7148 12492 7200
rect 13820 7216 13872 7268
rect 14740 7352 14792 7404
rect 15200 7352 15252 7404
rect 20444 7395 20496 7404
rect 14924 7327 14976 7336
rect 14924 7293 14933 7327
rect 14933 7293 14967 7327
rect 14967 7293 14976 7327
rect 14924 7284 14976 7293
rect 20444 7361 20462 7395
rect 20462 7361 20496 7395
rect 20444 7352 20496 7361
rect 19524 7216 19576 7268
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 1400 6944 1452 6996
rect 5816 6944 5868 6996
rect 7196 6944 7248 6996
rect 8392 6987 8444 6996
rect 8392 6953 8401 6987
rect 8401 6953 8435 6987
rect 8435 6953 8444 6987
rect 8392 6944 8444 6953
rect 9312 6987 9364 6996
rect 9312 6953 9321 6987
rect 9321 6953 9355 6987
rect 9355 6953 9364 6987
rect 9312 6944 9364 6953
rect 4068 6851 4120 6860
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 4068 6817 4077 6851
rect 4077 6817 4111 6851
rect 4111 6817 4120 6851
rect 4068 6808 4120 6817
rect 4804 6808 4856 6860
rect 4896 6808 4948 6860
rect 4436 6740 4488 6792
rect 5724 6740 5776 6792
rect 6000 6740 6052 6792
rect 6644 6740 6696 6792
rect 6828 6783 6880 6792
rect 6828 6749 6837 6783
rect 6837 6749 6871 6783
rect 6871 6749 6880 6783
rect 6828 6740 6880 6749
rect 7104 6851 7156 6860
rect 7104 6817 7113 6851
rect 7113 6817 7147 6851
rect 7147 6817 7156 6851
rect 7104 6808 7156 6817
rect 7932 6808 7984 6860
rect 8208 6876 8260 6928
rect 9956 6944 10008 6996
rect 10232 6944 10284 6996
rect 10416 6944 10468 6996
rect 12072 6944 12124 6996
rect 13820 6944 13872 6996
rect 9680 6876 9732 6928
rect 9220 6851 9272 6860
rect 9220 6817 9229 6851
rect 9229 6817 9263 6851
rect 9263 6817 9272 6851
rect 9220 6808 9272 6817
rect 10324 6808 10376 6860
rect 10784 6851 10836 6860
rect 10784 6817 10793 6851
rect 10793 6817 10827 6851
rect 10827 6817 10836 6851
rect 10784 6808 10836 6817
rect 14004 6876 14056 6928
rect 17776 6876 17828 6928
rect 11704 6808 11756 6860
rect 12716 6808 12768 6860
rect 14740 6851 14792 6860
rect 14740 6817 14749 6851
rect 14749 6817 14783 6851
rect 14783 6817 14792 6851
rect 14740 6808 14792 6817
rect 9680 6783 9732 6792
rect 9680 6749 9689 6783
rect 9689 6749 9723 6783
rect 9723 6749 9732 6783
rect 9680 6740 9732 6749
rect 10968 6740 11020 6792
rect 17868 6740 17920 6792
rect 2504 6604 2556 6656
rect 3976 6604 4028 6656
rect 9956 6672 10008 6724
rect 10508 6715 10560 6724
rect 10508 6681 10517 6715
rect 10517 6681 10551 6715
rect 10551 6681 10560 6715
rect 10508 6672 10560 6681
rect 16028 6672 16080 6724
rect 4712 6647 4764 6656
rect 4712 6613 4721 6647
rect 4721 6613 4755 6647
rect 4755 6613 4764 6647
rect 4712 6604 4764 6613
rect 4988 6604 5040 6656
rect 5540 6604 5592 6656
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 6644 6604 6696 6656
rect 7932 6647 7984 6656
rect 7932 6613 7941 6647
rect 7941 6613 7975 6647
rect 7975 6613 7984 6647
rect 7932 6604 7984 6613
rect 8392 6604 8444 6656
rect 9036 6604 9088 6656
rect 9588 6604 9640 6656
rect 10600 6647 10652 6656
rect 10600 6613 10609 6647
rect 10609 6613 10643 6647
rect 10643 6613 10652 6647
rect 10600 6604 10652 6613
rect 11152 6604 11204 6656
rect 12440 6604 12492 6656
rect 12992 6604 13044 6656
rect 13268 6604 13320 6656
rect 14280 6604 14332 6656
rect 14832 6604 14884 6656
rect 15016 6604 15068 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 4620 6400 4672 6452
rect 2136 6332 2188 6384
rect 7380 6400 7432 6452
rect 8300 6400 8352 6452
rect 9036 6400 9088 6452
rect 9956 6443 10008 6452
rect 9956 6409 9965 6443
rect 9965 6409 9999 6443
rect 9999 6409 10008 6443
rect 9956 6400 10008 6409
rect 10600 6400 10652 6452
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 2044 6196 2096 6248
rect 4160 6196 4212 6248
rect 4712 6196 4764 6248
rect 7472 6264 7524 6316
rect 8300 6307 8352 6316
rect 7196 6196 7248 6248
rect 8024 6196 8076 6248
rect 8300 6273 8309 6307
rect 8309 6273 8343 6307
rect 8343 6273 8352 6307
rect 8300 6264 8352 6273
rect 9128 6307 9180 6316
rect 9128 6273 9137 6307
rect 9137 6273 9171 6307
rect 9171 6273 9180 6307
rect 9128 6264 9180 6273
rect 8484 6196 8536 6248
rect 9312 6239 9364 6248
rect 9312 6205 9321 6239
rect 9321 6205 9355 6239
rect 9355 6205 9364 6239
rect 9312 6196 9364 6205
rect 5264 6128 5316 6180
rect 11520 6264 11572 6316
rect 12624 6307 12676 6316
rect 10692 6239 10744 6248
rect 10692 6205 10701 6239
rect 10701 6205 10735 6239
rect 10735 6205 10744 6239
rect 10692 6196 10744 6205
rect 10876 6239 10928 6248
rect 10876 6205 10885 6239
rect 10885 6205 10919 6239
rect 10919 6205 10928 6239
rect 10876 6196 10928 6205
rect 11796 6196 11848 6248
rect 12624 6273 12633 6307
rect 12633 6273 12667 6307
rect 12667 6273 12676 6307
rect 12624 6264 12676 6273
rect 12716 6239 12768 6248
rect 11060 6128 11112 6180
rect 8116 6060 8168 6112
rect 10140 6060 10192 6112
rect 12440 6128 12492 6180
rect 12716 6205 12725 6239
rect 12725 6205 12759 6239
rect 12759 6205 12768 6239
rect 12716 6196 12768 6205
rect 15568 6400 15620 6452
rect 21180 6400 21232 6452
rect 13268 6264 13320 6316
rect 14004 6239 14056 6248
rect 14004 6205 14013 6239
rect 14013 6205 14047 6239
rect 14047 6205 14056 6239
rect 14004 6196 14056 6205
rect 21548 6307 21600 6316
rect 11612 6060 11664 6112
rect 11704 6103 11756 6112
rect 11704 6069 11713 6103
rect 11713 6069 11747 6103
rect 11747 6069 11756 6103
rect 11704 6060 11756 6069
rect 12716 6060 12768 6112
rect 13544 6128 13596 6180
rect 21548 6273 21557 6307
rect 21557 6273 21591 6307
rect 21591 6273 21600 6307
rect 21548 6264 21600 6273
rect 15660 6128 15712 6180
rect 15844 6060 15896 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 1400 5856 1452 5908
rect 7196 5899 7248 5908
rect 7196 5865 7205 5899
rect 7205 5865 7239 5899
rect 7239 5865 7248 5899
rect 7196 5856 7248 5865
rect 7288 5856 7340 5908
rect 8484 5856 8536 5908
rect 8576 5856 8628 5908
rect 1584 5831 1636 5840
rect 1584 5797 1593 5831
rect 1593 5797 1627 5831
rect 1627 5797 1636 5831
rect 1584 5788 1636 5797
rect 5080 5788 5132 5840
rect 10876 5856 10928 5908
rect 12900 5856 12952 5908
rect 13268 5899 13320 5908
rect 13268 5865 13277 5899
rect 13277 5865 13311 5899
rect 13311 5865 13320 5899
rect 13268 5856 13320 5865
rect 5356 5720 5408 5772
rect 5816 5763 5868 5772
rect 5816 5729 5825 5763
rect 5825 5729 5859 5763
rect 5859 5729 5868 5763
rect 5816 5720 5868 5729
rect 6552 5720 6604 5772
rect 7288 5720 7340 5772
rect 8116 5763 8168 5772
rect 8116 5729 8125 5763
rect 8125 5729 8159 5763
rect 8159 5729 8168 5763
rect 8116 5720 8168 5729
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 5172 5652 5224 5704
rect 6736 5652 6788 5704
rect 6920 5652 6972 5704
rect 16580 5788 16632 5840
rect 8852 5720 8904 5772
rect 10416 5720 10468 5772
rect 11520 5763 11572 5772
rect 11520 5729 11529 5763
rect 11529 5729 11563 5763
rect 11563 5729 11572 5763
rect 11520 5720 11572 5729
rect 11612 5720 11664 5772
rect 11796 5695 11848 5704
rect 11796 5661 11805 5695
rect 11805 5661 11839 5695
rect 11839 5661 11848 5695
rect 11796 5652 11848 5661
rect 13084 5720 13136 5772
rect 13268 5720 13320 5772
rect 13636 5720 13688 5772
rect 20720 5856 20772 5908
rect 18788 5788 18840 5840
rect 17592 5763 17644 5772
rect 17592 5729 17601 5763
rect 17601 5729 17635 5763
rect 17635 5729 17644 5763
rect 17592 5720 17644 5729
rect 20076 5763 20128 5772
rect 20076 5729 20085 5763
rect 20085 5729 20119 5763
rect 20119 5729 20128 5763
rect 20076 5720 20128 5729
rect 16488 5652 16540 5704
rect 4804 5584 4856 5636
rect 2228 5559 2280 5568
rect 2228 5525 2237 5559
rect 2237 5525 2271 5559
rect 2271 5525 2280 5559
rect 2228 5516 2280 5525
rect 4712 5516 4764 5568
rect 4988 5516 5040 5568
rect 5724 5516 5776 5568
rect 6644 5516 6696 5568
rect 7012 5516 7064 5568
rect 7380 5516 7432 5568
rect 7932 5559 7984 5568
rect 7932 5525 7941 5559
rect 7941 5525 7975 5559
rect 7975 5525 7984 5559
rect 7932 5516 7984 5525
rect 8760 5516 8812 5568
rect 9036 5516 9088 5568
rect 9772 5584 9824 5636
rect 10876 5584 10928 5636
rect 9588 5559 9640 5568
rect 9588 5525 9597 5559
rect 9597 5525 9631 5559
rect 9631 5525 9640 5559
rect 10692 5559 10744 5568
rect 9588 5516 9640 5525
rect 10692 5525 10701 5559
rect 10701 5525 10735 5559
rect 10735 5525 10744 5559
rect 10692 5516 10744 5525
rect 11060 5516 11112 5568
rect 11336 5516 11388 5568
rect 12808 5559 12860 5568
rect 12808 5525 12817 5559
rect 12817 5525 12851 5559
rect 12851 5525 12860 5559
rect 12808 5516 12860 5525
rect 12900 5559 12952 5568
rect 12900 5525 12909 5559
rect 12909 5525 12943 5559
rect 12943 5525 12952 5559
rect 13544 5559 13596 5568
rect 12900 5516 12952 5525
rect 13544 5525 13553 5559
rect 13553 5525 13587 5559
rect 13587 5525 13596 5559
rect 13544 5516 13596 5525
rect 16580 5516 16632 5568
rect 17776 5559 17828 5568
rect 17776 5525 17785 5559
rect 17785 5525 17819 5559
rect 17819 5525 17828 5559
rect 17776 5516 17828 5525
rect 20260 5559 20312 5568
rect 20260 5525 20269 5559
rect 20269 5525 20303 5559
rect 20303 5525 20312 5559
rect 20260 5516 20312 5525
rect 20812 5516 20864 5568
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 2228 5355 2280 5364
rect 2228 5321 2237 5355
rect 2237 5321 2271 5355
rect 2271 5321 2280 5355
rect 2228 5312 2280 5321
rect 5264 5312 5316 5364
rect 6644 5355 6696 5364
rect 6644 5321 6653 5355
rect 6653 5321 6687 5355
rect 6687 5321 6696 5355
rect 6644 5312 6696 5321
rect 2320 5244 2372 5296
rect 4620 5287 4672 5296
rect 4620 5253 4629 5287
rect 4629 5253 4663 5287
rect 4663 5253 4672 5287
rect 4620 5244 4672 5253
rect 5724 5244 5776 5296
rect 7932 5312 7984 5364
rect 9312 5355 9364 5364
rect 9312 5321 9321 5355
rect 9321 5321 9355 5355
rect 9355 5321 9364 5355
rect 9680 5355 9732 5364
rect 9312 5312 9364 5321
rect 9680 5321 9689 5355
rect 9689 5321 9723 5355
rect 9723 5321 9732 5355
rect 9680 5312 9732 5321
rect 10692 5312 10744 5364
rect 12808 5312 12860 5364
rect 13360 5312 13412 5364
rect 17776 5312 17828 5364
rect 1492 5219 1544 5228
rect 1492 5185 1501 5219
rect 1501 5185 1535 5219
rect 1535 5185 1544 5219
rect 1492 5176 1544 5185
rect 5356 5176 5408 5228
rect 5816 5176 5868 5228
rect 12072 5244 12124 5296
rect 2044 5151 2096 5160
rect 2044 5117 2053 5151
rect 2053 5117 2087 5151
rect 2087 5117 2096 5151
rect 2044 5108 2096 5117
rect 4988 5108 5040 5160
rect 4712 5040 4764 5092
rect 5080 5083 5132 5092
rect 5080 5049 5089 5083
rect 5089 5049 5123 5083
rect 5123 5049 5132 5083
rect 5080 5040 5132 5049
rect 2044 4972 2096 5024
rect 5724 5108 5776 5160
rect 6000 5151 6052 5160
rect 6000 5117 6009 5151
rect 6009 5117 6043 5151
rect 6043 5117 6052 5151
rect 6000 5108 6052 5117
rect 6552 5151 6604 5160
rect 6552 5117 6561 5151
rect 6561 5117 6595 5151
rect 6595 5117 6604 5151
rect 6552 5108 6604 5117
rect 6920 5040 6972 5092
rect 7840 5040 7892 5092
rect 7012 4972 7064 5024
rect 7196 4972 7248 5024
rect 8484 5151 8536 5160
rect 8484 5117 8493 5151
rect 8493 5117 8527 5151
rect 8527 5117 8536 5151
rect 9404 5176 9456 5228
rect 9496 5151 9548 5160
rect 8484 5108 8536 5117
rect 9496 5117 9505 5151
rect 9505 5117 9539 5151
rect 9539 5117 9548 5151
rect 9496 5108 9548 5117
rect 10876 5176 10928 5228
rect 12624 5176 12676 5228
rect 15844 5219 15896 5228
rect 10324 5151 10376 5160
rect 9128 5040 9180 5092
rect 10324 5117 10333 5151
rect 10333 5117 10367 5151
rect 10367 5117 10376 5151
rect 10324 5108 10376 5117
rect 10508 5151 10560 5160
rect 10508 5117 10517 5151
rect 10517 5117 10551 5151
rect 10551 5117 10560 5151
rect 10508 5108 10560 5117
rect 11980 5108 12032 5160
rect 12532 5151 12584 5160
rect 12532 5117 12541 5151
rect 12541 5117 12575 5151
rect 12575 5117 12584 5151
rect 12532 5108 12584 5117
rect 12716 5151 12768 5160
rect 12716 5117 12725 5151
rect 12725 5117 12759 5151
rect 12759 5117 12768 5151
rect 12716 5108 12768 5117
rect 9956 5040 10008 5092
rect 10968 5040 11020 5092
rect 11612 5040 11664 5092
rect 8484 4972 8536 5024
rect 8760 4972 8812 5024
rect 9496 4972 9548 5024
rect 11980 4972 12032 5024
rect 15844 5185 15853 5219
rect 15853 5185 15887 5219
rect 15887 5185 15896 5219
rect 15844 5176 15896 5185
rect 20812 5219 20864 5228
rect 20812 5185 20821 5219
rect 20821 5185 20855 5219
rect 20855 5185 20864 5219
rect 20812 5176 20864 5185
rect 15476 5151 15528 5160
rect 15476 5117 15485 5151
rect 15485 5117 15519 5151
rect 15519 5117 15528 5151
rect 15476 5108 15528 5117
rect 15568 5151 15620 5160
rect 15568 5117 15577 5151
rect 15577 5117 15611 5151
rect 15611 5117 15620 5151
rect 15568 5108 15620 5117
rect 12900 4972 12952 5024
rect 13452 5015 13504 5024
rect 13452 4981 13461 5015
rect 13461 4981 13495 5015
rect 13495 4981 13504 5015
rect 13452 4972 13504 4981
rect 14832 4972 14884 5024
rect 17040 4972 17092 5024
rect 20720 4972 20772 5024
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 4712 4768 4764 4820
rect 5540 4768 5592 4820
rect 5816 4811 5868 4820
rect 5816 4777 5825 4811
rect 5825 4777 5859 4811
rect 5859 4777 5868 4811
rect 5816 4768 5868 4777
rect 5908 4768 5960 4820
rect 7104 4811 7156 4820
rect 7104 4777 7113 4811
rect 7113 4777 7147 4811
rect 7147 4777 7156 4811
rect 7104 4768 7156 4777
rect 8576 4768 8628 4820
rect 4252 4700 4304 4752
rect 7012 4700 7064 4752
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 5356 4632 5408 4684
rect 2228 4607 2280 4616
rect 2228 4573 2237 4607
rect 2237 4573 2271 4607
rect 2271 4573 2280 4607
rect 2228 4564 2280 4573
rect 6000 4564 6052 4616
rect 7932 4700 7984 4752
rect 9312 4768 9364 4820
rect 9772 4811 9824 4820
rect 9772 4777 9781 4811
rect 9781 4777 9815 4811
rect 9815 4777 9824 4811
rect 9772 4768 9824 4777
rect 10876 4768 10928 4820
rect 11428 4811 11480 4820
rect 11428 4777 11437 4811
rect 11437 4777 11471 4811
rect 11471 4777 11480 4811
rect 11428 4768 11480 4777
rect 11888 4768 11940 4820
rect 11980 4768 12032 4820
rect 7656 4632 7708 4684
rect 10048 4700 10100 4752
rect 9956 4632 10008 4684
rect 10324 4700 10376 4752
rect 10784 4700 10836 4752
rect 10968 4743 11020 4752
rect 10968 4709 10977 4743
rect 10977 4709 11011 4743
rect 11011 4709 11020 4743
rect 10968 4700 11020 4709
rect 11336 4700 11388 4752
rect 11612 4743 11664 4752
rect 11612 4709 11621 4743
rect 11621 4709 11655 4743
rect 11655 4709 11664 4743
rect 11612 4700 11664 4709
rect 12624 4768 12676 4820
rect 15476 4811 15528 4820
rect 15476 4777 15485 4811
rect 15485 4777 15519 4811
rect 15519 4777 15528 4811
rect 15476 4768 15528 4777
rect 17500 4768 17552 4820
rect 20260 4768 20312 4820
rect 9772 4564 9824 4616
rect 14832 4675 14884 4684
rect 14832 4641 14841 4675
rect 14841 4641 14875 4675
rect 14875 4641 14884 4675
rect 14832 4632 14884 4641
rect 10876 4564 10928 4616
rect 14740 4607 14792 4616
rect 14740 4573 14749 4607
rect 14749 4573 14783 4607
rect 14783 4573 14792 4607
rect 14740 4564 14792 4573
rect 16948 4700 17000 4752
rect 16028 4675 16080 4684
rect 16028 4641 16037 4675
rect 16037 4641 16071 4675
rect 16071 4641 16080 4675
rect 16028 4632 16080 4641
rect 17592 4632 17644 4684
rect 15936 4564 15988 4616
rect 16304 4564 16356 4616
rect 18788 4607 18840 4616
rect 18788 4573 18797 4607
rect 18797 4573 18831 4607
rect 18831 4573 18840 4607
rect 18788 4564 18840 4573
rect 4528 4496 4580 4548
rect 5540 4496 5592 4548
rect 6920 4496 6972 4548
rect 11336 4496 11388 4548
rect 5908 4471 5960 4480
rect 5908 4437 5917 4471
rect 5917 4437 5951 4471
rect 5951 4437 5960 4471
rect 6736 4471 6788 4480
rect 5908 4428 5960 4437
rect 6736 4437 6745 4471
rect 6745 4437 6779 4471
rect 6779 4437 6788 4471
rect 6736 4428 6788 4437
rect 8024 4428 8076 4480
rect 8208 4428 8260 4480
rect 9312 4428 9364 4480
rect 9496 4428 9548 4480
rect 9680 4428 9732 4480
rect 11704 4471 11756 4480
rect 11704 4437 11713 4471
rect 11713 4437 11747 4471
rect 11747 4437 11756 4471
rect 11704 4428 11756 4437
rect 12624 4496 12676 4548
rect 17960 4496 18012 4548
rect 11980 4428 12032 4480
rect 12716 4428 12768 4480
rect 13728 4428 13780 4480
rect 14372 4471 14424 4480
rect 14372 4437 14381 4471
rect 14381 4437 14415 4471
rect 14415 4437 14424 4471
rect 14372 4428 14424 4437
rect 15844 4471 15896 4480
rect 15844 4437 15853 4471
rect 15853 4437 15887 4471
rect 15887 4437 15896 4471
rect 15844 4428 15896 4437
rect 15936 4471 15988 4480
rect 15936 4437 15945 4471
rect 15945 4437 15979 4471
rect 15979 4437 15988 4471
rect 17592 4471 17644 4480
rect 15936 4428 15988 4437
rect 17592 4437 17601 4471
rect 17601 4437 17635 4471
rect 17635 4437 17644 4471
rect 17592 4428 17644 4437
rect 17684 4471 17736 4480
rect 17684 4437 17693 4471
rect 17693 4437 17727 4471
rect 17727 4437 17736 4471
rect 17684 4428 17736 4437
rect 19892 4428 19944 4480
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 5908 4224 5960 4276
rect 8392 4224 8444 4276
rect 2596 4156 2648 4208
rect 5356 4156 5408 4208
rect 5724 4156 5776 4208
rect 6828 4156 6880 4208
rect 7196 4156 7248 4208
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 1952 4088 2004 4097
rect 2044 4088 2096 4140
rect 2688 4088 2740 4140
rect 4068 4088 4120 4140
rect 7656 4131 7708 4140
rect 2228 4063 2280 4072
rect 2228 4029 2237 4063
rect 2237 4029 2271 4063
rect 2271 4029 2280 4063
rect 2228 4020 2280 4029
rect 4252 3952 4304 4004
rect 5724 4063 5776 4072
rect 5724 4029 5733 4063
rect 5733 4029 5767 4063
rect 5767 4029 5776 4063
rect 7656 4097 7665 4131
rect 7665 4097 7699 4131
rect 7699 4097 7708 4131
rect 7656 4088 7708 4097
rect 8484 4199 8536 4208
rect 8484 4165 8493 4199
rect 8493 4165 8527 4199
rect 8527 4165 8536 4199
rect 9128 4224 9180 4276
rect 9404 4224 9456 4276
rect 9680 4224 9732 4276
rect 10048 4267 10100 4276
rect 10048 4233 10057 4267
rect 10057 4233 10091 4267
rect 10091 4233 10100 4267
rect 10048 4224 10100 4233
rect 10324 4224 10376 4276
rect 10508 4267 10560 4276
rect 10508 4233 10517 4267
rect 10517 4233 10551 4267
rect 10551 4233 10560 4267
rect 10508 4224 10560 4233
rect 9312 4199 9364 4208
rect 8484 4156 8536 4165
rect 9312 4165 9321 4199
rect 9321 4165 9355 4199
rect 9355 4165 9364 4199
rect 9312 4156 9364 4165
rect 9496 4156 9548 4208
rect 5724 4020 5776 4029
rect 7012 4063 7064 4072
rect 7012 4029 7021 4063
rect 7021 4029 7055 4063
rect 7055 4029 7064 4063
rect 7012 4020 7064 4029
rect 6552 3952 6604 4004
rect 1308 3884 1360 3936
rect 2780 3927 2832 3936
rect 2780 3893 2789 3927
rect 2789 3893 2823 3927
rect 2823 3893 2832 3927
rect 2780 3884 2832 3893
rect 2964 3927 3016 3936
rect 2964 3893 2973 3927
rect 2973 3893 3007 3927
rect 3007 3893 3016 3927
rect 6184 3927 6236 3936
rect 2964 3884 3016 3893
rect 6184 3893 6193 3927
rect 6193 3893 6227 3927
rect 6227 3893 6236 3927
rect 6184 3884 6236 3893
rect 6736 3884 6788 3936
rect 8024 4020 8076 4072
rect 7932 3884 7984 3936
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 9036 4020 9088 4072
rect 9956 4020 10008 4072
rect 9588 3952 9640 4004
rect 10232 4063 10284 4072
rect 10232 4029 10241 4063
rect 10241 4029 10275 4063
rect 10275 4029 10284 4063
rect 10232 4020 10284 4029
rect 10508 4088 10560 4140
rect 11612 4224 11664 4276
rect 11888 4267 11940 4276
rect 11888 4233 11897 4267
rect 11897 4233 11931 4267
rect 11931 4233 11940 4267
rect 11888 4224 11940 4233
rect 11980 4267 12032 4276
rect 11980 4233 11989 4267
rect 11989 4233 12023 4267
rect 12023 4233 12032 4267
rect 11980 4224 12032 4233
rect 11060 4156 11112 4208
rect 10876 4131 10928 4140
rect 10876 4097 10885 4131
rect 10885 4097 10919 4131
rect 10919 4097 10928 4131
rect 10876 4088 10928 4097
rect 11336 4020 11388 4072
rect 12992 4224 13044 4276
rect 15936 4224 15988 4276
rect 17592 4267 17644 4276
rect 17592 4233 17601 4267
rect 17601 4233 17635 4267
rect 17635 4233 17644 4267
rect 17592 4224 17644 4233
rect 18512 4267 18564 4276
rect 18512 4233 18521 4267
rect 18521 4233 18555 4267
rect 18555 4233 18564 4267
rect 18512 4224 18564 4233
rect 14372 4131 14424 4140
rect 14372 4097 14381 4131
rect 14381 4097 14415 4131
rect 14415 4097 14424 4131
rect 14372 4088 14424 4097
rect 12348 4020 12400 4072
rect 13636 4020 13688 4072
rect 17868 4156 17920 4208
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 17224 4088 17276 4140
rect 17592 4088 17644 4140
rect 10048 3884 10100 3936
rect 15844 3952 15896 4004
rect 18512 4020 18564 4072
rect 20996 3952 21048 4004
rect 12624 3927 12676 3936
rect 12624 3893 12633 3927
rect 12633 3893 12667 3927
rect 12667 3893 12676 3927
rect 12624 3884 12676 3893
rect 12900 3927 12952 3936
rect 12900 3893 12909 3927
rect 12909 3893 12943 3927
rect 12943 3893 12952 3927
rect 12900 3884 12952 3893
rect 14924 3884 14976 3936
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 388 3680 440 3732
rect 2320 3680 2372 3732
rect 5080 3680 5132 3732
rect 1676 3655 1728 3664
rect 1676 3621 1685 3655
rect 1685 3621 1719 3655
rect 1719 3621 1728 3655
rect 1676 3612 1728 3621
rect 2412 3612 2464 3664
rect 2596 3655 2648 3664
rect 2596 3621 2605 3655
rect 2605 3621 2639 3655
rect 2639 3621 2648 3655
rect 2596 3612 2648 3621
rect 3976 3612 4028 3664
rect 2780 3544 2832 3596
rect 4252 3587 4304 3596
rect 4252 3553 4261 3587
rect 4261 3553 4295 3587
rect 4295 3553 4304 3587
rect 4252 3544 4304 3553
rect 1492 3519 1544 3528
rect 1492 3485 1501 3519
rect 1501 3485 1535 3519
rect 1535 3485 1544 3519
rect 1492 3476 1544 3485
rect 1308 3408 1360 3460
rect 2320 3476 2372 3528
rect 1860 3451 1912 3460
rect 1860 3417 1869 3451
rect 1869 3417 1903 3451
rect 1903 3417 1912 3451
rect 7012 3680 7064 3732
rect 6552 3587 6604 3596
rect 6552 3553 6561 3587
rect 6561 3553 6595 3587
rect 6595 3553 6604 3587
rect 6552 3544 6604 3553
rect 7656 3544 7708 3596
rect 8944 3544 8996 3596
rect 9128 3587 9180 3596
rect 9128 3553 9137 3587
rect 9137 3553 9171 3587
rect 9171 3553 9180 3587
rect 9128 3544 9180 3553
rect 6736 3519 6788 3528
rect 6736 3485 6745 3519
rect 6745 3485 6779 3519
rect 6779 3485 6788 3519
rect 6736 3476 6788 3485
rect 1860 3408 1912 3417
rect 2320 3383 2372 3392
rect 2320 3349 2329 3383
rect 2329 3349 2363 3383
rect 2363 3349 2372 3383
rect 2320 3340 2372 3349
rect 2780 3340 2832 3392
rect 3148 3340 3200 3392
rect 3424 3383 3476 3392
rect 3424 3349 3433 3383
rect 3433 3349 3467 3383
rect 3467 3349 3476 3383
rect 3424 3340 3476 3349
rect 4252 3340 4304 3392
rect 7196 3408 7248 3460
rect 8668 3476 8720 3528
rect 9312 3519 9364 3528
rect 9312 3485 9321 3519
rect 9321 3485 9355 3519
rect 9355 3485 9364 3519
rect 9312 3476 9364 3485
rect 10876 3680 10928 3732
rect 13820 3680 13872 3732
rect 14096 3723 14148 3732
rect 14096 3689 14105 3723
rect 14105 3689 14139 3723
rect 14139 3689 14148 3723
rect 14096 3680 14148 3689
rect 17224 3723 17276 3732
rect 17224 3689 17233 3723
rect 17233 3689 17267 3723
rect 17267 3689 17276 3723
rect 17224 3680 17276 3689
rect 17868 3680 17920 3732
rect 19524 3680 19576 3732
rect 20352 3680 20404 3732
rect 21364 3723 21416 3732
rect 21364 3689 21373 3723
rect 21373 3689 21407 3723
rect 21407 3689 21416 3723
rect 21364 3680 21416 3689
rect 9588 3544 9640 3596
rect 10048 3587 10100 3596
rect 10048 3553 10057 3587
rect 10057 3553 10091 3587
rect 10091 3553 10100 3587
rect 10048 3544 10100 3553
rect 10692 3587 10744 3596
rect 10692 3553 10701 3587
rect 10701 3553 10735 3587
rect 10735 3553 10744 3587
rect 10692 3544 10744 3553
rect 11520 3587 11572 3596
rect 11520 3553 11529 3587
rect 11529 3553 11563 3587
rect 11563 3553 11572 3587
rect 11520 3544 11572 3553
rect 11612 3544 11664 3596
rect 13084 3544 13136 3596
rect 13268 3544 13320 3596
rect 14556 3612 14608 3664
rect 16212 3612 16264 3664
rect 17592 3612 17644 3664
rect 18880 3612 18932 3664
rect 8392 3408 8444 3460
rect 9496 3408 9548 3460
rect 11888 3408 11940 3460
rect 5356 3383 5408 3392
rect 5356 3349 5365 3383
rect 5365 3349 5399 3383
rect 5399 3349 5408 3383
rect 5356 3340 5408 3349
rect 5448 3340 5500 3392
rect 6644 3383 6696 3392
rect 6644 3349 6653 3383
rect 6653 3349 6687 3383
rect 6687 3349 6696 3383
rect 6644 3340 6696 3349
rect 7288 3383 7340 3392
rect 7288 3349 7297 3383
rect 7297 3349 7331 3383
rect 7331 3349 7340 3383
rect 7288 3340 7340 3349
rect 7564 3383 7616 3392
rect 7564 3349 7573 3383
rect 7573 3349 7607 3383
rect 7607 3349 7616 3383
rect 7564 3340 7616 3349
rect 7748 3383 7800 3392
rect 7748 3349 7757 3383
rect 7757 3349 7791 3383
rect 7791 3349 7800 3383
rect 7748 3340 7800 3349
rect 8300 3340 8352 3392
rect 9680 3340 9732 3392
rect 10232 3340 10284 3392
rect 22468 3476 22520 3528
rect 12992 3340 13044 3392
rect 13636 3408 13688 3460
rect 13728 3383 13780 3392
rect 13728 3349 13737 3383
rect 13737 3349 13771 3383
rect 13771 3349 13780 3383
rect 13728 3340 13780 3349
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 2136 3136 2188 3188
rect 2780 3136 2832 3188
rect 4068 3136 4120 3188
rect 4252 3179 4304 3188
rect 4252 3145 4261 3179
rect 4261 3145 4295 3179
rect 4295 3145 4304 3179
rect 4252 3136 4304 3145
rect 4344 3136 4396 3188
rect 4620 3179 4672 3188
rect 4620 3145 4629 3179
rect 4629 3145 4663 3179
rect 4663 3145 4672 3179
rect 4620 3136 4672 3145
rect 1768 3000 1820 3052
rect 2688 3043 2740 3052
rect 2688 3009 2697 3043
rect 2697 3009 2731 3043
rect 2731 3009 2740 3043
rect 2688 3000 2740 3009
rect 2780 3000 2832 3052
rect 2044 2932 2096 2984
rect 2136 2932 2188 2984
rect 2320 2932 2372 2984
rect 848 2864 900 2916
rect 2504 2839 2556 2848
rect 2504 2805 2513 2839
rect 2513 2805 2547 2839
rect 2547 2805 2556 2839
rect 2504 2796 2556 2805
rect 2780 2796 2832 2848
rect 3884 2864 3936 2916
rect 4712 2975 4764 2984
rect 4712 2941 4721 2975
rect 4721 2941 4755 2975
rect 4755 2941 4764 2975
rect 4712 2932 4764 2941
rect 5080 3068 5132 3120
rect 6644 3136 6696 3188
rect 7656 3136 7708 3188
rect 8208 3136 8260 3188
rect 8484 3179 8536 3188
rect 8484 3145 8493 3179
rect 8493 3145 8527 3179
rect 8527 3145 8536 3179
rect 8484 3136 8536 3145
rect 8944 3179 8996 3188
rect 8944 3145 8953 3179
rect 8953 3145 8987 3179
rect 8987 3145 8996 3179
rect 8944 3136 8996 3145
rect 9404 3136 9456 3188
rect 7012 3068 7064 3120
rect 4988 2864 5040 2916
rect 5264 2932 5316 2984
rect 6552 2932 6604 2984
rect 7472 2932 7524 2984
rect 4252 2796 4304 2848
rect 5356 2796 5408 2848
rect 8300 3068 8352 3120
rect 9128 3068 9180 3120
rect 9588 3068 9640 3120
rect 10232 3136 10284 3188
rect 11888 3136 11940 3188
rect 12624 3136 12676 3188
rect 8576 3000 8628 3052
rect 9772 3000 9824 3052
rect 9956 3000 10008 3052
rect 10416 3043 10468 3052
rect 10416 3009 10425 3043
rect 10425 3009 10459 3043
rect 10459 3009 10468 3043
rect 10416 3000 10468 3009
rect 8760 2864 8812 2916
rect 9404 2975 9456 2984
rect 9404 2941 9413 2975
rect 9413 2941 9447 2975
rect 9447 2941 9456 2975
rect 9404 2932 9456 2941
rect 10048 2932 10100 2984
rect 13084 3068 13136 3120
rect 16120 3136 16172 3188
rect 17316 3136 17368 3188
rect 17960 3179 18012 3188
rect 11704 3000 11756 3052
rect 11796 3043 11848 3052
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 13452 3043 13504 3052
rect 11796 3000 11848 3009
rect 13452 3009 13461 3043
rect 13461 3009 13495 3043
rect 13495 3009 13504 3043
rect 13452 3000 13504 3009
rect 13544 3043 13596 3052
rect 13544 3009 13553 3043
rect 13553 3009 13587 3043
rect 13587 3009 13596 3043
rect 13544 3000 13596 3009
rect 13728 3000 13780 3052
rect 14096 3043 14148 3052
rect 14096 3009 14105 3043
rect 14105 3009 14139 3043
rect 14139 3009 14148 3043
rect 14096 3000 14148 3009
rect 15936 3111 15988 3120
rect 15936 3077 15945 3111
rect 15945 3077 15979 3111
rect 15979 3077 15988 3111
rect 15936 3068 15988 3077
rect 14924 3043 14976 3052
rect 12992 2975 13044 2984
rect 12992 2941 13001 2975
rect 13001 2941 13035 2975
rect 13035 2941 13044 2975
rect 12992 2932 13044 2941
rect 14924 3009 14933 3043
rect 14933 3009 14967 3043
rect 14967 3009 14976 3043
rect 14924 3000 14976 3009
rect 15108 3000 15160 3052
rect 17132 3068 17184 3120
rect 17040 3000 17092 3052
rect 17960 3145 17969 3179
rect 17969 3145 18003 3179
rect 18003 3145 18012 3179
rect 17960 3136 18012 3145
rect 19156 3136 19208 3188
rect 19432 3136 19484 3188
rect 19708 3136 19760 3188
rect 18880 3043 18932 3052
rect 14740 2864 14792 2916
rect 15292 2864 15344 2916
rect 16764 2864 16816 2916
rect 17500 2864 17552 2916
rect 17868 2864 17920 2916
rect 18880 3009 18889 3043
rect 18889 3009 18923 3043
rect 18923 3009 18932 3043
rect 18880 3000 18932 3009
rect 19340 3043 19392 3052
rect 19340 3009 19349 3043
rect 19349 3009 19383 3043
rect 19383 3009 19392 3043
rect 19340 3000 19392 3009
rect 19892 3043 19944 3052
rect 19892 3009 19901 3043
rect 19901 3009 19935 3043
rect 19935 3009 19944 3043
rect 19892 3000 19944 3009
rect 20352 3043 20404 3052
rect 20352 3009 20361 3043
rect 20361 3009 20395 3043
rect 20395 3009 20404 3043
rect 20352 3000 20404 3009
rect 20720 3043 20772 3052
rect 20720 3009 20729 3043
rect 20729 3009 20763 3043
rect 20763 3009 20772 3043
rect 20720 3000 20772 3009
rect 19708 2932 19760 2984
rect 18696 2864 18748 2916
rect 19248 2864 19300 2916
rect 9680 2796 9732 2848
rect 13360 2796 13412 2848
rect 13820 2796 13872 2848
rect 14464 2796 14516 2848
rect 16672 2796 16724 2848
rect 17132 2839 17184 2848
rect 17132 2805 17141 2839
rect 17141 2805 17175 2839
rect 17175 2805 17184 2839
rect 17132 2796 17184 2805
rect 18328 2839 18380 2848
rect 18328 2805 18337 2839
rect 18337 2805 18371 2839
rect 18371 2805 18380 2839
rect 18328 2796 18380 2805
rect 21180 2932 21232 2984
rect 19892 2864 19944 2916
rect 20720 2864 20772 2916
rect 22100 2864 22152 2916
rect 20444 2796 20496 2848
rect 21548 2796 21600 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 2228 2592 2280 2644
rect 3424 2524 3476 2576
rect 4252 2592 4304 2644
rect 4804 2635 4856 2644
rect 4804 2601 4813 2635
rect 4813 2601 4847 2635
rect 4847 2601 4856 2635
rect 4804 2592 4856 2601
rect 4896 2592 4948 2644
rect 5356 2592 5408 2644
rect 8576 2592 8628 2644
rect 9496 2592 9548 2644
rect 5540 2524 5592 2576
rect 11152 2592 11204 2644
rect 12440 2592 12492 2644
rect 13728 2592 13780 2644
rect 16672 2592 16724 2644
rect 4712 2456 4764 2508
rect 5356 2456 5408 2508
rect 5632 2456 5684 2508
rect 9220 2456 9272 2508
rect 9680 2499 9732 2508
rect 9680 2465 9689 2499
rect 9689 2465 9723 2499
rect 9723 2465 9732 2499
rect 9680 2456 9732 2465
rect 10140 2456 10192 2508
rect 10784 2456 10836 2508
rect 12440 2499 12492 2508
rect 12440 2465 12449 2499
rect 12449 2465 12483 2499
rect 12483 2465 12492 2499
rect 12440 2456 12492 2465
rect 12900 2456 12952 2508
rect 14188 2524 14240 2576
rect 19248 2524 19300 2576
rect 17684 2456 17736 2508
rect 2228 2431 2280 2440
rect 2228 2397 2237 2431
rect 2237 2397 2271 2431
rect 2271 2397 2280 2431
rect 2228 2388 2280 2397
rect 2320 2431 2372 2440
rect 2320 2397 2329 2431
rect 2329 2397 2363 2431
rect 2363 2397 2372 2431
rect 2320 2388 2372 2397
rect 2872 2388 2924 2440
rect 3148 2388 3200 2440
rect 3884 2388 3936 2440
rect 4068 2388 4120 2440
rect 4528 2388 4580 2440
rect 5448 2388 5500 2440
rect 2504 2295 2556 2304
rect 2504 2261 2513 2295
rect 2513 2261 2547 2295
rect 2547 2261 2556 2295
rect 2504 2252 2556 2261
rect 4252 2252 4304 2304
rect 5908 2320 5960 2372
rect 6828 2388 6880 2440
rect 7748 2388 7800 2440
rect 9864 2388 9916 2440
rect 10876 2388 10928 2440
rect 11060 2431 11112 2440
rect 11060 2397 11069 2431
rect 11069 2397 11103 2431
rect 11103 2397 11112 2431
rect 11060 2388 11112 2397
rect 12348 2431 12400 2440
rect 12348 2397 12357 2431
rect 12357 2397 12391 2431
rect 12391 2397 12400 2431
rect 12348 2388 12400 2397
rect 13360 2431 13412 2440
rect 8208 2320 8260 2372
rect 8392 2320 8444 2372
rect 9588 2320 9640 2372
rect 12164 2320 12216 2372
rect 13360 2397 13369 2431
rect 13369 2397 13403 2431
rect 13403 2397 13412 2431
rect 13360 2388 13412 2397
rect 12808 2320 12860 2372
rect 13636 2320 13688 2372
rect 13820 2388 13872 2440
rect 14464 2431 14516 2440
rect 14464 2397 14473 2431
rect 14473 2397 14507 2431
rect 14507 2397 14516 2431
rect 14464 2388 14516 2397
rect 14740 2388 14792 2440
rect 15292 2388 15344 2440
rect 16120 2431 16172 2440
rect 14556 2320 14608 2372
rect 16120 2397 16129 2431
rect 16129 2397 16163 2431
rect 16163 2397 16172 2431
rect 16120 2388 16172 2397
rect 16948 2388 17000 2440
rect 17132 2388 17184 2440
rect 17500 2431 17552 2440
rect 17500 2397 17509 2431
rect 17509 2397 17543 2431
rect 17543 2397 17552 2431
rect 17500 2388 17552 2397
rect 18328 2388 18380 2440
rect 18696 2431 18748 2440
rect 18696 2397 18705 2431
rect 18705 2397 18739 2431
rect 18739 2397 18748 2431
rect 18696 2388 18748 2397
rect 20260 2456 20312 2508
rect 19892 2431 19944 2440
rect 19892 2397 19901 2431
rect 19901 2397 19935 2431
rect 19935 2397 19944 2431
rect 19892 2388 19944 2397
rect 20720 2431 20772 2440
rect 16764 2320 16816 2372
rect 20720 2397 20729 2431
rect 20729 2397 20763 2431
rect 20763 2397 20772 2431
rect 20720 2388 20772 2397
rect 21180 2431 21232 2440
rect 21180 2397 21189 2431
rect 21189 2397 21223 2431
rect 21223 2397 21232 2431
rect 21180 2388 21232 2397
rect 6736 2295 6788 2304
rect 6736 2261 6745 2295
rect 6745 2261 6779 2295
rect 6779 2261 6788 2295
rect 6736 2252 6788 2261
rect 9220 2295 9272 2304
rect 9220 2261 9229 2295
rect 9229 2261 9263 2295
rect 9263 2261 9272 2295
rect 9220 2252 9272 2261
rect 9496 2252 9548 2304
rect 13268 2252 13320 2304
rect 14280 2252 14332 2304
rect 14740 2252 14792 2304
rect 15108 2252 15160 2304
rect 15568 2252 15620 2304
rect 16028 2252 16080 2304
rect 16396 2252 16448 2304
rect 16948 2252 17000 2304
rect 17408 2252 17460 2304
rect 17868 2252 17920 2304
rect 18328 2252 18380 2304
rect 18788 2252 18840 2304
rect 19708 2252 19760 2304
rect 20260 2252 20312 2304
rect 20628 2252 20680 2304
rect 21088 2252 21140 2304
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
rect 2504 2048 2556 2100
rect 6644 2048 6696 2100
rect 11060 2048 11112 2100
rect 14372 2048 14424 2100
rect 9220 1980 9272 2032
rect 17776 1980 17828 2032
rect 6736 1912 6788 1964
rect 15016 1912 15068 1964
<< metal2 >>
rect 202 22200 258 23000
rect 662 22200 718 23000
rect 1122 22200 1178 23000
rect 1582 22200 1638 23000
rect 2042 22200 2098 23000
rect 2502 22200 2558 23000
rect 2962 22200 3018 23000
rect 3422 22200 3478 23000
rect 3882 22200 3938 23000
rect 4342 22200 4398 23000
rect 4802 22200 4858 23000
rect 5262 22200 5318 23000
rect 5722 22200 5778 23000
rect 6182 22200 6238 23000
rect 6642 22200 6698 23000
rect 7102 22200 7158 23000
rect 7562 22200 7618 23000
rect 8022 22200 8078 23000
rect 8482 22200 8538 23000
rect 8942 22200 8998 23000
rect 9402 22200 9458 23000
rect 9862 22200 9918 23000
rect 10322 22200 10378 23000
rect 10782 22200 10838 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12162 22200 12218 23000
rect 12622 22200 12678 23000
rect 12728 22222 13032 22250
rect 216 19310 244 22200
rect 204 19304 256 19310
rect 204 19246 256 19252
rect 676 18834 704 22200
rect 1136 19242 1164 22200
rect 1492 20256 1544 20262
rect 1490 20224 1492 20233
rect 1544 20224 1546 20233
rect 1490 20159 1546 20168
rect 1596 19786 1624 22200
rect 1858 20632 1914 20641
rect 2056 20618 2084 22200
rect 2226 21040 2282 21049
rect 2226 20975 2282 20984
rect 2056 20590 2176 20618
rect 2240 20602 2268 20975
rect 1858 20567 1860 20576
rect 1912 20567 1914 20576
rect 1860 20538 1912 20544
rect 1768 20460 1820 20466
rect 1768 20402 1820 20408
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 1676 19848 1728 19854
rect 1676 19790 1728 19796
rect 1584 19780 1636 19786
rect 1584 19722 1636 19728
rect 1492 19712 1544 19718
rect 1492 19654 1544 19660
rect 1504 19417 1532 19654
rect 1490 19408 1546 19417
rect 1490 19343 1546 19352
rect 1124 19236 1176 19242
rect 1124 19178 1176 19184
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1504 19009 1532 19110
rect 1490 19000 1546 19009
rect 1490 18935 1546 18944
rect 1688 18850 1716 19790
rect 664 18828 716 18834
rect 664 18770 716 18776
rect 1596 18822 1716 18850
rect 1492 18624 1544 18630
rect 1490 18592 1492 18601
rect 1544 18592 1546 18601
rect 1490 18527 1546 18536
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1504 17785 1532 18022
rect 1490 17776 1546 17785
rect 1490 17711 1546 17720
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 17377 1532 17478
rect 1490 17368 1546 17377
rect 1490 17303 1546 17312
rect 1596 16998 1624 18822
rect 1676 18760 1728 18766
rect 1676 18702 1728 18708
rect 1688 18057 1716 18702
rect 1674 18048 1730 18057
rect 1674 17983 1730 17992
rect 1780 17338 1808 20402
rect 1858 19816 1914 19825
rect 1858 19751 1914 19760
rect 1872 19718 1900 19751
rect 1860 19712 1912 19718
rect 1860 19654 1912 19660
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1964 19417 1992 19450
rect 1950 19408 2006 19417
rect 1860 19372 1912 19378
rect 1950 19343 2006 19352
rect 1860 19314 1912 19320
rect 1872 19242 1900 19314
rect 1860 19236 1912 19242
rect 1860 19178 1912 19184
rect 2056 18426 2084 20402
rect 2148 19990 2176 20590
rect 2228 20596 2280 20602
rect 2228 20538 2280 20544
rect 2516 20466 2544 22200
rect 2976 20602 3004 22200
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 3436 20466 3464 22200
rect 3896 20466 3924 22200
rect 4160 20596 4212 20602
rect 4160 20538 4212 20544
rect 2412 20460 2464 20466
rect 2412 20402 2464 20408
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 3424 20460 3476 20466
rect 3424 20402 3476 20408
rect 3884 20460 3936 20466
rect 3884 20402 3936 20408
rect 2424 20058 2452 20402
rect 2412 20052 2464 20058
rect 2412 19994 2464 20000
rect 2136 19984 2188 19990
rect 2136 19926 2188 19932
rect 2148 19854 2176 19926
rect 2136 19848 2188 19854
rect 2136 19790 2188 19796
rect 2320 19712 2372 19718
rect 2318 19680 2320 19689
rect 2372 19680 2374 19689
rect 2318 19615 2374 19624
rect 2516 19514 2544 20402
rect 3436 20058 3464 20402
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3896 20058 3924 20402
rect 3976 20256 4028 20262
rect 3976 20198 4028 20204
rect 3424 20052 3476 20058
rect 3424 19994 3476 20000
rect 3884 20052 3936 20058
rect 3884 19994 3936 20000
rect 2596 19916 2648 19922
rect 2596 19858 2648 19864
rect 2504 19508 2556 19514
rect 2504 19450 2556 19456
rect 2044 18420 2096 18426
rect 2044 18362 2096 18368
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 2228 18284 2280 18290
rect 2228 18226 2280 18232
rect 1858 18184 1914 18193
rect 1858 18119 1860 18128
rect 1912 18119 1914 18128
rect 1860 18090 1912 18096
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1492 16992 1544 16998
rect 1490 16960 1492 16969
rect 1584 16992 1636 16998
rect 1544 16960 1546 16969
rect 1584 16934 1636 16940
rect 1490 16895 1546 16904
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 1504 16153 1532 16390
rect 1490 16144 1546 16153
rect 1490 16079 1546 16088
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 15745 1532 15846
rect 1490 15736 1546 15745
rect 1490 15671 1546 15680
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 12968 1440 15438
rect 1492 15360 1544 15366
rect 1490 15328 1492 15337
rect 1544 15328 1546 15337
rect 1490 15263 1546 15272
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1504 14521 1532 14758
rect 1490 14512 1546 14521
rect 1490 14447 1546 14456
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1504 14113 1532 14214
rect 1490 14104 1546 14113
rect 1490 14039 1546 14048
rect 1492 13728 1544 13734
rect 1490 13696 1492 13705
rect 1544 13696 1546 13705
rect 1490 13631 1546 13640
rect 1490 13288 1546 13297
rect 1490 13223 1546 13232
rect 1504 13190 1532 13223
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 1412 12940 1532 12968
rect 1398 12880 1454 12889
rect 1398 12815 1400 12824
rect 1452 12815 1454 12824
rect 1400 12786 1452 12792
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1412 12073 1440 12174
rect 1398 12064 1454 12073
rect 1398 11999 1454 12008
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1412 11665 1440 11698
rect 1398 11656 1454 11665
rect 1398 11591 1454 11600
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10849 1440 11086
rect 1398 10840 1454 10849
rect 1398 10775 1454 10784
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1412 10441 1440 10610
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 1400 10056 1452 10062
rect 1398 10024 1400 10033
rect 1452 10024 1454 10033
rect 1398 9959 1454 9968
rect 1412 9722 1440 9959
rect 1400 9716 1452 9722
rect 1400 9658 1452 9664
rect 1504 9450 1532 12940
rect 1596 12442 1624 16526
rect 1688 15706 1716 17138
rect 1858 16552 1914 16561
rect 1858 16487 1914 16496
rect 1872 16454 1900 16487
rect 1860 16448 1912 16454
rect 1860 16390 1912 16396
rect 1964 15706 1992 18226
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 2056 15162 2084 16526
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1688 12481 1716 12786
rect 1674 12472 1730 12481
rect 1584 12436 1636 12442
rect 1674 12407 1730 12416
rect 1584 12378 1636 12384
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1596 10606 1624 11494
rect 1688 11257 1716 11698
rect 1780 11354 1808 14962
rect 1858 14920 1914 14929
rect 1858 14855 1860 14864
rect 1912 14855 1914 14864
rect 1860 14826 1912 14832
rect 1860 14408 1912 14414
rect 1860 14350 1912 14356
rect 1768 11348 1820 11354
rect 1768 11290 1820 11296
rect 1674 11248 1730 11257
rect 1674 11183 1730 11192
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1596 10033 1624 10406
rect 1676 10056 1728 10062
rect 1582 10024 1638 10033
rect 1676 9998 1728 10004
rect 1582 9959 1638 9968
rect 1688 9625 1716 9998
rect 1674 9616 1730 9625
rect 1674 9551 1730 9560
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 1492 9444 1544 9450
rect 1492 9386 1544 9392
rect 1398 9208 1454 9217
rect 1398 9143 1454 9152
rect 1412 8974 1440 9143
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1688 8809 1716 8910
rect 1674 8800 1730 8809
rect 1674 8735 1730 8744
rect 1688 8634 1716 8735
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8401 1440 8434
rect 1398 8392 1454 8401
rect 1454 8350 1624 8378
rect 1398 8327 1454 8336
rect 1398 7984 1454 7993
rect 1398 7919 1454 7928
rect 1412 7886 1440 7919
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 7698 1440 7822
rect 1412 7670 1532 7698
rect 1398 7576 1454 7585
rect 1504 7546 1532 7670
rect 1398 7511 1454 7520
rect 1492 7540 1544 7546
rect 1412 7410 1440 7511
rect 1492 7482 1544 7488
rect 1596 7478 1624 8350
rect 1780 8090 1808 9522
rect 1872 9450 1900 14350
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1964 9450 1992 13874
rect 2056 10266 2084 14962
rect 2148 11354 2176 16050
rect 2240 15162 2268 18226
rect 2504 17672 2556 17678
rect 2504 17614 2556 17620
rect 2516 15706 2544 17614
rect 2608 17338 2636 19858
rect 2688 19712 2740 19718
rect 2688 19654 2740 19660
rect 2700 19553 2728 19654
rect 2686 19544 2742 19553
rect 2686 19479 2742 19488
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 2700 17338 2728 19314
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 2872 18284 2924 18290
rect 2872 18226 2924 18232
rect 2596 17332 2648 17338
rect 2596 17274 2648 17280
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 2884 16250 2912 18226
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 3516 17196 3568 17202
rect 3516 17138 3568 17144
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 2976 16794 3004 17070
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 3068 16250 3096 17138
rect 3528 17082 3556 17138
rect 3436 17054 3556 17082
rect 3436 16794 3464 17054
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 3056 16244 3108 16250
rect 3056 16186 3108 16192
rect 3160 16114 3188 16390
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 2228 15156 2280 15162
rect 2228 15098 2280 15104
rect 2884 14890 2912 15302
rect 3896 15162 3924 15302
rect 3884 15156 3936 15162
rect 3884 15098 3936 15104
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 3424 14952 3476 14958
rect 3988 14906 4016 20198
rect 4172 17270 4200 20538
rect 4356 20466 4384 22200
rect 4816 20466 4844 22200
rect 4344 20460 4396 20466
rect 4344 20402 4396 20408
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 4356 20058 4384 20402
rect 4436 20324 4488 20330
rect 4436 20266 4488 20272
rect 4344 20052 4396 20058
rect 4344 19994 4396 20000
rect 4342 19544 4398 19553
rect 4342 19479 4398 19488
rect 4250 19408 4306 19417
rect 4250 19343 4306 19352
rect 4160 17264 4212 17270
rect 4160 17206 4212 17212
rect 4264 16658 4292 19343
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 4356 16590 4384 19479
rect 4448 17338 4476 20266
rect 4816 20058 4844 20402
rect 4988 20392 5040 20398
rect 4988 20334 5040 20340
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 5000 19417 5028 20334
rect 5276 20058 5304 22200
rect 5736 20466 5764 22200
rect 6196 20856 6224 22200
rect 6012 20828 6224 20856
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 5264 20052 5316 20058
rect 5264 19994 5316 20000
rect 5276 19854 5304 19994
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 5540 19712 5592 19718
rect 5592 19672 5672 19700
rect 5540 19654 5592 19660
rect 4986 19408 5042 19417
rect 4986 19343 5042 19352
rect 5540 19236 5592 19242
rect 5540 19178 5592 19184
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 5264 18352 5316 18358
rect 5264 18294 5316 18300
rect 4988 18216 5040 18222
rect 4988 18158 5040 18164
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4436 17332 4488 17338
rect 4488 17292 4568 17320
rect 4436 17274 4488 17280
rect 4436 17128 4488 17134
rect 4436 17070 4488 17076
rect 4448 16726 4476 17070
rect 4436 16720 4488 16726
rect 4436 16662 4488 16668
rect 4160 16584 4212 16590
rect 4158 16552 4160 16561
rect 4344 16584 4396 16590
rect 4212 16552 4214 16561
rect 4344 16526 4396 16532
rect 4158 16487 4214 16496
rect 4356 16130 4384 16526
rect 4172 16102 4384 16130
rect 4068 15564 4120 15570
rect 4068 15506 4120 15512
rect 3424 14894 3476 14900
rect 2872 14884 2924 14890
rect 2872 14826 2924 14832
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2320 10600 2372 10606
rect 2320 10542 2372 10548
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 1952 9444 2004 9450
rect 1952 9386 2004 9392
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1964 8480 1992 8774
rect 2056 8634 2084 9522
rect 2148 9178 2176 9522
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 2044 8492 2096 8498
rect 1964 8452 2044 8480
rect 2044 8434 2096 8440
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1584 7472 1636 7478
rect 1584 7414 1636 7420
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1412 7002 1440 7346
rect 1582 7304 1638 7313
rect 1582 7239 1584 7248
rect 1636 7239 1638 7248
rect 1584 7210 1636 7216
rect 1688 7177 1716 7346
rect 1674 7168 1730 7177
rect 1674 7103 1730 7112
rect 1400 6996 1452 7002
rect 1400 6938 1452 6944
rect 1400 6792 1452 6798
rect 1398 6760 1400 6769
rect 1676 6792 1728 6798
rect 1452 6760 1454 6769
rect 1676 6734 1728 6740
rect 1398 6695 1454 6704
rect 1688 6361 1716 6734
rect 1674 6352 1730 6361
rect 1400 6316 1452 6322
rect 1674 6287 1730 6296
rect 1400 6258 1452 6264
rect 1412 5953 1440 6258
rect 1398 5944 1454 5953
rect 1398 5879 1400 5888
rect 1452 5879 1454 5888
rect 1400 5850 1452 5856
rect 1412 5819 1440 5850
rect 1584 5840 1636 5846
rect 1582 5808 1584 5817
rect 1636 5808 1638 5817
rect 1582 5743 1638 5752
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1412 5545 1440 5646
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 1504 4729 1532 5170
rect 1688 5137 1716 5646
rect 1674 5128 1730 5137
rect 1674 5063 1730 5072
rect 1490 4720 1546 4729
rect 1490 4655 1546 4664
rect 1964 4146 1992 7686
rect 2056 6458 2084 8434
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2148 6390 2176 8366
rect 2240 6769 2268 9454
rect 2226 6760 2282 6769
rect 2226 6695 2282 6704
rect 2136 6384 2188 6390
rect 2136 6326 2188 6332
rect 2044 6248 2096 6254
rect 2044 6190 2096 6196
rect 2056 5166 2084 6190
rect 2240 5760 2268 6695
rect 2148 5732 2268 5760
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 2056 5030 2084 5102
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 1308 3936 1360 3942
rect 1308 3878 1360 3884
rect 388 3732 440 3738
rect 388 3674 440 3680
rect 400 800 428 3674
rect 1320 3466 1348 3878
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1492 3528 1544 3534
rect 1490 3496 1492 3505
rect 1688 3505 1716 3606
rect 1544 3496 1546 3505
rect 1308 3460 1360 3466
rect 1490 3431 1546 3440
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 1860 3460 1912 3466
rect 1308 3402 1360 3408
rect 1860 3402 1912 3408
rect 848 2916 900 2922
rect 848 2858 900 2864
rect 860 800 888 2858
rect 1320 800 1348 3402
rect 1872 3097 1900 3402
rect 1858 3088 1914 3097
rect 1768 3052 1820 3058
rect 1858 3023 1914 3032
rect 1768 2994 1820 3000
rect 1780 800 1808 2994
rect 2056 2990 2084 4082
rect 2148 3754 2176 5732
rect 2228 5568 2280 5574
rect 2228 5510 2280 5516
rect 2240 5370 2268 5510
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2332 5302 2360 10542
rect 2700 9926 2728 12038
rect 2884 10169 2912 14826
rect 2976 11898 3004 14894
rect 3436 14346 3464 14894
rect 3896 14878 4016 14906
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3424 14340 3476 14346
rect 3424 14282 3476 14288
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3160 12986 3188 13262
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2870 10160 2926 10169
rect 2870 10095 2926 10104
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2410 9480 2466 9489
rect 2410 9415 2412 9424
rect 2464 9415 2466 9424
rect 2504 9444 2556 9450
rect 2412 9386 2464 9392
rect 2504 9386 2556 9392
rect 2516 8974 2544 9386
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2608 8974 2636 9114
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2412 8016 2464 8022
rect 2412 7958 2464 7964
rect 2424 7546 2452 7958
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2410 7440 2466 7449
rect 2410 7375 2466 7384
rect 2320 5296 2372 5302
rect 2320 5238 2372 5244
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 2240 4321 2268 4558
rect 2226 4312 2282 4321
rect 2226 4247 2282 4256
rect 2228 4072 2280 4078
rect 2228 4014 2280 4020
rect 2240 3913 2268 4014
rect 2226 3904 2282 3913
rect 2226 3839 2282 3848
rect 2148 3726 2268 3754
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 2148 2990 2176 3130
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 2148 1873 2176 2926
rect 2240 2650 2268 3726
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2332 3534 2360 3674
rect 2424 3670 2452 7375
rect 2516 6662 2544 8774
rect 2608 7886 2636 8910
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2700 7818 2728 9862
rect 2792 9722 2820 9862
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2792 8906 2820 9318
rect 2976 9110 3004 10406
rect 3068 9178 3096 11018
rect 3148 10736 3200 10742
rect 3148 10678 3200 10684
rect 3160 10266 3188 10678
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3146 10160 3202 10169
rect 3146 10095 3202 10104
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 2964 9104 3016 9110
rect 2964 9046 3016 9052
rect 2780 8900 2832 8906
rect 2780 8842 2832 8848
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2792 8362 2820 8570
rect 3160 8498 3188 10095
rect 3252 8537 3280 12174
rect 3436 10266 3464 14282
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3896 12850 3924 14878
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3988 12889 4016 14758
rect 3974 12880 4030 12889
rect 3884 12844 3936 12850
rect 3974 12815 4030 12824
rect 3884 12786 3936 12792
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 4080 12442 4108 15506
rect 4172 14414 4200 16102
rect 4436 15496 4488 15502
rect 4436 15438 4488 15444
rect 4252 15428 4304 15434
rect 4252 15370 4304 15376
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4264 12986 4292 15370
rect 4344 15088 4396 15094
rect 4344 15030 4396 15036
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 4172 12646 4200 12854
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 4172 11286 4200 11698
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3424 10260 3476 10266
rect 3344 10220 3424 10248
rect 3344 10130 3372 10220
rect 3424 10202 3476 10208
rect 3790 10160 3846 10169
rect 3332 10124 3384 10130
rect 3790 10095 3792 10104
rect 3332 10066 3384 10072
rect 3844 10095 3846 10104
rect 3792 10066 3844 10072
rect 3344 9178 3372 10066
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3436 9178 3464 9998
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3238 8528 3294 8537
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 3148 8492 3200 8498
rect 3238 8463 3294 8472
rect 3148 8434 3200 8440
rect 2884 8401 2912 8434
rect 2870 8392 2926 8401
rect 2780 8356 2832 8362
rect 2870 8327 2926 8336
rect 2780 8298 2832 8304
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 3896 8090 3924 11086
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4080 10130 4108 10542
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3988 8634 4016 9998
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 4080 7857 4108 8910
rect 4172 8634 4200 10610
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4066 7848 4122 7857
rect 2688 7812 2740 7818
rect 4066 7783 4122 7792
rect 2688 7754 2740 7760
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 4068 6860 4120 6866
rect 4120 6820 4200 6848
rect 4068 6802 4120 6808
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 2778 6352 2834 6361
rect 2778 6287 2834 6296
rect 2792 5522 2820 6287
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 2700 5494 2820 5522
rect 2596 4208 2648 4214
rect 2596 4150 2648 4156
rect 2608 3670 2636 4150
rect 2700 4146 2728 5494
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2412 3664 2464 3670
rect 2596 3664 2648 3670
rect 2412 3606 2464 3612
rect 2502 3632 2558 3641
rect 2596 3606 2648 3612
rect 2792 3602 2820 3878
rect 2502 3567 2558 3576
rect 2780 3596 2832 3602
rect 2320 3528 2372 3534
rect 2320 3470 2372 3476
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2332 3097 2360 3334
rect 2318 3088 2374 3097
rect 2318 3023 2374 3032
rect 2320 2984 2372 2990
rect 2320 2926 2372 2932
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 2332 2446 2360 2926
rect 2516 2854 2544 3567
rect 2780 3538 2832 3544
rect 2780 3392 2832 3398
rect 2700 3352 2780 3380
rect 2700 3058 2728 3352
rect 2780 3334 2832 3340
rect 2780 3188 2832 3194
rect 2976 3176 3004 3878
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 3988 3670 4016 6598
rect 4172 6254 4200 6820
rect 4160 6248 4212 6254
rect 4160 6190 4212 6196
rect 4264 4758 4292 11018
rect 4356 10266 4384 15030
rect 4448 13530 4476 15438
rect 4540 15434 4568 17292
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 4632 16674 4660 17206
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4724 16794 4752 17138
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4632 16646 4752 16674
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4632 15502 4660 16526
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4528 15428 4580 15434
rect 4528 15370 4580 15376
rect 4528 14952 4580 14958
rect 4528 14894 4580 14900
rect 4540 14278 4568 14894
rect 4632 14890 4660 15438
rect 4620 14884 4672 14890
rect 4620 14826 4672 14832
rect 4618 14648 4674 14657
rect 4618 14583 4674 14592
rect 4632 14482 4660 14583
rect 4724 14550 4752 16646
rect 4816 15094 4844 17614
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4908 17338 4936 17478
rect 4896 17332 4948 17338
rect 4896 17274 4948 17280
rect 5000 16726 5028 18158
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5184 17649 5212 17682
rect 5170 17640 5226 17649
rect 5170 17575 5226 17584
rect 5184 17134 5212 17575
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 4988 16720 5040 16726
rect 4988 16662 5040 16668
rect 4896 15904 4948 15910
rect 4896 15846 4948 15852
rect 4908 15638 4936 15846
rect 4896 15632 4948 15638
rect 4896 15574 4948 15580
rect 4804 15088 4856 15094
rect 4804 15030 4856 15036
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 4908 14618 4936 14894
rect 4896 14612 4948 14618
rect 4896 14554 4948 14560
rect 4712 14544 4764 14550
rect 5000 14498 5028 16662
rect 5276 16153 5304 18294
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5368 17746 5396 18022
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 5460 17678 5488 18566
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5262 16144 5318 16153
rect 5080 16108 5132 16114
rect 5262 16079 5318 16088
rect 5080 16050 5132 16056
rect 5092 15609 5120 16050
rect 5172 15972 5224 15978
rect 5172 15914 5224 15920
rect 5184 15706 5212 15914
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5078 15600 5134 15609
rect 5276 15570 5304 16079
rect 5368 15910 5396 16730
rect 5552 16538 5580 19178
rect 5460 16510 5580 16538
rect 5460 15994 5488 16510
rect 5460 15966 5580 15994
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 5368 15570 5396 15846
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 5078 15535 5134 15544
rect 5264 15564 5316 15570
rect 5264 15506 5316 15512
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 4712 14486 4764 14492
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4816 14470 5028 14498
rect 5080 14476 5132 14482
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4528 12708 4580 12714
rect 4528 12650 4580 12656
rect 4540 12434 4568 12650
rect 4448 12406 4568 12434
rect 4448 10674 4476 12406
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4436 10668 4488 10674
rect 4436 10610 4488 10616
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4448 9654 4476 9862
rect 4436 9648 4488 9654
rect 4436 9590 4488 9596
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4356 8430 4384 8978
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4448 6798 4476 9590
rect 4540 9382 4568 11494
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 4540 4554 4568 9318
rect 4632 6458 4660 11018
rect 4816 10538 4844 14470
rect 5080 14418 5132 14424
rect 5092 14385 5120 14418
rect 5264 14408 5316 14414
rect 5078 14376 5134 14385
rect 5264 14350 5316 14356
rect 5078 14311 5134 14320
rect 5276 14006 5304 14350
rect 5368 14074 5396 14894
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5264 14000 5316 14006
rect 5264 13942 5316 13948
rect 5460 13938 5488 15574
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5552 13870 5580 15966
rect 5644 15570 5672 19672
rect 5736 19514 5764 20402
rect 5816 20324 5868 20330
rect 5816 20266 5868 20272
rect 5724 19508 5776 19514
rect 5724 19450 5776 19456
rect 5722 19408 5778 19417
rect 5722 19343 5778 19352
rect 5736 18358 5764 19343
rect 5828 18426 5856 20266
rect 5908 20256 5960 20262
rect 5908 20198 5960 20204
rect 5920 18426 5948 20198
rect 6012 20058 6040 20828
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 6656 20398 6684 22200
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 6644 20392 6696 20398
rect 6644 20334 6696 20340
rect 6000 20052 6052 20058
rect 6000 19994 6052 20000
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 6564 19417 6592 19790
rect 6656 19786 6684 20334
rect 6736 20256 6788 20262
rect 6736 20198 6788 20204
rect 6644 19780 6696 19786
rect 6644 19722 6696 19728
rect 6550 19408 6606 19417
rect 6000 19372 6052 19378
rect 6550 19343 6606 19352
rect 6000 19314 6052 19320
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 5724 18352 5776 18358
rect 5724 18294 5776 18300
rect 5828 17626 5856 18362
rect 6012 17746 6040 19314
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 6000 17740 6052 17746
rect 6000 17682 6052 17688
rect 6552 17672 6604 17678
rect 5828 17598 6040 17626
rect 6552 17614 6604 17620
rect 5724 17536 5776 17542
rect 5724 17478 5776 17484
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5736 17270 5764 17478
rect 5816 17332 5868 17338
rect 5920 17320 5948 17478
rect 5868 17292 5948 17320
rect 5816 17274 5868 17280
rect 5724 17264 5776 17270
rect 5724 17206 5776 17212
rect 5724 17128 5776 17134
rect 5724 17070 5776 17076
rect 5736 15638 5764 17070
rect 6012 16538 6040 17598
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 6182 17096 6238 17105
rect 6182 17031 6238 17040
rect 6196 16658 6224 17031
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 5828 16510 6040 16538
rect 5724 15632 5776 15638
rect 5724 15574 5776 15580
rect 5632 15564 5684 15570
rect 5632 15506 5684 15512
rect 5828 15162 5856 16510
rect 5908 16448 5960 16454
rect 5908 16390 5960 16396
rect 6000 16448 6052 16454
rect 6000 16390 6052 16396
rect 5920 16250 5948 16390
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 5906 16144 5962 16153
rect 6012 16130 6040 16390
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6564 16182 6592 17614
rect 6748 16402 6776 20198
rect 6656 16374 6776 16402
rect 6368 16176 6420 16182
rect 6012 16102 6132 16130
rect 6368 16118 6420 16124
rect 6552 16176 6604 16182
rect 6552 16118 6604 16124
rect 5906 16079 5908 16088
rect 5960 16079 5962 16088
rect 5908 16050 5960 16056
rect 6000 15972 6052 15978
rect 6000 15914 6052 15920
rect 5908 15904 5960 15910
rect 5908 15846 5960 15852
rect 5816 15156 5868 15162
rect 5816 15098 5868 15104
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4908 11082 4936 12582
rect 5000 12442 5028 12786
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 5000 11150 5028 11630
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4710 10432 4766 10441
rect 4710 10367 4766 10376
rect 4724 10169 4752 10367
rect 4908 10198 4936 10542
rect 4896 10192 4948 10198
rect 4710 10160 4766 10169
rect 4896 10134 4948 10140
rect 4710 10095 4766 10104
rect 4724 10062 4752 10095
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4816 6866 4844 9454
rect 4908 8974 4936 10134
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5000 9489 5028 9998
rect 4986 9480 5042 9489
rect 4986 9415 5042 9424
rect 5092 9042 5120 12038
rect 5184 10810 5212 13806
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5262 13288 5318 13297
rect 5262 13223 5318 13232
rect 5276 12782 5304 13223
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5276 10810 5304 11290
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 4988 8016 5040 8022
rect 4988 7958 5040 7964
rect 4908 7410 4936 7958
rect 5000 7750 5028 7958
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4988 7336 5040 7342
rect 4988 7278 5040 7284
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4724 6254 4752 6598
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4724 5574 4752 6190
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4620 5296 4672 5302
rect 4724 5273 4752 5510
rect 4620 5238 4672 5244
rect 4710 5264 4766 5273
rect 4528 4548 4580 4554
rect 4528 4490 4580 4496
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 2832 3148 3004 3176
rect 2780 3130 2832 3136
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2792 2854 2820 2994
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2792 2689 2820 2790
rect 3160 2774 3188 3334
rect 2884 2746 3188 2774
rect 2778 2680 2834 2689
rect 2778 2615 2834 2624
rect 2884 2446 2912 2746
rect 3436 2582 3464 3334
rect 4080 3194 4108 4082
rect 4252 4004 4304 4010
rect 4252 3946 4304 3952
rect 4264 3602 4292 3946
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4264 3194 4292 3334
rect 4632 3194 4660 5238
rect 4710 5199 4766 5208
rect 4712 5092 4764 5098
rect 4712 5034 4764 5040
rect 4724 4826 4752 5034
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 3884 2916 3936 2922
rect 3884 2858 3936 2864
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 3424 2576 3476 2582
rect 3424 2518 3476 2524
rect 3896 2446 3924 2858
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4264 2650 4292 2790
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2872 2440 2924 2446
rect 2872 2382 2924 2388
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 2240 2281 2268 2382
rect 2226 2272 2282 2281
rect 2226 2207 2282 2216
rect 2134 1864 2190 1873
rect 2134 1799 2190 1808
rect 2332 1714 2360 2382
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 2516 2106 2544 2246
rect 2504 2100 2556 2106
rect 2504 2042 2556 2048
rect 2884 1986 2912 2382
rect 2240 1686 2360 1714
rect 2700 1958 2912 1986
rect 2240 800 2268 1686
rect 2700 800 2728 1958
rect 3160 800 3188 2382
rect 3620 870 3740 898
rect 3620 800 3648 870
rect 386 0 442 800
rect 846 0 902 800
rect 1306 0 1362 800
rect 1766 0 1822 800
rect 2226 0 2282 800
rect 2686 0 2742 800
rect 3146 0 3202 800
rect 3606 0 3662 800
rect 3712 762 3740 870
rect 3896 762 3924 2382
rect 4080 800 4108 2382
rect 4252 2304 4304 2310
rect 4356 2292 4384 3130
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4724 2514 4752 2926
rect 4816 2650 4844 5578
rect 4908 2650 4936 6802
rect 5000 6662 5028 7278
rect 5092 7274 5120 8978
rect 5184 8906 5212 9386
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5170 8392 5226 8401
rect 5170 8327 5172 8336
rect 5224 8327 5226 8336
rect 5172 8298 5224 8304
rect 5172 7812 5224 7818
rect 5172 7754 5224 7760
rect 5184 7274 5212 7754
rect 5276 7478 5304 10746
rect 5368 9518 5396 13398
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5460 11218 5488 11766
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5460 9654 5488 11154
rect 5552 9654 5580 13806
rect 5644 13530 5672 14214
rect 5736 14074 5764 14962
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5828 14550 5856 14758
rect 5816 14544 5868 14550
rect 5816 14486 5868 14492
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5724 13252 5776 13258
rect 5724 13194 5776 13200
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5644 11082 5672 12242
rect 5736 11354 5764 13194
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5722 11248 5778 11257
rect 5722 11183 5778 11192
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5736 10606 5764 11183
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5644 9897 5672 10066
rect 5630 9888 5686 9897
rect 5630 9823 5686 9832
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5460 9178 5488 9454
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5264 7472 5316 7478
rect 5264 7414 5316 7420
rect 5080 7268 5132 7274
rect 5080 7210 5132 7216
rect 5172 7268 5224 7274
rect 5172 7210 5224 7216
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 5000 5574 5028 6598
rect 5264 6180 5316 6186
rect 5264 6122 5316 6128
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 5000 5166 5028 5510
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5092 5098 5120 5782
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 5184 4690 5212 5646
rect 5276 5370 5304 6122
rect 5368 5778 5396 8774
rect 5460 8294 5488 9114
rect 5552 8430 5580 9318
rect 5736 9042 5764 10542
rect 5828 10266 5856 12786
rect 5920 11218 5948 15846
rect 6012 15706 6040 15914
rect 6104 15706 6132 16102
rect 6380 15910 6408 16118
rect 6368 15904 6420 15910
rect 6366 15872 6368 15881
rect 6420 15872 6422 15881
rect 6366 15807 6422 15816
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 6380 15638 6408 15807
rect 6368 15632 6420 15638
rect 6368 15574 6420 15580
rect 6564 15434 6592 16118
rect 6552 15428 6604 15434
rect 6552 15370 6604 15376
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 6012 14822 6040 15302
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 6012 12374 6040 14758
rect 6274 14512 6330 14521
rect 6274 14447 6330 14456
rect 6288 14414 6316 14447
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6564 14074 6592 14214
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6458 13968 6514 13977
rect 6458 13903 6514 13912
rect 6182 13560 6238 13569
rect 6182 13495 6238 13504
rect 6196 13394 6224 13495
rect 6472 13394 6500 13903
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 6460 13388 6512 13394
rect 6460 13330 6512 13336
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 6550 13016 6606 13025
rect 6460 12980 6512 12986
rect 6550 12951 6606 12960
rect 6460 12922 6512 12928
rect 6276 12776 6328 12782
rect 6276 12718 6328 12724
rect 6000 12368 6052 12374
rect 6000 12310 6052 12316
rect 6288 12306 6316 12718
rect 6472 12628 6500 12922
rect 6564 12782 6592 12951
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6472 12600 6592 12628
rect 6564 12345 6592 12600
rect 6550 12336 6606 12345
rect 6276 12300 6328 12306
rect 6656 12306 6684 16374
rect 6734 16280 6790 16289
rect 6734 16215 6790 16224
rect 6748 15570 6776 16215
rect 6736 15564 6788 15570
rect 6736 15506 6788 15512
rect 6840 15094 6868 20538
rect 7116 20466 7144 22200
rect 7576 20466 7604 22200
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7564 20460 7616 20466
rect 7564 20402 7616 20408
rect 7012 20392 7064 20398
rect 7012 20334 7064 20340
rect 7024 19417 7052 20334
rect 7116 20058 7144 20402
rect 7470 20360 7526 20369
rect 7380 20324 7432 20330
rect 7470 20295 7526 20304
rect 7380 20266 7432 20272
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7010 19408 7066 19417
rect 7010 19343 7066 19352
rect 7116 19174 7144 19790
rect 7196 19236 7248 19242
rect 7196 19178 7248 19184
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 6920 18896 6972 18902
rect 6920 18838 6972 18844
rect 6932 18358 6960 18838
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 6932 17882 6960 18294
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6918 17776 6974 17785
rect 6918 17711 6974 17720
rect 6932 17134 6960 17711
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 6932 16266 6960 17070
rect 6932 16238 7052 16266
rect 6918 16144 6974 16153
rect 6918 16079 6974 16088
rect 6932 15978 6960 16079
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 7024 15858 7052 16238
rect 6932 15830 7052 15858
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 6932 14958 6960 15830
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6736 14952 6788 14958
rect 6736 14894 6788 14900
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6748 14822 6776 14894
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6748 14074 6776 14758
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6734 13560 6790 13569
rect 6734 13495 6790 13504
rect 6748 12986 6776 13495
rect 6840 13258 6868 14826
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6932 13138 6960 13806
rect 6840 13110 6960 13138
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6840 12866 6868 13110
rect 6748 12838 6868 12866
rect 6550 12271 6606 12280
rect 6644 12300 6696 12306
rect 6276 12242 6328 12248
rect 6644 12242 6696 12248
rect 6748 12220 6776 12838
rect 6920 12640 6972 12646
rect 6826 12608 6882 12617
rect 6920 12582 6972 12588
rect 6826 12543 6882 12552
rect 6840 12442 6868 12543
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6748 12192 6868 12220
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6734 12064 6790 12073
rect 6012 11354 6040 12038
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 6564 11898 6592 12038
rect 6734 11999 6790 12008
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6092 11756 6144 11762
rect 6092 11698 6144 11704
rect 6104 11558 6132 11698
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6104 11234 6132 11494
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 6012 11206 6132 11234
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5920 9625 5948 9862
rect 5906 9616 5962 9625
rect 5816 9580 5868 9586
rect 5906 9551 5962 9560
rect 5816 9522 5868 9528
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5724 8832 5776 8838
rect 5644 8792 5724 8820
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5460 7478 5488 7890
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5552 7342 5580 8366
rect 5644 7546 5672 8792
rect 5724 8774 5776 8780
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5736 8090 5764 8366
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5722 7984 5778 7993
rect 5722 7919 5724 7928
rect 5776 7919 5778 7928
rect 5724 7890 5776 7896
rect 5632 7540 5684 7546
rect 5828 7528 5856 9522
rect 6012 9353 6040 11206
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6090 10160 6146 10169
rect 6090 10095 6092 10104
rect 6144 10095 6146 10104
rect 6092 10066 6144 10072
rect 6472 9926 6500 10542
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6092 9648 6144 9654
rect 6092 9590 6144 9596
rect 5998 9344 6054 9353
rect 5998 9279 6054 9288
rect 6104 9194 6132 9590
rect 6012 9166 6132 9194
rect 6564 9178 6592 10950
rect 6656 10810 6684 10950
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6642 10704 6698 10713
rect 6642 10639 6698 10648
rect 6656 10130 6684 10639
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6748 9382 6776 11999
rect 6840 10606 6868 12192
rect 6932 11830 6960 12582
rect 6920 11824 6972 11830
rect 6920 11766 6972 11772
rect 7024 11354 7052 15302
rect 7116 14482 7144 19110
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 7116 13462 7144 13942
rect 7104 13456 7156 13462
rect 7104 13398 7156 13404
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 7116 11558 7144 12378
rect 7208 12170 7236 19178
rect 7392 19174 7420 20266
rect 7484 20058 7512 20295
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 7380 19168 7432 19174
rect 7380 19110 7432 19116
rect 7576 18970 7604 20402
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 8036 20346 8064 22200
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 7656 19848 7708 19854
rect 7656 19790 7708 19796
rect 7564 18964 7616 18970
rect 7564 18906 7616 18912
rect 7668 18698 7696 19790
rect 7656 18692 7708 18698
rect 7656 18634 7708 18640
rect 7656 18284 7708 18290
rect 7656 18226 7708 18232
rect 7668 18086 7696 18226
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7288 17740 7340 17746
rect 7288 17682 7340 17688
rect 7300 15042 7328 17682
rect 7472 17604 7524 17610
rect 7472 17546 7524 17552
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7392 17338 7420 17478
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7484 15162 7512 17546
rect 7564 16652 7616 16658
rect 7564 16594 7616 16600
rect 7576 15162 7604 16594
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7300 15014 7420 15042
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 7300 14074 7328 14894
rect 7392 14822 7420 15014
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7392 12782 7420 13330
rect 7288 12776 7340 12782
rect 7380 12776 7432 12782
rect 7288 12718 7340 12724
rect 7378 12744 7380 12753
rect 7432 12744 7434 12753
rect 7196 12164 7248 12170
rect 7196 12106 7248 12112
rect 7300 11898 7328 12718
rect 7378 12679 7434 12688
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7300 11694 7328 11834
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 7300 11354 7328 11630
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7194 11248 7250 11257
rect 6920 11212 6972 11218
rect 7300 11218 7328 11290
rect 7194 11183 7250 11192
rect 7288 11212 7340 11218
rect 6920 11154 6972 11160
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6840 10266 6868 10542
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6932 10198 6960 11154
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7010 10296 7066 10305
rect 7010 10231 7066 10240
rect 6920 10192 6972 10198
rect 6920 10134 6972 10140
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6552 9172 6604 9178
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 5920 8430 5948 8978
rect 6012 8634 6040 9166
rect 6840 9160 6868 10066
rect 6932 9654 6960 10134
rect 7024 10130 7052 10231
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 7024 9450 7052 10066
rect 7012 9444 7064 9450
rect 7012 9386 7064 9392
rect 6840 9132 6960 9160
rect 6552 9114 6604 9120
rect 6826 9072 6882 9081
rect 6826 9007 6828 9016
rect 6880 9007 6882 9016
rect 6828 8978 6880 8984
rect 6932 8922 6960 9132
rect 6840 8894 6960 8922
rect 7012 8900 7064 8906
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6564 8634 6592 8774
rect 6000 8628 6052 8634
rect 6552 8628 6604 8634
rect 6052 8588 6132 8616
rect 6000 8570 6052 8576
rect 6104 8498 6132 8588
rect 6552 8570 6604 8576
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5632 7482 5684 7488
rect 5736 7500 5856 7528
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5460 5817 5488 7142
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5446 5808 5502 5817
rect 5356 5772 5408 5778
rect 5446 5743 5502 5752
rect 5356 5714 5408 5720
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5368 5234 5396 5714
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5552 4826 5580 6598
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5368 4214 5396 4626
rect 5540 4548 5592 4554
rect 5540 4490 5592 4496
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 5262 4040 5318 4049
rect 5262 3975 5318 3984
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5092 3126 5120 3674
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 5276 2990 5304 3975
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 4988 2916 5040 2922
rect 4988 2858 5040 2864
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4304 2264 4384 2292
rect 4252 2246 4304 2252
rect 4540 800 4568 2382
rect 5000 800 5028 2858
rect 5368 2854 5396 3334
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5368 2514 5396 2586
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 5460 2446 5488 3334
rect 5552 2582 5580 4490
rect 5644 4026 5672 7346
rect 5736 6798 5764 7500
rect 5920 7449 5948 7686
rect 5906 7440 5962 7449
rect 5816 7404 5868 7410
rect 5906 7375 5962 7384
rect 5816 7346 5868 7352
rect 5828 7002 5856 7346
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5828 5681 5856 5714
rect 5814 5672 5870 5681
rect 5814 5607 5870 5616
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5736 5302 5764 5510
rect 5724 5296 5776 5302
rect 5724 5238 5776 5244
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5736 4214 5764 5102
rect 5828 4826 5856 5170
rect 5920 4826 5948 7278
rect 6012 7274 6040 8434
rect 6090 8392 6146 8401
rect 6090 8327 6146 8336
rect 6104 8022 6132 8327
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 6366 7984 6422 7993
rect 6366 7919 6422 7928
rect 6550 7984 6606 7993
rect 6550 7919 6606 7928
rect 6380 7818 6408 7919
rect 6564 7886 6592 7919
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 6656 7546 6684 8774
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6276 7336 6328 7342
rect 6276 7278 6328 7284
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6012 5250 6040 6734
rect 6288 6662 6316 7278
rect 6550 6896 6606 6905
rect 6550 6831 6606 6840
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6564 5953 6592 6831
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6656 6662 6684 6734
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6550 5944 6606 5953
rect 6550 5879 6606 5888
rect 6564 5778 6592 5879
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6748 5710 6776 8434
rect 6840 6905 6868 8894
rect 7012 8842 7064 8848
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 6932 8090 6960 8570
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6932 7342 6960 8026
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6826 6896 6882 6905
rect 6826 6831 6882 6840
rect 6828 6792 6880 6798
rect 6826 6760 6828 6769
rect 6880 6760 6882 6769
rect 6826 6695 6882 6704
rect 7024 6644 7052 8842
rect 7116 7721 7144 10610
rect 7208 10266 7236 11183
rect 7288 11154 7340 11160
rect 7288 10532 7340 10538
rect 7288 10474 7340 10480
rect 7300 10441 7328 10474
rect 7286 10432 7342 10441
rect 7286 10367 7342 10376
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7288 8900 7340 8906
rect 7392 8888 7420 12242
rect 7340 8860 7420 8888
rect 7288 8842 7340 8848
rect 7484 8650 7512 14418
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7576 14006 7604 14214
rect 7564 14000 7616 14006
rect 7564 13942 7616 13948
rect 7668 13954 7696 18022
rect 7760 17814 7788 20334
rect 8036 20318 8156 20346
rect 8128 19854 8156 20318
rect 8024 19848 8076 19854
rect 8024 19790 8076 19796
rect 8116 19848 8168 19854
rect 8116 19790 8168 19796
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 7748 17808 7800 17814
rect 7748 17750 7800 17756
rect 7852 17270 7880 18022
rect 7944 17338 7972 18158
rect 8036 17338 8064 19790
rect 8128 19514 8156 19790
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 8312 19310 8340 20402
rect 8496 19786 8524 22200
rect 8956 20466 8984 22200
rect 9128 20596 9180 20602
rect 9128 20538 9180 20544
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 8574 19952 8630 19961
rect 8574 19887 8630 19896
rect 8484 19780 8536 19786
rect 8484 19722 8536 19728
rect 8392 19372 8444 19378
rect 8392 19314 8444 19320
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 8208 18692 8260 18698
rect 8208 18634 8260 18640
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 7840 17264 7892 17270
rect 7746 17232 7802 17241
rect 7840 17206 7892 17212
rect 8116 17264 8168 17270
rect 8116 17206 8168 17212
rect 7746 17167 7802 17176
rect 7760 17134 7788 17167
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 8128 16794 8156 17206
rect 8116 16788 8168 16794
rect 8116 16730 8168 16736
rect 8128 16658 8156 16730
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8220 16590 8248 18634
rect 8312 18465 8340 18702
rect 8298 18456 8354 18465
rect 8298 18391 8354 18400
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 8128 16182 8156 16390
rect 8220 16289 8248 16526
rect 8206 16280 8262 16289
rect 8206 16215 8262 16224
rect 8116 16176 8168 16182
rect 8116 16118 8168 16124
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7748 16040 7800 16046
rect 7746 16008 7748 16017
rect 7800 16008 7802 16017
rect 7746 15943 7802 15952
rect 7852 15706 7880 16050
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7944 15570 7972 15846
rect 7748 15564 7800 15570
rect 7748 15506 7800 15512
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 7760 15434 7788 15506
rect 7748 15428 7800 15434
rect 7748 15370 7800 15376
rect 8128 15201 8156 16118
rect 8312 15638 8340 18022
rect 8404 16658 8432 19314
rect 8496 18970 8524 19722
rect 8588 19174 8616 19887
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8576 18828 8628 18834
rect 8680 18816 8708 19790
rect 9140 19394 9168 20538
rect 9218 20496 9274 20505
rect 9416 20466 9444 22200
rect 9496 20596 9548 20602
rect 9496 20538 9548 20544
rect 9404 20460 9456 20466
rect 9218 20431 9274 20440
rect 9232 20058 9260 20431
rect 9324 20420 9404 20448
rect 9220 20052 9272 20058
rect 9220 19994 9272 20000
rect 9220 19780 9272 19786
rect 9220 19722 9272 19728
rect 9232 19417 9260 19722
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 9048 19366 9168 19394
rect 9218 19408 9274 19417
rect 8956 19174 8984 19314
rect 9048 19281 9076 19366
rect 9218 19343 9274 19352
rect 9034 19272 9090 19281
rect 9324 19242 9352 20420
rect 9404 20402 9456 20408
rect 9404 19848 9456 19854
rect 9404 19790 9456 19796
rect 9034 19207 9090 19216
rect 9312 19236 9364 19242
rect 9312 19178 9364 19184
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 9310 19136 9366 19145
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 9140 18970 9168 19110
rect 9310 19071 9366 19080
rect 9128 18964 9180 18970
rect 9128 18906 9180 18912
rect 9324 18902 9352 19071
rect 9312 18896 9364 18902
rect 9312 18838 9364 18844
rect 8628 18788 8708 18816
rect 8576 18770 8628 18776
rect 8482 18728 8538 18737
rect 8482 18663 8538 18672
rect 8496 18630 8524 18663
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8484 18148 8536 18154
rect 8484 18090 8536 18096
rect 8496 17338 8524 18090
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 8390 16280 8446 16289
rect 8390 16215 8392 16224
rect 8444 16215 8446 16224
rect 8392 16186 8444 16192
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8300 15632 8352 15638
rect 8300 15574 8352 15580
rect 8114 15192 8170 15201
rect 7932 15156 7984 15162
rect 8114 15127 8170 15136
rect 8298 15192 8354 15201
rect 8298 15127 8354 15136
rect 7932 15098 7984 15104
rect 7944 14890 7972 15098
rect 8114 15056 8170 15065
rect 8114 14991 8170 15000
rect 8208 15020 8260 15026
rect 8128 14958 8156 14991
rect 8208 14962 8260 14968
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 7932 14884 7984 14890
rect 7932 14826 7984 14832
rect 8024 14884 8076 14890
rect 8024 14826 8076 14832
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 7944 14346 7972 14418
rect 7932 14340 7984 14346
rect 7932 14282 7984 14288
rect 7840 14000 7892 14006
rect 7668 13926 7788 13954
rect 7840 13942 7892 13948
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7576 10266 7604 13126
rect 7668 13025 7696 13670
rect 7654 13016 7710 13025
rect 7654 12951 7710 12960
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7668 9450 7696 12854
rect 7656 9444 7708 9450
rect 7656 9386 7708 9392
rect 7760 9178 7788 13926
rect 7852 12442 7880 13942
rect 7932 13864 7984 13870
rect 7932 13806 7984 13812
rect 7944 13530 7972 13806
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 8036 12646 8064 14826
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8128 14482 8156 14758
rect 8116 14476 8168 14482
rect 8116 14418 8168 14424
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 7930 11928 7986 11937
rect 7930 11863 7986 11872
rect 7944 11830 7972 11863
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 7932 11688 7984 11694
rect 7932 11630 7984 11636
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7484 8622 7604 8650
rect 7472 8560 7524 8566
rect 7472 8502 7524 8508
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7196 7948 7248 7954
rect 7196 7890 7248 7896
rect 7102 7712 7158 7721
rect 7102 7647 7158 7656
rect 7116 7313 7144 7647
rect 7208 7410 7236 7890
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7300 7546 7328 7686
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7102 7304 7158 7313
rect 7102 7239 7158 7248
rect 7208 7002 7236 7346
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 6840 6616 7052 6644
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 6656 5370 6684 5510
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6012 5222 6132 5250
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 6012 4622 6040 5102
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 5908 4480 5960 4486
rect 6104 4468 6132 5222
rect 6552 5160 6604 5166
rect 6550 5128 6552 5137
rect 6840 5148 6868 6616
rect 7010 6080 7066 6089
rect 7010 6015 7066 6024
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6604 5128 6606 5137
rect 6550 5063 6606 5072
rect 6748 5120 6868 5148
rect 6748 4486 6776 5120
rect 6932 5098 6960 5646
rect 7024 5574 7052 6015
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7010 5400 7066 5409
rect 7010 5335 7066 5344
rect 6920 5092 6972 5098
rect 6920 5034 6972 5040
rect 7024 5030 7052 5335
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 7116 4826 7144 6802
rect 7392 6458 7420 8366
rect 7484 7546 7512 8502
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7472 6316 7524 6322
rect 7576 6304 7604 8622
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7524 6276 7604 6304
rect 7472 6258 7524 6264
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7208 5914 7236 6190
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7300 5778 7328 5850
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7012 4752 7064 4758
rect 7208 4706 7236 4966
rect 7064 4700 7236 4706
rect 7012 4694 7236 4700
rect 7024 4678 7236 4694
rect 6840 4554 6960 4570
rect 6840 4548 6972 4554
rect 6840 4542 6920 4548
rect 5908 4422 5960 4428
rect 6012 4440 6132 4468
rect 6736 4480 6788 4486
rect 5920 4282 5948 4422
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 5724 4208 5776 4214
rect 5724 4150 5776 4156
rect 5724 4072 5776 4078
rect 5644 4020 5724 4026
rect 5644 4014 5776 4020
rect 5644 3998 5764 4014
rect 6012 2774 6040 4440
rect 6736 4422 6788 4428
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 6840 4214 6868 4542
rect 6920 4490 6972 4496
rect 6828 4208 6880 4214
rect 6550 4176 6606 4185
rect 6828 4150 6880 4156
rect 7196 4208 7248 4214
rect 7196 4150 7248 4156
rect 6550 4111 6606 4120
rect 6564 4010 6592 4111
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6196 3641 6224 3878
rect 6182 3632 6238 3641
rect 6564 3602 6592 3946
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6182 3567 6238 3576
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6748 3534 6776 3878
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 6656 3194 6684 3334
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 5644 2746 6040 2774
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 5644 2514 5672 2746
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5460 800 5488 2382
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 5920 800 5948 2314
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 6564 1442 6592 2926
rect 6840 2774 6868 4150
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 7024 3738 7052 4014
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7024 3126 7052 3674
rect 7208 3466 7236 4150
rect 7196 3460 7248 3466
rect 7196 3402 7248 3408
rect 7288 3392 7340 3398
rect 7392 3369 7420 5510
rect 7288 3334 7340 3340
rect 7378 3360 7434 3369
rect 7012 3120 7064 3126
rect 7012 3062 7064 3068
rect 6656 2746 6868 2774
rect 6656 2106 6684 2746
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 6748 1970 6776 2246
rect 6736 1964 6788 1970
rect 6736 1906 6788 1912
rect 6380 1414 6592 1442
rect 6380 800 6408 1414
rect 6840 800 6868 2382
rect 7300 800 7328 3334
rect 7378 3295 7434 3304
rect 7484 2990 7512 6258
rect 7562 6216 7618 6225
rect 7562 6151 7618 6160
rect 7576 3398 7604 6151
rect 7668 4690 7696 8230
rect 7760 8090 7788 8774
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7852 7970 7880 11494
rect 7944 10810 7972 11630
rect 7932 10804 7984 10810
rect 7932 10746 7984 10752
rect 7932 10600 7984 10606
rect 7930 10568 7932 10577
rect 7984 10568 7986 10577
rect 7930 10503 7986 10512
rect 7944 10266 7972 10503
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 8036 10062 8064 12378
rect 8128 12306 8156 14418
rect 8220 12442 8248 14962
rect 8312 14550 8340 15127
rect 8300 14544 8352 14550
rect 8300 14486 8352 14492
rect 8404 13938 8432 15846
rect 8496 14074 8524 17138
rect 8588 16114 8616 18770
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 8772 18170 8800 18702
rect 9220 18624 9272 18630
rect 8680 18142 8800 18170
rect 9140 18584 9220 18612
rect 9140 18154 9168 18584
rect 9416 18601 9444 19790
rect 9508 19242 9536 20538
rect 9876 19922 9904 22200
rect 10336 20466 10364 22200
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10140 20392 10192 20398
rect 10140 20334 10192 20340
rect 9956 20324 10008 20330
rect 9956 20266 10008 20272
rect 9864 19916 9916 19922
rect 9864 19858 9916 19864
rect 9770 19816 9826 19825
rect 9770 19751 9826 19760
rect 9586 19680 9642 19689
rect 9586 19615 9642 19624
rect 9600 19514 9628 19615
rect 9784 19514 9812 19751
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9680 19440 9732 19446
rect 9680 19382 9732 19388
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9496 19236 9548 19242
rect 9496 19178 9548 19184
rect 9600 19122 9628 19314
rect 9508 19094 9628 19122
rect 9508 18630 9536 19094
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 9496 18624 9548 18630
rect 9220 18566 9272 18572
rect 9402 18592 9458 18601
rect 9496 18566 9548 18572
rect 9402 18527 9458 18536
rect 9600 18306 9628 18906
rect 9692 18426 9720 19382
rect 9864 19236 9916 19242
rect 9864 19178 9916 19184
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 9784 18873 9812 19110
rect 9770 18864 9826 18873
rect 9770 18799 9826 18808
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9600 18278 9720 18306
rect 9220 18268 9272 18274
rect 9220 18210 9272 18216
rect 9128 18148 9180 18154
rect 8680 16538 8708 18142
rect 9232 18136 9260 18210
rect 9496 18148 9548 18154
rect 9232 18108 9352 18136
rect 9128 18090 9180 18096
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 9324 17864 9352 18108
rect 9496 18090 9548 18096
rect 9404 18080 9456 18086
rect 9402 18048 9404 18057
rect 9456 18048 9458 18057
rect 9402 17983 9458 17992
rect 9508 17882 9536 18090
rect 9586 18048 9642 18057
rect 9586 17983 9642 17992
rect 9232 17836 9352 17864
rect 9496 17876 9548 17882
rect 9128 17536 9180 17542
rect 9128 17478 9180 17484
rect 9140 17338 9168 17478
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 9232 16674 9260 17836
rect 9496 17818 9548 17824
rect 9404 17672 9456 17678
rect 9600 17649 9628 17983
rect 9692 17882 9720 18278
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9678 17776 9734 17785
rect 9678 17711 9680 17720
rect 9732 17711 9734 17720
rect 9680 17682 9732 17688
rect 9404 17614 9456 17620
rect 9586 17640 9642 17649
rect 9416 17134 9444 17614
rect 9586 17575 9642 17584
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9232 16646 9536 16674
rect 9692 16658 9720 16934
rect 9220 16584 9272 16590
rect 8680 16510 8800 16538
rect 9220 16526 9272 16532
rect 8668 16448 8720 16454
rect 8668 16390 8720 16396
rect 8576 16108 8628 16114
rect 8576 16050 8628 16056
rect 8576 15972 8628 15978
rect 8576 15914 8628 15920
rect 8588 15162 8616 15914
rect 8680 15366 8708 16390
rect 8772 16250 8800 16510
rect 9128 16516 9180 16522
rect 9128 16458 9180 16464
rect 8760 16244 8812 16250
rect 8760 16186 8812 16192
rect 9140 16182 9168 16458
rect 9128 16176 9180 16182
rect 9128 16118 9180 16124
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 9034 15192 9090 15201
rect 8576 15156 8628 15162
rect 9034 15127 9036 15136
rect 8576 15098 8628 15104
rect 9088 15127 9090 15136
rect 9036 15098 9088 15104
rect 9128 14952 9180 14958
rect 9128 14894 9180 14900
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 9140 14618 9168 14894
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 8760 14544 8812 14550
rect 8758 14512 8760 14521
rect 8812 14512 8814 14521
rect 8758 14447 8814 14456
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8864 14006 8892 14350
rect 8852 14000 8904 14006
rect 8852 13942 8904 13948
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 9232 13530 9260 16526
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9324 16250 9352 16390
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9416 16114 9444 16390
rect 9404 16108 9456 16114
rect 9404 16050 9456 16056
rect 9402 16008 9458 16017
rect 9324 15966 9402 15994
rect 9324 15502 9352 15966
rect 9402 15943 9458 15952
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9416 15609 9444 15846
rect 9402 15600 9458 15609
rect 9402 15535 9458 15544
rect 9312 15496 9364 15502
rect 9404 15496 9456 15502
rect 9312 15438 9364 15444
rect 9402 15464 9404 15473
rect 9456 15464 9458 15473
rect 9402 15399 9458 15408
rect 9508 15162 9536 16646
rect 9680 16652 9732 16658
rect 9680 16594 9732 16600
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9310 14920 9366 14929
rect 9310 14855 9366 14864
rect 9324 14482 9352 14855
rect 9404 14816 9456 14822
rect 9404 14758 9456 14764
rect 9416 14482 9444 14758
rect 9312 14476 9364 14482
rect 9312 14418 9364 14424
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 8760 13456 8812 13462
rect 8666 13424 8722 13433
rect 8760 13398 8812 13404
rect 8666 13359 8668 13368
rect 8720 13359 8722 13368
rect 8668 13330 8720 13336
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8404 12986 8432 13126
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8772 12850 8800 13398
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 8404 12594 8432 12786
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8312 12566 8432 12594
rect 8208 12436 8260 12442
rect 8312 12434 8340 12566
rect 8588 12442 8616 12718
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8680 12442 8708 12582
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 8576 12436 8628 12442
rect 8312 12406 8432 12434
rect 8208 12378 8260 12384
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8116 11824 8168 11830
rect 8116 11766 8168 11772
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 7932 8900 7984 8906
rect 7932 8842 7984 8848
rect 7944 8430 7972 8842
rect 8036 8634 8064 9114
rect 8128 9110 8156 11766
rect 8116 9104 8168 9110
rect 8116 9046 8168 9052
rect 8220 9042 8248 12242
rect 8298 10160 8354 10169
rect 8298 10095 8354 10104
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7760 7942 7880 7970
rect 7760 6089 7788 7942
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7746 6080 7802 6089
rect 7746 6015 7802 6024
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 7668 3602 7696 4082
rect 7760 3777 7788 6015
rect 7852 5098 7880 7346
rect 7944 6866 7972 8366
rect 8220 8362 8248 8774
rect 8312 8430 8340 10095
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8036 7818 8064 8026
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 8128 7342 8156 8230
rect 8404 7970 8432 12406
rect 8576 12378 8628 12384
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 9324 12374 9352 12786
rect 9312 12368 9364 12374
rect 9312 12310 9364 12316
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8588 10062 8616 10678
rect 8680 10266 8708 11698
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 8772 10810 8800 10950
rect 8760 10804 8812 10810
rect 8760 10746 8812 10752
rect 9036 10804 9088 10810
rect 9140 10792 9168 12038
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 9088 10764 9168 10792
rect 9036 10746 9088 10752
rect 9126 10568 9182 10577
rect 9126 10503 9182 10512
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8484 9920 8536 9926
rect 8482 9888 8484 9897
rect 8536 9888 8538 9897
rect 8482 9823 8538 9832
rect 8484 9376 8536 9382
rect 8482 9344 8484 9353
rect 8536 9344 8538 9353
rect 8482 9279 8538 9288
rect 8588 9042 8616 9998
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 8666 9616 8722 9625
rect 8666 9551 8722 9560
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8220 7954 8432 7970
rect 8496 7954 8524 8978
rect 8680 8945 8708 9551
rect 9048 9382 9076 9862
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 8760 9036 8812 9042
rect 8760 8978 8812 8984
rect 8666 8936 8722 8945
rect 8666 8871 8722 8880
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8588 8634 8616 8774
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8680 8514 8708 8871
rect 8772 8838 8800 8978
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8588 8486 8708 8514
rect 8208 7948 8432 7954
rect 8260 7942 8432 7948
rect 8484 7948 8536 7954
rect 8208 7890 8260 7896
rect 8484 7890 8536 7896
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7932 6656 7984 6662
rect 7930 6624 7932 6633
rect 7984 6624 7986 6633
rect 7930 6559 7986 6568
rect 7944 6100 7972 6559
rect 8024 6248 8076 6254
rect 8128 6236 8156 7278
rect 8220 6934 8248 7414
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 8076 6208 8156 6236
rect 8024 6190 8076 6196
rect 8116 6112 8168 6118
rect 7944 6072 8064 6100
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7944 5370 7972 5510
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 7930 5264 7986 5273
rect 7930 5199 7986 5208
rect 7840 5092 7892 5098
rect 7840 5034 7892 5040
rect 7944 4758 7972 5199
rect 7932 4752 7984 4758
rect 7932 4694 7984 4700
rect 7944 3942 7972 4694
rect 8036 4593 8064 6072
rect 8116 6054 8168 6060
rect 8128 5778 8156 6054
rect 8220 5930 8248 6870
rect 8312 6458 8340 7346
rect 8404 7002 8432 7686
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8298 6352 8354 6361
rect 8298 6287 8300 6296
rect 8352 6287 8354 6296
rect 8300 6258 8352 6264
rect 8404 6089 8432 6598
rect 8588 6361 8616 8486
rect 8668 8424 8720 8430
rect 8772 8412 8800 8774
rect 9140 8430 9168 10503
rect 8720 8384 8800 8412
rect 9128 8424 9180 8430
rect 8668 8366 8720 8372
rect 9128 8366 9180 8372
rect 8680 7886 8708 8366
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 9140 8090 9168 8366
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 9140 7886 9168 8026
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8574 6352 8630 6361
rect 8574 6287 8630 6296
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8390 6080 8446 6089
rect 8390 6015 8446 6024
rect 8220 5902 8432 5930
rect 8496 5914 8524 6190
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8298 5672 8354 5681
rect 8298 5607 8354 5616
rect 8022 4584 8078 4593
rect 8022 4519 8078 4528
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8036 4078 8064 4422
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 8114 4040 8170 4049
rect 8114 3975 8170 3984
rect 8128 3942 8156 3975
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 7746 3768 7802 3777
rect 7746 3703 7802 3712
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7668 3097 7696 3130
rect 7654 3088 7710 3097
rect 7654 3023 7710 3032
rect 7472 2984 7524 2990
rect 7472 2926 7524 2932
rect 7760 2446 7788 3334
rect 8220 3194 8248 4422
rect 8312 4321 8340 5607
rect 8298 4312 8354 4321
rect 8404 4282 8432 5902
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8496 5166 8524 5850
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8496 4706 8524 4966
rect 8588 4826 8616 5850
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8496 4678 8616 4706
rect 8298 4247 8354 4256
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8484 4208 8536 4214
rect 8484 4150 8536 4156
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8312 3126 8340 3334
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7760 800 7788 2382
rect 8404 2378 8432 3402
rect 8496 3194 8524 4150
rect 8588 3233 8616 4678
rect 8680 3618 8708 7346
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 9126 6896 9182 6905
rect 9232 6866 9260 11698
rect 9324 11626 9352 12174
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9416 11257 9444 13262
rect 9508 11762 9536 13874
rect 9600 12986 9628 16526
rect 9692 15366 9720 16594
rect 9784 16250 9812 18702
rect 9876 18154 9904 19178
rect 9968 18714 9996 20266
rect 10048 19780 10100 19786
rect 10048 19722 10100 19728
rect 10060 19514 10088 19722
rect 10152 19553 10180 20334
rect 10232 19848 10284 19854
rect 10232 19790 10284 19796
rect 10138 19544 10194 19553
rect 10048 19508 10100 19514
rect 10138 19479 10194 19488
rect 10048 19450 10100 19456
rect 10244 19417 10272 19790
rect 10230 19408 10286 19417
rect 10140 19372 10192 19378
rect 10230 19343 10286 19352
rect 10140 19314 10192 19320
rect 10152 19258 10180 19314
rect 10152 19230 10272 19258
rect 10048 18896 10100 18902
rect 10100 18844 10180 18850
rect 10048 18838 10180 18844
rect 10060 18822 10180 18838
rect 9968 18686 10088 18714
rect 9956 18624 10008 18630
rect 9954 18592 9956 18601
rect 10008 18592 10010 18601
rect 9954 18527 10010 18536
rect 9864 18148 9916 18154
rect 9864 18090 9916 18096
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9876 16402 9904 17750
rect 9956 17536 10008 17542
rect 9956 17478 10008 17484
rect 9968 17202 9996 17478
rect 10060 17338 10088 18686
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9968 16969 9996 17138
rect 9954 16960 10010 16969
rect 9954 16895 10010 16904
rect 10046 16552 10102 16561
rect 10046 16487 10048 16496
rect 10100 16487 10102 16496
rect 10048 16458 10100 16464
rect 9876 16374 10088 16402
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9784 15706 9812 15846
rect 9772 15700 9824 15706
rect 9772 15642 9824 15648
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9692 14890 9720 15302
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9692 12714 9720 13874
rect 9680 12708 9732 12714
rect 9680 12650 9732 12656
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9600 12209 9628 12242
rect 9586 12200 9642 12209
rect 9586 12135 9642 12144
rect 9784 11914 9812 14962
rect 9876 14618 9904 16050
rect 9956 16040 10008 16046
rect 9954 16008 9956 16017
rect 10008 16008 10010 16017
rect 9954 15943 10010 15952
rect 9968 15473 9996 15943
rect 9954 15464 10010 15473
rect 9954 15399 10010 15408
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9876 13938 9904 14214
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 9864 13184 9916 13190
rect 9862 13152 9864 13161
rect 9916 13152 9918 13161
rect 9862 13087 9918 13096
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 9692 11898 9812 11914
rect 9680 11892 9812 11898
rect 9732 11886 9812 11892
rect 9680 11834 9732 11840
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9402 11248 9458 11257
rect 9402 11183 9458 11192
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9324 9450 9352 11018
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9416 10810 9444 10950
rect 9494 10840 9550 10849
rect 9404 10804 9456 10810
rect 9692 10810 9720 11698
rect 9770 10840 9826 10849
rect 9494 10775 9496 10784
rect 9404 10746 9456 10752
rect 9548 10775 9550 10784
rect 9680 10804 9732 10810
rect 9496 10746 9548 10752
rect 9770 10775 9826 10784
rect 9680 10746 9732 10752
rect 9508 10690 9536 10746
rect 9508 10662 9720 10690
rect 9784 10674 9812 10775
rect 9496 10600 9548 10606
rect 9494 10568 9496 10577
rect 9548 10568 9550 10577
rect 9494 10503 9550 10512
rect 9402 10024 9458 10033
rect 9402 9959 9458 9968
rect 9416 9926 9444 9959
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9402 9616 9458 9625
rect 9508 9586 9536 10503
rect 9402 9551 9458 9560
rect 9496 9580 9548 9586
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 9324 7002 9352 7754
rect 9416 7342 9444 9551
rect 9496 9522 9548 9528
rect 9586 9480 9642 9489
rect 9586 9415 9642 9424
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9126 6831 9182 6840
rect 9220 6860 9272 6866
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9048 6458 9076 6598
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9140 6322 9168 6831
rect 9220 6802 9272 6808
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8772 5030 8800 5510
rect 8864 5409 8892 5714
rect 9036 5568 9088 5574
rect 9140 5556 9168 6258
rect 9088 5528 9168 5556
rect 9036 5510 9088 5516
rect 8850 5400 8906 5409
rect 8850 5335 8906 5344
rect 9128 5092 9180 5098
rect 9128 5034 9180 5040
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 9034 4312 9090 4321
rect 9140 4282 9168 5034
rect 9034 4247 9090 4256
rect 9128 4276 9180 4282
rect 9048 4078 9076 4247
rect 9128 4218 9180 4224
rect 9036 4072 9088 4078
rect 9036 4014 9088 4020
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 9126 3768 9182 3777
rect 9126 3703 9182 3712
rect 8680 3590 8800 3618
rect 9140 3602 9168 3703
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8574 3224 8630 3233
rect 8484 3188 8536 3194
rect 8574 3159 8630 3168
rect 8484 3130 8536 3136
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8588 2650 8616 2994
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8208 2372 8260 2378
rect 8208 2314 8260 2320
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8220 800 8248 2314
rect 8680 800 8708 3470
rect 8772 2922 8800 3590
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 9128 3596 9180 3602
rect 9128 3538 9180 3544
rect 8956 3194 8984 3538
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9128 3120 9180 3126
rect 9128 3062 9180 3068
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 9140 800 9168 3062
rect 9232 2514 9260 6802
rect 9310 6624 9366 6633
rect 9310 6559 9366 6568
rect 9324 6254 9352 6559
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9310 5400 9366 5409
rect 9310 5335 9312 5344
rect 9364 5335 9366 5344
rect 9312 5306 9364 5312
rect 9508 5273 9536 9318
rect 9600 9178 9628 9415
rect 9692 9364 9720 10662
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9876 10554 9904 12786
rect 9968 12442 9996 13194
rect 9956 12436 10008 12442
rect 10060 12434 10088 16374
rect 10152 14006 10180 18822
rect 10244 18193 10272 19230
rect 10336 18426 10364 20402
rect 10416 19440 10468 19446
rect 10416 19382 10468 19388
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10230 18184 10286 18193
rect 10230 18119 10286 18128
rect 10244 18086 10272 18119
rect 10428 18086 10456 19382
rect 10520 18601 10548 20946
rect 10692 19916 10744 19922
rect 10692 19858 10744 19864
rect 10600 19712 10652 19718
rect 10600 19654 10652 19660
rect 10506 18592 10562 18601
rect 10506 18527 10562 18536
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10416 18080 10468 18086
rect 10416 18022 10468 18028
rect 10232 17876 10284 17882
rect 10232 17818 10284 17824
rect 10416 17876 10468 17882
rect 10416 17818 10468 17824
rect 10244 16590 10272 17818
rect 10428 16658 10456 17818
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 10244 12646 10272 16526
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10336 14414 10364 16390
rect 10428 15706 10456 16594
rect 10506 16552 10562 16561
rect 10506 16487 10562 16496
rect 10520 16046 10548 16487
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10612 15638 10640 19654
rect 10704 18290 10732 19858
rect 10796 19310 10824 22200
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 10796 18358 10824 19246
rect 10876 19168 10928 19174
rect 10968 19168 11020 19174
rect 10876 19110 10928 19116
rect 10966 19136 10968 19145
rect 11020 19136 11022 19145
rect 10784 18352 10836 18358
rect 10784 18294 10836 18300
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10704 16017 10732 18022
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10796 16182 10824 16390
rect 10888 16250 10916 19110
rect 10966 19071 11022 19080
rect 11072 18698 11100 20198
rect 11256 19922 11284 22200
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 11716 20466 11744 22200
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11808 20058 11836 20878
rect 11888 20868 11940 20874
rect 11888 20810 11940 20816
rect 11900 20330 11928 20810
rect 12176 20806 12204 22200
rect 12636 22114 12664 22200
rect 12728 22114 12756 22222
rect 12636 22086 12756 22114
rect 12808 20868 12860 20874
rect 12808 20810 12860 20816
rect 12164 20800 12216 20806
rect 12164 20742 12216 20748
rect 12622 20632 12678 20641
rect 12622 20567 12678 20576
rect 12636 20534 12664 20567
rect 12820 20534 12848 20810
rect 12624 20528 12676 20534
rect 12624 20470 12676 20476
rect 12808 20528 12860 20534
rect 12808 20470 12860 20476
rect 12072 20460 12124 20466
rect 12072 20402 12124 20408
rect 11888 20324 11940 20330
rect 11888 20266 11940 20272
rect 11796 20052 11848 20058
rect 11796 19994 11848 20000
rect 11888 20052 11940 20058
rect 11888 19994 11940 20000
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11152 19848 11204 19854
rect 11152 19790 11204 19796
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 11072 16538 11100 18634
rect 10980 16510 11100 16538
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 10784 16176 10836 16182
rect 10784 16118 10836 16124
rect 10690 16008 10746 16017
rect 10690 15943 10746 15952
rect 10600 15632 10652 15638
rect 10600 15574 10652 15580
rect 10980 15434 11008 16510
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11072 16250 11100 16390
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11164 16130 11192 19790
rect 11256 19514 11284 19858
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11244 19236 11296 19242
rect 11244 19178 11296 19184
rect 11256 18630 11284 19178
rect 11244 18624 11296 18630
rect 11244 18566 11296 18572
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11716 18290 11744 19314
rect 11808 18714 11836 19654
rect 11900 19378 11928 19994
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11808 18698 11928 18714
rect 11808 18692 11940 18698
rect 11808 18686 11888 18692
rect 11808 18329 11836 18686
rect 11888 18634 11940 18640
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11794 18320 11850 18329
rect 11704 18284 11756 18290
rect 11794 18255 11850 18264
rect 11704 18226 11756 18232
rect 11520 18080 11572 18086
rect 11518 18048 11520 18057
rect 11572 18048 11574 18057
rect 11518 17983 11574 17992
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11624 16658 11652 16934
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 11072 16102 11192 16130
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10704 15162 10732 15302
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10416 15020 10468 15026
rect 10416 14962 10468 14968
rect 10428 14822 10456 14962
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10060 12406 10272 12434
rect 9956 12378 10008 12384
rect 9954 12336 10010 12345
rect 9954 12271 10010 12280
rect 9968 11694 9996 12271
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9954 11384 10010 11393
rect 9954 11319 10010 11328
rect 9968 11218 9996 11319
rect 10060 11286 10088 12038
rect 10048 11280 10100 11286
rect 10048 11222 10100 11228
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9784 10526 9904 10554
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9784 10470 9812 10526
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9784 9654 9812 9862
rect 9772 9648 9824 9654
rect 9772 9590 9824 9596
rect 9772 9512 9824 9518
rect 9770 9480 9772 9489
rect 9824 9480 9826 9489
rect 9770 9415 9826 9424
rect 9772 9376 9824 9382
rect 9692 9344 9772 9364
rect 9824 9344 9826 9353
rect 9692 9336 9770 9344
rect 9770 9279 9826 9288
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9678 8936 9734 8945
rect 9784 8906 9812 9114
rect 9678 8871 9734 8880
rect 9772 8900 9824 8906
rect 9692 8566 9720 8871
rect 9772 8842 9824 8848
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9784 8498 9812 8842
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9784 7970 9812 8434
rect 9876 8430 9904 10406
rect 9968 10062 9996 10542
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 10060 8922 10088 9930
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10152 9042 10180 9318
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 9968 8634 9996 8910
rect 10060 8894 10180 8922
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 10060 8634 10088 8774
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10152 8566 10180 8894
rect 10140 8560 10192 8566
rect 10140 8502 10192 8508
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 10060 8362 10088 8434
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 9692 7942 9812 7970
rect 10048 7948 10100 7954
rect 9692 6934 9720 7942
rect 10048 7890 10100 7896
rect 9770 7848 9826 7857
rect 9770 7783 9826 7792
rect 9784 7750 9812 7783
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9864 7200 9916 7206
rect 9864 7142 9916 7148
rect 9954 7168 10010 7177
rect 9680 6928 9732 6934
rect 9586 6896 9642 6905
rect 9680 6870 9732 6876
rect 9586 6831 9642 6840
rect 9600 6662 9628 6831
rect 9680 6792 9732 6798
rect 9678 6760 9680 6769
rect 9732 6760 9734 6769
rect 9678 6695 9734 6704
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9772 5636 9824 5642
rect 9772 5578 9824 5584
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9494 5264 9550 5273
rect 9404 5228 9456 5234
rect 9494 5199 9550 5208
rect 9404 5170 9456 5176
rect 9310 4992 9366 5001
rect 9310 4927 9366 4936
rect 9324 4826 9352 4927
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9312 4480 9364 4486
rect 9416 4468 9444 5170
rect 9496 5160 9548 5166
rect 9496 5102 9548 5108
rect 9508 5030 9536 5102
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9364 4440 9444 4468
rect 9312 4422 9364 4428
rect 9416 4282 9444 4440
rect 9496 4480 9548 4486
rect 9496 4422 9548 4428
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9508 4214 9536 4422
rect 9312 4208 9364 4214
rect 9312 4150 9364 4156
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9324 4026 9352 4150
rect 9324 3998 9444 4026
rect 9310 3632 9366 3641
rect 9310 3567 9366 3576
rect 9324 3534 9352 3567
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 9416 3194 9444 3998
rect 9508 3890 9536 4150
rect 9600 4010 9628 5510
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9692 4729 9720 5306
rect 9784 4826 9812 5578
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9678 4720 9734 4729
rect 9678 4655 9734 4664
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9692 4282 9720 4422
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9588 4004 9640 4010
rect 9588 3946 9640 3952
rect 9508 3862 9628 3890
rect 9494 3632 9550 3641
rect 9600 3602 9628 3862
rect 9494 3567 9550 3576
rect 9588 3596 9640 3602
rect 9508 3466 9536 3567
rect 9588 3538 9640 3544
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9416 2990 9444 3130
rect 9600 3126 9628 3538
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9692 2854 9720 3334
rect 9784 3058 9812 4558
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 9218 2408 9274 2417
rect 9218 2343 9274 2352
rect 9232 2310 9260 2343
rect 9508 2310 9536 2586
rect 9692 2514 9720 2790
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9876 2446 9904 7142
rect 9954 7103 10010 7112
rect 9968 7002 9996 7103
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 9956 6724 10008 6730
rect 9956 6666 10008 6672
rect 9968 6458 9996 6666
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9956 5092 10008 5098
rect 9956 5034 10008 5040
rect 9968 4690 9996 5034
rect 10060 4758 10088 7890
rect 10152 6118 10180 8502
rect 10244 7834 10272 12406
rect 10336 11898 10364 14010
rect 10428 13841 10456 14758
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 10520 13977 10548 14418
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 10692 14000 10744 14006
rect 10506 13968 10562 13977
rect 10692 13942 10744 13948
rect 10506 13903 10562 13912
rect 10704 13870 10732 13942
rect 10692 13864 10744 13870
rect 10414 13832 10470 13841
rect 10692 13806 10744 13812
rect 10414 13767 10470 13776
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10428 12986 10456 13126
rect 10506 13016 10562 13025
rect 10416 12980 10468 12986
rect 10506 12951 10562 12960
rect 10416 12922 10468 12928
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10336 11286 10364 11834
rect 10324 11280 10376 11286
rect 10428 11257 10456 12106
rect 10324 11222 10376 11228
rect 10414 11248 10470 11257
rect 10414 11183 10470 11192
rect 10428 11150 10456 11183
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10414 10840 10470 10849
rect 10414 10775 10470 10784
rect 10428 9722 10456 10775
rect 10520 9926 10548 12951
rect 10612 12918 10640 13670
rect 10600 12912 10652 12918
rect 10600 12854 10652 12860
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10612 12102 10640 12582
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10612 10742 10640 11154
rect 10600 10736 10652 10742
rect 10600 10678 10652 10684
rect 10704 10010 10732 13806
rect 10784 13796 10836 13802
rect 10784 13738 10836 13744
rect 10796 12442 10824 13738
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10888 13326 10916 13670
rect 10980 13394 11008 14282
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10876 13184 10928 13190
rect 10874 13152 10876 13161
rect 10928 13152 10930 13161
rect 10874 13087 10930 13096
rect 10980 13025 11008 13330
rect 10966 13016 11022 13025
rect 10876 12980 10928 12986
rect 10966 12951 11022 12960
rect 10876 12922 10928 12928
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10784 12164 10836 12170
rect 10784 12106 10836 12112
rect 10796 11830 10824 12106
rect 10784 11824 10836 11830
rect 10784 11766 10836 11772
rect 10784 11688 10836 11694
rect 10782 11656 10784 11665
rect 10836 11656 10838 11665
rect 10782 11591 10838 11600
rect 10796 10588 10824 11591
rect 10888 11218 10916 12922
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 10980 12306 11008 12650
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 11072 12238 11100 16102
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11164 15502 11192 15982
rect 11256 15570 11284 16186
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11348 15348 11376 15642
rect 11164 15320 11376 15348
rect 11164 14482 11192 15320
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11716 15026 11744 17478
rect 11796 17060 11848 17066
rect 11796 17002 11848 17008
rect 11808 15706 11836 17002
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11796 15700 11848 15706
rect 11796 15642 11848 15648
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11256 14618 11284 14894
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11242 14512 11298 14521
rect 11152 14476 11204 14482
rect 11242 14447 11298 14456
rect 11152 14418 11204 14424
rect 11256 14074 11284 14447
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11244 14068 11296 14074
rect 11244 14010 11296 14016
rect 11900 13530 11928 16526
rect 11992 15065 12020 18566
rect 11978 15056 12034 15065
rect 11978 14991 12034 15000
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11612 13320 11664 13326
rect 11664 13280 11744 13308
rect 11612 13262 11664 13268
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11152 12368 11204 12374
rect 11152 12310 11204 12316
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10980 11694 11008 12038
rect 11072 11778 11100 12174
rect 11164 12102 11192 12310
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11256 11898 11284 13126
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11716 12889 11744 13280
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11702 12880 11758 12889
rect 11702 12815 11758 12824
rect 11808 12714 11836 13194
rect 11796 12708 11848 12714
rect 11796 12650 11848 12656
rect 11704 12164 11756 12170
rect 11704 12106 11756 12112
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11426 11792 11482 11801
rect 11072 11750 11192 11778
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 10876 10600 10928 10606
rect 10796 10560 10876 10588
rect 10876 10542 10928 10548
rect 10980 10418 11008 10678
rect 11072 10538 11100 11562
rect 11164 11558 11192 11750
rect 11716 11762 11744 12106
rect 11992 12050 12020 13330
rect 12084 12170 12112 20402
rect 12900 20392 12952 20398
rect 12900 20334 12952 20340
rect 12912 20058 12940 20334
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 12912 19854 12940 19994
rect 13004 19922 13032 22222
rect 13082 22200 13138 23000
rect 13542 22200 13598 23000
rect 14002 22200 14058 23000
rect 14462 22200 14518 23000
rect 14922 22200 14978 23000
rect 15382 22200 15438 23000
rect 15842 22200 15898 23000
rect 16302 22200 16358 23000
rect 16762 22200 16818 23000
rect 17222 22200 17278 23000
rect 17682 22200 17738 23000
rect 18142 22200 18198 23000
rect 18602 22200 18658 23000
rect 19062 22200 19118 23000
rect 19522 22200 19578 23000
rect 19982 22200 20038 23000
rect 20442 22200 20498 23000
rect 20902 22200 20958 23000
rect 21362 22200 21418 23000
rect 21822 22200 21878 23000
rect 22282 22200 22338 23000
rect 22742 22200 22798 23000
rect 13096 20058 13124 22200
rect 13556 20482 13584 22200
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13556 20454 13676 20482
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13648 20346 13676 20454
rect 13924 20398 13952 20742
rect 13912 20392 13964 20398
rect 13464 20074 13492 20334
rect 13648 20318 13860 20346
rect 13912 20334 13964 20340
rect 14016 20330 14044 22200
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 14108 20466 14136 20878
rect 14278 20632 14334 20641
rect 14476 20618 14504 22200
rect 14476 20602 14596 20618
rect 14476 20596 14608 20602
rect 14476 20590 14556 20596
rect 14278 20567 14334 20576
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 13832 20262 13860 20318
rect 14004 20324 14056 20330
rect 14004 20266 14056 20272
rect 13728 20256 13780 20262
rect 13728 20198 13780 20204
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13084 20052 13136 20058
rect 13084 19994 13136 20000
rect 13372 20046 13492 20074
rect 13740 20058 13768 20198
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 13728 20052 13780 20058
rect 12992 19916 13044 19922
rect 12992 19858 13044 19864
rect 12900 19848 12952 19854
rect 12900 19790 12952 19796
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 12624 19780 12676 19786
rect 12624 19722 12676 19728
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12452 19378 12480 19450
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12176 18057 12204 19314
rect 12532 18352 12584 18358
rect 12532 18294 12584 18300
rect 12162 18048 12218 18057
rect 12162 17983 12218 17992
rect 12346 17640 12402 17649
rect 12164 17604 12216 17610
rect 12346 17575 12402 17584
rect 12164 17546 12216 17552
rect 12176 15978 12204 17546
rect 12360 16794 12388 17575
rect 12440 17264 12492 17270
rect 12440 17206 12492 17212
rect 12452 16969 12480 17206
rect 12438 16960 12494 16969
rect 12438 16895 12494 16904
rect 12544 16794 12572 18294
rect 12636 17762 12664 19722
rect 12912 18766 12940 19790
rect 13188 19378 13216 19790
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 13268 19236 13320 19242
rect 13268 19178 13320 19184
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 12912 18290 12940 18702
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 12806 18048 12862 18057
rect 12806 17983 12862 17992
rect 12820 17882 12848 17983
rect 12912 17882 12940 18226
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 13004 17762 13032 18022
rect 12636 17734 13032 17762
rect 12728 17649 12756 17734
rect 12714 17640 12770 17649
rect 12714 17575 12770 17584
rect 12992 17604 13044 17610
rect 12992 17546 13044 17552
rect 13004 17490 13032 17546
rect 12820 17462 13032 17490
rect 12820 17338 12848 17462
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 13004 16794 13032 17138
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12532 16788 12584 16794
rect 12532 16730 12584 16736
rect 12992 16788 13044 16794
rect 12992 16730 13044 16736
rect 12900 16516 12952 16522
rect 12900 16458 12952 16464
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12164 15972 12216 15978
rect 12164 15914 12216 15920
rect 12176 14550 12204 15914
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12164 14544 12216 14550
rect 12164 14486 12216 14492
rect 12164 14272 12216 14278
rect 12164 14214 12216 14220
rect 12176 14006 12204 14214
rect 12164 14000 12216 14006
rect 12164 13942 12216 13948
rect 12176 12782 12204 13942
rect 12452 13841 12480 15846
rect 12544 13938 12572 16390
rect 12912 16114 12940 16458
rect 13096 16182 13124 18566
rect 13280 17921 13308 19178
rect 13266 17912 13322 17921
rect 13266 17847 13322 17856
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 13188 17338 13216 17682
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 13176 16992 13228 16998
rect 13174 16960 13176 16969
rect 13228 16960 13230 16969
rect 13174 16895 13230 16904
rect 13084 16176 13136 16182
rect 13084 16118 13136 16124
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12728 14822 12756 14962
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12532 13932 12584 13938
rect 12532 13874 12584 13880
rect 12438 13832 12494 13841
rect 12438 13767 12494 13776
rect 12452 13394 12480 13767
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 12544 12481 12572 13874
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12636 13326 12664 13670
rect 12820 13326 12848 15302
rect 13096 15094 13124 16118
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12912 13938 12940 14962
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12636 12646 12664 13262
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12530 12472 12586 12481
rect 12530 12407 12586 12416
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12532 12232 12584 12238
rect 12636 12220 12664 12582
rect 12584 12192 12664 12220
rect 12532 12174 12584 12180
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 11992 12022 12112 12050
rect 11978 11792 12034 11801
rect 11426 11727 11482 11736
rect 11704 11756 11756 11762
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11256 10742 11284 11086
rect 11440 11082 11468 11727
rect 11704 11698 11756 11704
rect 11888 11756 11940 11762
rect 11978 11727 12034 11736
rect 11888 11698 11940 11704
rect 11716 11642 11744 11698
rect 11624 11614 11744 11642
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11624 11393 11652 11614
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11610 11384 11666 11393
rect 11610 11319 11666 11328
rect 11520 11280 11572 11286
rect 11624 11268 11652 11319
rect 11572 11240 11652 11268
rect 11520 11222 11572 11228
rect 11610 11112 11666 11121
rect 11428 11076 11480 11082
rect 11610 11047 11612 11056
rect 11428 11018 11480 11024
rect 11664 11047 11666 11056
rect 11612 11018 11664 11024
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11716 10810 11744 11494
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 10612 9982 10732 10010
rect 10796 10390 11008 10418
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10322 9480 10378 9489
rect 10322 9415 10378 9424
rect 10336 9042 10364 9415
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10428 8480 10456 9658
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10520 9110 10548 9318
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 10508 8968 10560 8974
rect 10506 8936 10508 8945
rect 10560 8936 10562 8945
rect 10506 8871 10562 8880
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10336 8452 10456 8480
rect 10336 7954 10364 8452
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10324 7948 10376 7954
rect 10324 7890 10376 7896
rect 10244 7806 10364 7834
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 7002 10272 7686
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10336 6866 10364 7806
rect 10428 7313 10456 8298
rect 10520 7886 10548 8774
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10414 7304 10470 7313
rect 10414 7239 10470 7248
rect 10612 7206 10640 9982
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10600 7200 10652 7206
rect 10520 7160 10600 7188
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10322 5944 10378 5953
rect 10322 5879 10378 5888
rect 10336 5166 10364 5879
rect 10428 5778 10456 6938
rect 10520 6730 10548 7160
rect 10600 7142 10652 7148
rect 10508 6724 10560 6730
rect 10508 6666 10560 6672
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10612 6458 10640 6598
rect 10600 6452 10652 6458
rect 10600 6394 10652 6400
rect 10704 6254 10732 9862
rect 10796 9382 10824 10390
rect 11256 10062 11284 10678
rect 11244 10056 11296 10062
rect 11150 10024 11206 10033
rect 11244 9998 11296 10004
rect 11150 9959 11206 9968
rect 10968 9648 11020 9654
rect 10968 9590 11020 9596
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10796 8634 10824 8978
rect 10888 8945 10916 9454
rect 10874 8936 10930 8945
rect 10874 8871 10930 8880
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10796 6866 10824 8570
rect 10888 8362 10916 8871
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10980 8106 11008 9590
rect 11058 8528 11114 8537
rect 11058 8463 11114 8472
rect 10888 8078 11008 8106
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10888 6338 10916 8078
rect 11072 7970 11100 8463
rect 10980 7954 11100 7970
rect 10968 7948 11100 7954
rect 11020 7942 11100 7948
rect 10968 7890 11020 7896
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10980 6798 11008 7414
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10796 6310 10916 6338
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10414 5672 10470 5681
rect 10414 5607 10470 5616
rect 10324 5160 10376 5166
rect 10322 5128 10324 5137
rect 10376 5128 10378 5137
rect 10322 5063 10378 5072
rect 10048 4752 10100 4758
rect 10324 4752 10376 4758
rect 10048 4694 10100 4700
rect 10244 4712 10324 4740
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 9968 4162 9996 4626
rect 10060 4282 10088 4694
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 9968 4134 10180 4162
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 9968 3058 9996 4014
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10060 3602 10088 3878
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 9968 2774 9996 2994
rect 10060 2990 10088 3538
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 9968 2746 10088 2774
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9588 2372 9640 2378
rect 9588 2314 9640 2320
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 9232 2038 9260 2246
rect 9220 2032 9272 2038
rect 9220 1974 9272 1980
rect 9600 800 9628 2314
rect 10060 800 10088 2746
rect 10152 2514 10180 4134
rect 10244 4078 10272 4712
rect 10324 4694 10376 4700
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 10244 3194 10272 3334
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10336 3097 10364 4218
rect 10322 3088 10378 3097
rect 10428 3058 10456 5607
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10704 5370 10732 5510
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10598 5128 10654 5137
rect 10520 4282 10548 5102
rect 10598 5063 10654 5072
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10520 3913 10548 4082
rect 10506 3904 10562 3913
rect 10506 3839 10562 3848
rect 10612 3641 10640 5063
rect 10796 4758 10824 6310
rect 11072 6304 11100 7822
rect 11164 7818 11192 9959
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11704 9376 11756 9382
rect 11808 9364 11836 11630
rect 11900 9518 11928 11698
rect 11992 11694 12020 11727
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 11992 10985 12020 11630
rect 11978 10976 12034 10985
rect 11978 10911 12034 10920
rect 11978 10704 12034 10713
rect 12084 10690 12112 12022
rect 12360 11898 12388 12174
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12544 11558 12572 12174
rect 12624 11620 12676 11626
rect 12624 11562 12676 11568
rect 12532 11552 12584 11558
rect 12532 11494 12584 11500
rect 12636 11286 12664 11562
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12622 11112 12678 11121
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12176 10713 12204 11018
rect 12034 10662 12112 10690
rect 12162 10704 12218 10713
rect 11978 10639 12034 10648
rect 12162 10639 12218 10648
rect 12176 10554 12204 10639
rect 11992 10526 12204 10554
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11808 9336 11928 9364
rect 11704 9318 11756 9324
rect 11716 9042 11744 9318
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11336 7880 11388 7886
rect 11334 7848 11336 7857
rect 11388 7848 11390 7857
rect 11152 7812 11204 7818
rect 11334 7783 11390 7792
rect 11152 7754 11204 7760
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11716 7206 11744 7278
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11716 7041 11744 7142
rect 11702 7032 11758 7041
rect 11702 6967 11758 6976
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 10980 6276 11100 6304
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 10888 5914 10916 6190
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10874 5808 10930 5817
rect 10874 5743 10930 5752
rect 10888 5642 10916 5743
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10888 4826 10916 5170
rect 10980 5098 11008 6276
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 11072 5681 11100 6122
rect 11058 5672 11114 5681
rect 11058 5607 11114 5616
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10784 4752 10836 4758
rect 10784 4694 10836 4700
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10888 4298 10916 4558
rect 10796 4270 10916 4298
rect 10690 4176 10746 4185
rect 10690 4111 10746 4120
rect 10598 3632 10654 3641
rect 10704 3602 10732 4111
rect 10598 3567 10654 3576
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10322 3023 10378 3032
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10796 2514 10824 4270
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10888 3738 10916 4082
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10520 870 10640 898
rect 10520 800 10548 870
rect 3712 734 3924 762
rect 4066 0 4122 800
rect 4526 0 4582 800
rect 4986 0 5042 800
rect 5446 0 5502 800
rect 5906 0 5962 800
rect 6366 0 6422 800
rect 6826 0 6882 800
rect 7286 0 7342 800
rect 7746 0 7802 800
rect 8206 0 8262 800
rect 8666 0 8722 800
rect 9126 0 9182 800
rect 9586 0 9642 800
rect 10046 0 10102 800
rect 10506 0 10562 800
rect 10612 762 10640 870
rect 10796 762 10824 2450
rect 10876 2440 10928 2446
rect 10980 2428 11008 4694
rect 11072 4321 11100 5510
rect 11058 4312 11114 4321
rect 11058 4247 11114 4256
rect 11072 4214 11100 4247
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 11164 2650 11192 6598
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 11334 6080 11390 6089
rect 11334 6015 11390 6024
rect 11348 5574 11376 6015
rect 11532 5778 11560 6258
rect 11716 6118 11744 6802
rect 11808 6361 11836 7686
rect 11794 6352 11850 6361
rect 11794 6287 11850 6296
rect 11796 6248 11848 6254
rect 11796 6190 11848 6196
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11624 5778 11652 6054
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11808 5710 11836 6190
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11336 5568 11388 5574
rect 11900 5556 11928 9336
rect 11336 5510 11388 5516
rect 11808 5528 11928 5556
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 11426 5264 11482 5273
rect 11426 5199 11482 5208
rect 11334 4856 11390 4865
rect 11440 4826 11468 5199
rect 11612 5092 11664 5098
rect 11612 5034 11664 5040
rect 11334 4791 11390 4800
rect 11428 4820 11480 4826
rect 11348 4758 11376 4791
rect 11428 4762 11480 4768
rect 11624 4758 11652 5034
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11612 4752 11664 4758
rect 11612 4694 11664 4700
rect 11348 4554 11376 4694
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 11348 3913 11376 4014
rect 11334 3904 11390 3913
rect 11334 3839 11390 3848
rect 11518 3768 11574 3777
rect 11518 3703 11574 3712
rect 11532 3602 11560 3703
rect 11624 3602 11652 4218
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 11716 3058 11744 4422
rect 11808 3058 11836 5528
rect 11886 5400 11942 5409
rect 11886 5335 11942 5344
rect 11900 5001 11928 5335
rect 11992 5166 12020 10526
rect 12164 9376 12216 9382
rect 12164 9318 12216 9324
rect 12176 8498 12204 9318
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 12084 7546 12112 7686
rect 12072 7540 12124 7546
rect 12072 7482 12124 7488
rect 12176 7426 12204 8434
rect 12084 7398 12204 7426
rect 12084 7002 12112 7398
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12070 6216 12126 6225
rect 12070 6151 12126 6160
rect 12084 5817 12112 6151
rect 12070 5808 12126 5817
rect 12070 5743 12126 5752
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 11980 5160 12032 5166
rect 11980 5102 12032 5108
rect 11980 5024 12032 5030
rect 11886 4992 11942 5001
rect 11980 4966 12032 4972
rect 11886 4927 11942 4936
rect 11992 4826 12020 4966
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 11900 4282 11928 4762
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11992 4282 12020 4422
rect 11888 4276 11940 4282
rect 11888 4218 11940 4224
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11992 3777 12020 4218
rect 12084 4049 12112 5238
rect 12070 4040 12126 4049
rect 12070 3975 12126 3984
rect 11978 3768 12034 3777
rect 11978 3703 12034 3712
rect 11888 3460 11940 3466
rect 11888 3402 11940 3408
rect 11900 3194 11928 3402
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 10928 2400 11008 2428
rect 10876 2382 10928 2388
rect 10980 800 11008 2400
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 11072 2106 11100 2382
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11060 2100 11112 2106
rect 11060 2042 11112 2048
rect 11440 870 11560 898
rect 11440 800 11468 870
rect 10612 734 10824 762
rect 10966 0 11022 800
rect 11426 0 11482 800
rect 11532 762 11560 870
rect 11716 762 11744 2994
rect 12176 2378 12204 7142
rect 12268 5386 12296 11086
rect 12622 11047 12678 11056
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12360 8106 12388 9454
rect 12452 8242 12480 10746
rect 12544 9722 12572 10950
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12636 9586 12664 11047
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12544 9353 12572 9522
rect 12530 9344 12586 9353
rect 12530 9279 12586 9288
rect 12532 8900 12584 8906
rect 12532 8842 12584 8848
rect 12544 8809 12572 8842
rect 12530 8800 12586 8809
rect 12530 8735 12586 8744
rect 12452 8214 12572 8242
rect 12360 8078 12480 8106
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12360 7857 12388 7890
rect 12346 7848 12402 7857
rect 12346 7783 12402 7792
rect 12452 7206 12480 8078
rect 12544 7886 12572 8214
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12544 7018 12572 7686
rect 12452 6990 12572 7018
rect 12452 6662 12480 6990
rect 12636 6882 12664 9522
rect 12728 8294 12756 12582
rect 12820 11354 12848 13262
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12820 10674 12848 10746
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12912 9081 12940 13874
rect 13280 13190 13308 17206
rect 13268 13184 13320 13190
rect 13268 13126 13320 13132
rect 13280 12986 13308 13126
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 13004 12170 13032 12582
rect 13372 12434 13400 20046
rect 13728 19994 13780 20000
rect 13452 19984 13504 19990
rect 13452 19926 13504 19932
rect 13464 19718 13492 19926
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 13556 19310 13584 19858
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 14108 19718 14136 19790
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13452 19236 13504 19242
rect 13452 19178 13504 19184
rect 13464 18834 13492 19178
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13464 18290 13492 18770
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13648 16810 13676 19654
rect 13818 19136 13874 19145
rect 13818 19071 13874 19080
rect 13832 18290 13860 19071
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13726 18048 13782 18057
rect 13726 17983 13782 17992
rect 13740 17882 13768 17983
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 13464 16782 13676 16810
rect 13464 15162 13492 16782
rect 13636 16652 13688 16658
rect 13740 16640 13768 17206
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 13688 16612 13768 16640
rect 13636 16594 13688 16600
rect 13648 16454 13676 16594
rect 14292 16454 14320 20567
rect 14556 20538 14608 20544
rect 14648 20528 14700 20534
rect 14648 20470 14700 20476
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14384 16998 14412 17138
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 13648 16114 13676 16390
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13648 15570 13676 16050
rect 14292 16017 14320 16390
rect 14278 16008 14334 16017
rect 14278 15943 14334 15952
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 13648 15366 13676 15506
rect 14476 15473 14504 19790
rect 14568 19786 14596 20402
rect 14660 20369 14688 20470
rect 14646 20360 14702 20369
rect 14936 20330 14964 22200
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 15212 20466 15240 20946
rect 15396 20602 15424 22200
rect 15856 20602 15884 22200
rect 16316 20602 16344 22200
rect 16776 20890 16804 22200
rect 16776 20862 16988 20890
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 16304 20596 16356 20602
rect 16304 20538 16356 20544
rect 16026 20496 16082 20505
rect 15200 20460 15252 20466
rect 16026 20431 16028 20440
rect 15200 20402 15252 20408
rect 16080 20431 16082 20440
rect 16028 20402 16080 20408
rect 16960 20330 16988 20862
rect 17236 20602 17264 22200
rect 17696 20618 17724 22200
rect 17696 20602 18000 20618
rect 18156 20602 18184 22200
rect 18616 20602 18644 22200
rect 17224 20596 17276 20602
rect 17696 20596 18012 20602
rect 17696 20590 17960 20596
rect 17224 20538 17276 20544
rect 17960 20538 18012 20544
rect 18144 20596 18196 20602
rect 18144 20538 18196 20544
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 18236 20460 18288 20466
rect 18236 20402 18288 20408
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 14646 20295 14702 20304
rect 14924 20324 14976 20330
rect 14924 20266 14976 20272
rect 16948 20324 17000 20330
rect 16948 20266 17000 20272
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 14832 19712 14884 19718
rect 14832 19654 14884 19660
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 14648 19236 14700 19242
rect 14648 19178 14700 19184
rect 14660 18766 14688 19178
rect 14648 18760 14700 18766
rect 14648 18702 14700 18708
rect 14660 18358 14688 18702
rect 14648 18352 14700 18358
rect 14648 18294 14700 18300
rect 14648 18080 14700 18086
rect 14648 18022 14700 18028
rect 14660 17338 14688 18022
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14462 15464 14518 15473
rect 13728 15428 13780 15434
rect 14462 15399 14518 15408
rect 14556 15428 14608 15434
rect 13728 15370 13780 15376
rect 14556 15370 14608 15376
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13648 14890 13676 15302
rect 13636 14884 13688 14890
rect 13636 14826 13688 14832
rect 13648 14482 13676 14826
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13556 12918 13584 14214
rect 13544 12912 13596 12918
rect 13544 12854 13596 12860
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13188 12406 13400 12434
rect 13464 12434 13492 12582
rect 13464 12406 13676 12434
rect 12992 12164 13044 12170
rect 12992 12106 13044 12112
rect 12992 10532 13044 10538
rect 12992 10474 13044 10480
rect 12898 9072 12954 9081
rect 12898 9007 12954 9016
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12820 7954 12848 8026
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12728 7342 12756 7822
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12544 6854 12664 6882
rect 12728 6866 12756 7278
rect 13004 7177 13032 10474
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 12990 7168 13046 7177
rect 12990 7103 13046 7112
rect 12716 6860 12768 6866
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12440 6180 12492 6186
rect 12440 6122 12492 6128
rect 12452 5545 12480 6122
rect 12544 5953 12572 6854
rect 12716 6802 12768 6808
rect 12992 6656 13044 6662
rect 12992 6598 13044 6604
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12530 5944 12586 5953
rect 12530 5879 12586 5888
rect 12636 5817 12664 6258
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12728 6118 12756 6190
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12622 5808 12678 5817
rect 12622 5743 12678 5752
rect 12438 5536 12494 5545
rect 12438 5471 12494 5480
rect 12268 5358 12480 5386
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 12360 2446 12388 4014
rect 12452 2650 12480 5358
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12544 5001 12572 5102
rect 12530 4992 12586 5001
rect 12530 4927 12586 4936
rect 12636 4865 12664 5170
rect 12728 5166 12756 6054
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 12912 5574 12940 5850
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 12820 5370 12848 5510
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12622 4856 12678 4865
rect 12622 4791 12624 4800
rect 12676 4791 12678 4800
rect 12624 4762 12676 4768
rect 12636 4554 12664 4762
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 12728 4486 12756 5102
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12912 4162 12940 4966
rect 13004 4282 13032 6598
rect 13096 5778 13124 10406
rect 13188 9874 13216 12406
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13280 11014 13308 11494
rect 13358 11248 13414 11257
rect 13358 11183 13414 11192
rect 13372 11014 13400 11183
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13280 10606 13308 10950
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13280 10130 13308 10542
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 13188 9846 13308 9874
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13084 5772 13136 5778
rect 13084 5714 13136 5720
rect 12992 4276 13044 4282
rect 12992 4218 13044 4224
rect 12912 4134 13032 4162
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12636 3505 12664 3878
rect 12622 3496 12678 3505
rect 12622 3431 12678 3440
rect 12636 3194 12664 3431
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12912 2514 12940 3878
rect 13004 3398 13032 4134
rect 13188 3618 13216 9658
rect 13280 9353 13308 9846
rect 13266 9344 13322 9353
rect 13266 9279 13322 9288
rect 13266 8800 13322 8809
rect 13266 8735 13322 8744
rect 13280 6662 13308 8735
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13280 5914 13308 6258
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13096 3602 13216 3618
rect 13280 3602 13308 5714
rect 13372 5370 13400 10746
rect 13464 10130 13492 12038
rect 13556 10169 13584 12038
rect 13648 11762 13676 12406
rect 13740 12374 13768 15370
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13832 14414 13860 15302
rect 14280 14884 14332 14890
rect 14280 14826 14332 14832
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 13912 14476 13964 14482
rect 13912 14418 13964 14424
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13924 14260 13952 14418
rect 13832 14232 13952 14260
rect 13832 13938 13860 14232
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13832 13802 13860 13874
rect 13820 13796 13872 13802
rect 13820 13738 13872 13744
rect 13832 13172 13860 13738
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 14096 13184 14148 13190
rect 13832 13144 14096 13172
rect 14096 13126 14148 13132
rect 14108 12850 14136 13126
rect 14292 13002 14320 14826
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14384 13161 14412 14758
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14476 14074 14504 14214
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14370 13152 14426 13161
rect 14370 13087 14426 13096
rect 14200 12986 14504 13002
rect 14188 12980 14504 12986
rect 14240 12974 14504 12980
rect 14188 12922 14240 12928
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 13728 12368 13780 12374
rect 13728 12310 13780 12316
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 13542 10160 13598 10169
rect 13452 10124 13504 10130
rect 13542 10095 13598 10104
rect 13452 10066 13504 10072
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13464 9110 13492 9318
rect 13648 9178 13676 11698
rect 13740 10577 13768 12310
rect 14188 12096 14240 12102
rect 14292 12084 14320 12786
rect 14476 12434 14504 12974
rect 14240 12056 14320 12084
rect 14384 12406 14504 12434
rect 14188 12038 14240 12044
rect 14200 11694 14228 12038
rect 14188 11688 14240 11694
rect 14240 11648 14320 11676
rect 14188 11630 14240 11636
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 14292 11218 14320 11648
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 13726 10568 13782 10577
rect 13726 10503 13782 10512
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13464 8072 13492 9046
rect 13556 8634 13584 9046
rect 13636 8832 13688 8838
rect 13634 8800 13636 8809
rect 13688 8800 13690 8809
rect 13634 8735 13690 8744
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13740 8430 13768 9862
rect 13832 9722 13860 10406
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 14280 9988 14332 9994
rect 14280 9930 14332 9936
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13832 8974 13860 9454
rect 13924 9382 13952 9590
rect 14292 9382 14320 9930
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 13820 8968 13872 8974
rect 13820 8910 13872 8916
rect 13832 8634 13860 8910
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13464 8044 13584 8072
rect 13450 7984 13506 7993
rect 13450 7919 13506 7928
rect 13464 7546 13492 7919
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13556 7392 13584 8044
rect 13464 7364 13584 7392
rect 13464 6089 13492 7364
rect 13542 7304 13598 7313
rect 13542 7239 13598 7248
rect 13556 6186 13584 7239
rect 13544 6180 13596 6186
rect 13544 6122 13596 6128
rect 13450 6080 13506 6089
rect 13450 6015 13506 6024
rect 13648 5778 13676 8298
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13372 5001 13400 5306
rect 13452 5024 13504 5030
rect 13358 4992 13414 5001
rect 13452 4966 13504 4972
rect 13358 4927 13414 4936
rect 13084 3596 13216 3602
rect 13136 3590 13216 3596
rect 13268 3596 13320 3602
rect 13084 3538 13136 3544
rect 13268 3538 13320 3544
rect 12992 3392 13044 3398
rect 12992 3334 13044 3340
rect 13004 2990 13032 3334
rect 13096 3233 13124 3538
rect 13082 3224 13138 3233
rect 13082 3159 13138 3168
rect 13096 3126 13124 3159
rect 13084 3120 13136 3126
rect 13084 3062 13136 3068
rect 13464 3058 13492 4966
rect 13556 3058 13584 5510
rect 13740 4706 13768 7754
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14292 7546 14320 7686
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13832 7002 13860 7210
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 14004 6928 14056 6934
rect 14004 6870 14056 6876
rect 14016 6254 14044 6870
rect 14384 6769 14412 12406
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14476 8906 14504 10202
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 14370 6760 14426 6769
rect 14370 6695 14426 6704
rect 14280 6656 14332 6662
rect 14280 6598 14332 6604
rect 14004 6248 14056 6254
rect 14004 6190 14056 6196
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 13648 4678 13768 4706
rect 13648 4078 13676 4678
rect 13726 4584 13782 4593
rect 13726 4519 13782 4528
rect 13740 4486 13768 4519
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13818 3768 13874 3777
rect 13945 3771 14253 3780
rect 13818 3703 13820 3712
rect 13872 3703 13874 3712
rect 14096 3732 14148 3738
rect 13820 3674 13872 3680
rect 14096 3674 14148 3680
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12900 2508 12952 2514
rect 12900 2450 12952 2456
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12164 2372 12216 2378
rect 12164 2314 12216 2320
rect 12360 2258 12388 2382
rect 12268 2230 12388 2258
rect 11900 870 12020 898
rect 11900 800 11928 870
rect 11532 734 11744 762
rect 11886 0 11942 800
rect 11992 762 12020 870
rect 12268 762 12296 2230
rect 12452 2122 12480 2450
rect 13372 2446 13400 2790
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13648 2378 13676 3402
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13740 3058 13768 3334
rect 14108 3058 14136 3674
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 12808 2372 12860 2378
rect 12808 2314 12860 2320
rect 13636 2372 13688 2378
rect 13636 2314 13688 2320
rect 12360 2094 12480 2122
rect 12360 800 12388 2094
rect 12820 800 12848 2314
rect 13268 2304 13320 2310
rect 13268 2246 13320 2252
rect 13280 800 13308 2246
rect 13740 800 13768 2586
rect 13832 2446 13860 2790
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 14188 2576 14240 2582
rect 14188 2518 14240 2524
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 14200 800 14228 2518
rect 14292 2310 14320 6598
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14384 4146 14412 4422
rect 14476 4185 14504 8842
rect 14568 8090 14596 15370
rect 14660 12209 14688 17138
rect 14844 14521 14872 19654
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 16132 17105 16160 18566
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 16224 18086 16252 18226
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16224 17678 16252 18022
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16224 17270 16252 17478
rect 16212 17264 16264 17270
rect 16212 17206 16264 17212
rect 16118 17096 16174 17105
rect 16118 17031 16174 17040
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 15488 16522 15516 16730
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15476 16516 15528 16522
rect 15476 16458 15528 16464
rect 15764 16454 15792 16526
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15752 16448 15804 16454
rect 15752 16390 15804 16396
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 14936 15434 14964 16186
rect 15212 16182 15240 16390
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 15212 16046 15240 16118
rect 15568 16108 15620 16114
rect 15568 16050 15620 16056
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 15212 15484 15240 15982
rect 15580 15910 15608 16050
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 16028 15904 16080 15910
rect 16028 15846 16080 15852
rect 15384 15496 15436 15502
rect 15212 15456 15384 15484
rect 14924 15428 14976 15434
rect 14924 15370 14976 15376
rect 14830 14512 14886 14521
rect 14830 14447 14886 14456
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14844 12850 14872 14350
rect 14936 14006 14964 15370
rect 15212 15026 15240 15456
rect 15384 15438 15436 15444
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15028 14385 15056 14962
rect 15212 14618 15240 14962
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15764 14414 15792 14758
rect 15752 14408 15804 14414
rect 15014 14376 15070 14385
rect 15070 14334 15240 14362
rect 15752 14350 15804 14356
rect 15014 14311 15070 14320
rect 14924 14000 14976 14006
rect 14924 13942 14976 13948
rect 15212 13462 15240 14334
rect 16040 13802 16068 15846
rect 16224 15706 16252 16730
rect 16212 15700 16264 15706
rect 16212 15642 16264 15648
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15948 12918 15976 13126
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 14646 12200 14702 12209
rect 15304 12170 15332 12786
rect 14646 12135 14702 12144
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 15028 11558 15056 12038
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14830 10976 14886 10985
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14660 7970 14688 10950
rect 14830 10911 14886 10920
rect 14568 7942 14688 7970
rect 14740 8016 14792 8022
rect 14740 7958 14792 7964
rect 14462 4176 14518 4185
rect 14372 4140 14424 4146
rect 14462 4111 14518 4120
rect 14372 4082 14424 4088
rect 14568 4026 14596 7942
rect 14752 7546 14780 7958
rect 14740 7540 14792 7546
rect 14740 7482 14792 7488
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14752 6866 14780 7346
rect 14844 7188 14872 10911
rect 14924 8560 14976 8566
rect 14924 8502 14976 8508
rect 14936 7342 14964 8502
rect 15028 7857 15056 11494
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15212 10742 15240 11154
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15120 9586 15148 10610
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15120 8634 15148 9522
rect 15212 8974 15240 9522
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15014 7848 15070 7857
rect 15014 7783 15070 7792
rect 15120 7546 15148 8026
rect 15212 7732 15240 8774
rect 15304 7886 15332 11086
rect 15382 10704 15438 10713
rect 15382 10639 15384 10648
rect 15436 10639 15438 10648
rect 15384 10610 15436 10616
rect 15488 8809 15516 11494
rect 15936 11348 15988 11354
rect 16040 11336 16068 13738
rect 15988 11308 16068 11336
rect 16120 11348 16172 11354
rect 15936 11290 15988 11296
rect 16120 11290 16172 11296
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15580 9926 15608 11018
rect 15936 9988 15988 9994
rect 15936 9930 15988 9936
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15474 8800 15530 8809
rect 15474 8735 15530 8744
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15212 7704 15332 7732
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 15212 7188 15240 7346
rect 14844 7160 15240 7188
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14844 6662 14872 7160
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 14738 5536 14794 5545
rect 14738 5471 14794 5480
rect 14752 4622 14780 5471
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 14844 4690 14872 4966
rect 14832 4684 14884 4690
rect 14832 4626 14884 4632
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14384 3998 14596 4026
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 14384 2106 14412 3998
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 14556 3664 14608 3670
rect 14556 3606 14608 3612
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 14476 2446 14504 2790
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 14568 2378 14596 3606
rect 14936 3058 14964 3878
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14740 2916 14792 2922
rect 14740 2858 14792 2864
rect 14752 2446 14780 2858
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 14556 2372 14608 2378
rect 14556 2314 14608 2320
rect 14740 2304 14792 2310
rect 14660 2264 14740 2292
rect 14372 2100 14424 2106
rect 14372 2042 14424 2048
rect 14660 800 14688 2264
rect 14740 2246 14792 2252
rect 15028 1970 15056 6598
rect 15304 3641 15332 7704
rect 15580 6458 15608 9862
rect 15672 9654 15700 9862
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15672 6186 15700 9590
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15764 8634 15792 8910
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15660 6180 15712 6186
rect 15660 6122 15712 6128
rect 15566 5672 15622 5681
rect 15566 5607 15622 5616
rect 15580 5166 15608 5607
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15568 5160 15620 5166
rect 15764 5137 15792 7686
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15856 5234 15884 6054
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 15568 5102 15620 5108
rect 15750 5128 15806 5137
rect 15488 4826 15516 5102
rect 15750 5063 15806 5072
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 15948 4622 15976 9930
rect 16132 9178 16160 11290
rect 16224 9489 16252 14554
rect 16316 11898 16344 19654
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 17052 19530 17080 20402
rect 16960 19502 17080 19530
rect 16960 19174 16988 19502
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 16408 17814 16436 18566
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 16960 18290 16988 18702
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16396 17808 16448 17814
rect 16396 17750 16448 17756
rect 16592 17678 16620 18226
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 17052 17610 17080 19314
rect 17144 18970 17172 20402
rect 17788 20058 17816 20402
rect 17776 20052 17828 20058
rect 17776 19994 17828 20000
rect 18248 19446 18276 20402
rect 18328 20392 18380 20398
rect 18328 20334 18380 20340
rect 18236 19440 18288 19446
rect 18236 19382 18288 19388
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 17696 18766 17724 19110
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 18144 18692 18196 18698
rect 18144 18634 18196 18640
rect 18156 18578 18184 18634
rect 18156 18550 18276 18578
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 16396 17604 16448 17610
rect 16396 17546 16448 17552
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 16408 15910 16436 17546
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16488 17128 16540 17134
rect 16488 17070 16540 17076
rect 16500 16590 16528 17070
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16408 15434 16436 15846
rect 16396 15428 16448 15434
rect 16396 15370 16448 15376
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16960 15094 16988 17138
rect 17420 16998 17448 18226
rect 18156 18170 18184 18226
rect 17788 18142 18184 18170
rect 17788 17814 17816 18142
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 18144 18080 18196 18086
rect 18248 18034 18276 18550
rect 18196 18028 18276 18034
rect 18144 18022 18276 18028
rect 17776 17808 17828 17814
rect 17774 17776 17776 17785
rect 17828 17776 17830 17785
rect 17774 17711 17830 17720
rect 17880 17678 17908 18022
rect 18156 18006 18276 18022
rect 17868 17672 17920 17678
rect 18156 17626 18184 18006
rect 18340 17882 18368 20334
rect 18708 19961 18736 20402
rect 19076 19990 19104 22200
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 19536 19990 19564 22200
rect 19616 20460 19668 20466
rect 19616 20402 19668 20408
rect 19628 20058 19656 20402
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 19064 19984 19116 19990
rect 18694 19952 18750 19961
rect 19064 19926 19116 19932
rect 19524 19984 19576 19990
rect 19524 19926 19576 19932
rect 18694 19887 18750 19896
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19996 19802 20024 22200
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 19536 18737 19564 19790
rect 19996 19774 20116 19802
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 19522 18728 19578 18737
rect 19522 18663 19578 18672
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19536 18154 19564 18362
rect 19628 18358 19656 19654
rect 19996 19446 20024 19654
rect 20088 19514 20116 19774
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 19984 19440 20036 19446
rect 19984 19382 20036 19388
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 19904 18426 19932 19314
rect 20076 18624 20128 18630
rect 20076 18566 20128 18572
rect 19892 18420 19944 18426
rect 19892 18362 19944 18368
rect 19616 18352 19668 18358
rect 19616 18294 19668 18300
rect 19524 18148 19576 18154
rect 19524 18090 19576 18096
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 18328 17876 18380 17882
rect 18328 17818 18380 17824
rect 17868 17614 17920 17620
rect 17880 17338 17908 17614
rect 18064 17598 18184 17626
rect 20088 17610 20116 18566
rect 20076 17604 20128 17610
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17880 16810 17908 17274
rect 17880 16794 18000 16810
rect 17880 16788 18012 16794
rect 17880 16782 17960 16788
rect 17960 16730 18012 16736
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 16948 15088 17000 15094
rect 16948 15030 17000 15036
rect 17604 15008 17632 15438
rect 17684 15020 17736 15026
rect 17604 14980 17684 15008
rect 17604 14414 17632 14980
rect 17684 14962 17736 14968
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17500 14340 17552 14346
rect 17500 14282 17552 14288
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 17512 14074 17540 14282
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 16394 13832 16450 13841
rect 16394 13767 16450 13776
rect 16408 12918 16436 13767
rect 17328 13530 17356 13874
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 16684 12306 16712 12786
rect 17038 12744 17094 12753
rect 17038 12679 17094 12688
rect 16672 12300 16724 12306
rect 16408 12260 16672 12288
rect 16304 11892 16356 11898
rect 16408 11880 16436 12260
rect 16672 12242 16724 12248
rect 17052 12238 17080 12679
rect 17512 12434 17540 14010
rect 17604 13530 17632 14350
rect 17972 13870 18000 16458
rect 18064 16153 18092 17598
rect 20076 17546 20128 17552
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 18050 16144 18106 16153
rect 18050 16079 18106 16088
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17604 12986 17632 13466
rect 17684 13320 17736 13326
rect 17972 13297 18000 13806
rect 17684 13262 17736 13268
rect 17958 13288 18014 13297
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 17696 12714 17724 13262
rect 18064 13258 18092 14758
rect 18156 14618 18184 17070
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 18236 16516 18288 16522
rect 18236 16458 18288 16464
rect 18248 15706 18276 16458
rect 19064 16448 19116 16454
rect 19064 16390 19116 16396
rect 19076 16114 19104 16390
rect 19352 16114 19380 16594
rect 20088 16182 20116 17546
rect 20180 16998 20208 19654
rect 20456 19446 20484 22200
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 20824 19786 20852 20334
rect 20812 19780 20864 19786
rect 20812 19722 20864 19728
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20718 19408 20774 19417
rect 20718 19343 20720 19352
rect 20772 19343 20774 19352
rect 20720 19314 20772 19320
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20364 16998 20392 18702
rect 20444 18692 20496 18698
rect 20444 18634 20496 18640
rect 20456 18290 20484 18634
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 20732 17241 20760 19110
rect 20824 18766 20852 19722
rect 20916 18970 20944 22200
rect 21376 20058 21404 22200
rect 21836 20890 21864 22200
rect 21652 20862 21864 20890
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 21178 19816 21234 19825
rect 21178 19751 21234 19760
rect 21272 19780 21324 19786
rect 21192 19378 21220 19751
rect 21272 19722 21324 19728
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 21284 19258 21312 19722
rect 21192 19230 21312 19258
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 20994 18864 21050 18873
rect 20994 18799 21050 18808
rect 21008 18766 21036 18799
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 20824 18426 20852 18702
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 21192 17542 21220 19230
rect 21652 18426 21680 20862
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 22296 20466 22324 22200
rect 22756 20534 22784 22200
rect 22744 20528 22796 20534
rect 22744 20470 22796 20476
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 21640 18420 21692 18426
rect 21640 18362 21692 18368
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 20718 17232 20774 17241
rect 20718 17167 20774 17176
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20076 16176 20128 16182
rect 20076 16118 20128 16124
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 19076 14929 19104 16050
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19812 15094 19840 15302
rect 19800 15088 19852 15094
rect 19800 15030 19852 15036
rect 19800 14952 19852 14958
rect 19062 14920 19118 14929
rect 19800 14894 19852 14900
rect 19062 14855 19118 14864
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 18340 13938 18368 14758
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19812 14278 19840 14894
rect 20364 14346 20392 16934
rect 21192 16561 21220 17478
rect 21284 17241 21312 17614
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21468 17241 21496 17478
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21270 17232 21326 17241
rect 21270 17167 21326 17176
rect 21454 17232 21510 17241
rect 21454 17167 21510 17176
rect 21456 16584 21508 16590
rect 21178 16552 21234 16561
rect 21456 16526 21508 16532
rect 21178 16487 21234 16496
rect 21468 16114 21496 16526
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 20628 15360 20680 15366
rect 20628 15302 20680 15308
rect 20352 14340 20404 14346
rect 20352 14282 20404 14288
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 18328 13932 18380 13938
rect 18328 13874 18380 13880
rect 17958 13223 18014 13232
rect 18052 13252 18104 13258
rect 18052 13194 18104 13200
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17684 12708 17736 12714
rect 17684 12650 17736 12656
rect 17880 12442 17908 12922
rect 17420 12406 17540 12434
rect 17868 12436 17920 12442
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16408 11852 16528 11880
rect 16304 11834 16356 11840
rect 16500 11762 16528 11852
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16408 11218 16436 11698
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16500 11354 16528 11562
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16948 11280 17000 11286
rect 16948 11222 17000 11228
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16500 9994 16528 10406
rect 16488 9988 16540 9994
rect 16488 9930 16540 9936
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16210 9480 16266 9489
rect 16210 9415 16266 9424
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 16210 9072 16266 9081
rect 16210 9007 16266 9016
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 16040 6730 16068 7686
rect 16028 6724 16080 6730
rect 16028 6666 16080 6672
rect 16026 5400 16082 5409
rect 16132 5386 16160 8570
rect 16082 5358 16160 5386
rect 16026 5335 16082 5344
rect 16040 4690 16068 5335
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 15856 4185 15884 4422
rect 15948 4282 15976 4422
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 15842 4176 15898 4185
rect 15842 4111 15898 4120
rect 15856 4010 15884 4111
rect 15844 4004 15896 4010
rect 15844 3946 15896 3952
rect 16224 3670 16252 9007
rect 16408 8838 16436 9862
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16670 9616 16726 9625
rect 16670 9551 16726 9560
rect 16684 9450 16712 9551
rect 16672 9444 16724 9450
rect 16672 9386 16724 9392
rect 16960 8906 16988 11222
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 17052 9586 17080 9998
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 17420 8945 17448 12406
rect 17868 12378 17920 12384
rect 18340 12345 18368 13874
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 19536 13530 19564 13806
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 18972 13456 19024 13462
rect 18970 13424 18972 13433
rect 19024 13424 19026 13433
rect 18970 13359 19026 13368
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 19536 12434 19564 12582
rect 19536 12406 19748 12434
rect 18326 12336 18382 12345
rect 18236 12300 18288 12306
rect 18326 12271 18382 12280
rect 18236 12242 18288 12248
rect 18248 11558 18276 12242
rect 19524 12164 19576 12170
rect 19524 12106 19576 12112
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 17960 11076 18012 11082
rect 17960 11018 18012 11024
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 17406 8936 17462 8945
rect 16948 8900 17000 8906
rect 17406 8871 17462 8880
rect 16948 8842 17000 8848
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 16486 6352 16542 6361
rect 16486 6287 16542 6296
rect 16500 5710 16528 6287
rect 16580 5840 16632 5846
rect 16580 5782 16632 5788
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16592 5574 16620 5782
rect 16960 5681 16988 8842
rect 17512 8838 17540 10678
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17788 10062 17816 10406
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 16946 5672 17002 5681
rect 16946 5607 17002 5616
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 17040 5024 17092 5030
rect 17040 4966 17092 4972
rect 16948 4752 17000 4758
rect 16948 4694 17000 4700
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 16316 4321 16344 4558
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16302 4312 16358 4321
rect 16544 4315 16852 4324
rect 16302 4247 16358 4256
rect 16316 4146 16344 4247
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16212 3664 16264 3670
rect 15290 3632 15346 3641
rect 16212 3606 16264 3612
rect 15290 3567 15346 3576
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 15934 3224 15990 3233
rect 16544 3227 16852 3236
rect 15934 3159 15990 3168
rect 16120 3188 16172 3194
rect 15948 3126 15976 3159
rect 16120 3130 16172 3136
rect 15936 3120 15988 3126
rect 15106 3088 15162 3097
rect 15936 3062 15988 3068
rect 15106 3023 15108 3032
rect 15160 3023 15162 3032
rect 15108 2994 15160 3000
rect 15292 2916 15344 2922
rect 15292 2858 15344 2864
rect 15304 2446 15332 2858
rect 16132 2446 16160 3130
rect 16764 2916 16816 2922
rect 16764 2858 16816 2864
rect 16672 2848 16724 2854
rect 16672 2790 16724 2796
rect 16684 2650 16712 2790
rect 16672 2644 16724 2650
rect 16672 2586 16724 2592
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16776 2378 16804 2858
rect 16960 2446 16988 4694
rect 17052 3058 17080 4966
rect 17130 4584 17186 4593
rect 17130 4519 17186 4528
rect 17144 3126 17172 4519
rect 17236 4146 17264 7482
rect 17328 5148 17356 7686
rect 17420 5273 17448 7686
rect 17406 5264 17462 5273
rect 17406 5199 17462 5208
rect 17328 5120 17448 5148
rect 17420 4729 17448 5120
rect 17512 4826 17540 8774
rect 17592 8084 17644 8090
rect 17592 8026 17644 8032
rect 17604 5778 17632 8026
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17592 5772 17644 5778
rect 17592 5714 17644 5720
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17406 4720 17462 4729
rect 17604 4690 17632 5714
rect 17696 5250 17724 7686
rect 17788 6934 17816 9998
rect 17880 9625 17908 10610
rect 17866 9616 17922 9625
rect 17866 9551 17922 9560
rect 17868 9376 17920 9382
rect 17972 9364 18000 11018
rect 18432 11014 18460 11494
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 18432 10606 18460 10950
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18432 9994 18460 10542
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 18052 9988 18104 9994
rect 18052 9930 18104 9936
rect 18420 9988 18472 9994
rect 18420 9930 18472 9936
rect 18064 9518 18092 9930
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 17920 9336 18000 9364
rect 17868 9318 17920 9324
rect 17972 8634 18000 9336
rect 18064 8974 18092 9454
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 18064 8498 18092 8910
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17776 6928 17828 6934
rect 17776 6870 17828 6876
rect 17880 6798 17908 7686
rect 18248 7478 18276 9522
rect 18524 8362 18552 9862
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19536 8838 19564 12106
rect 19616 11552 19668 11558
rect 19616 11494 19668 11500
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19430 8528 19486 8537
rect 19430 8463 19432 8472
rect 19484 8463 19486 8472
rect 19432 8434 19484 8440
rect 18512 8356 18564 8362
rect 18512 8298 18564 8304
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18236 7472 18288 7478
rect 18236 7414 18288 7420
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17788 5370 17816 5510
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 17696 5222 17816 5250
rect 17406 4655 17462 4664
rect 17592 4684 17644 4690
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17236 3738 17264 4082
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17236 3176 17264 3674
rect 17316 3188 17368 3194
rect 17236 3148 17316 3176
rect 17316 3130 17368 3136
rect 17132 3120 17184 3126
rect 17420 3097 17448 4655
rect 17592 4626 17644 4632
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17684 4480 17736 4486
rect 17684 4422 17736 4428
rect 17604 4282 17632 4422
rect 17592 4276 17644 4282
rect 17592 4218 17644 4224
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17604 3670 17632 4082
rect 17592 3664 17644 3670
rect 17592 3606 17644 3612
rect 17132 3062 17184 3068
rect 17406 3088 17462 3097
rect 17040 3052 17092 3058
rect 17406 3023 17462 3032
rect 17040 2994 17092 3000
rect 17500 2916 17552 2922
rect 17500 2858 17552 2864
rect 17132 2848 17184 2854
rect 17132 2790 17184 2796
rect 17144 2446 17172 2790
rect 17512 2446 17540 2858
rect 17696 2514 17724 4422
rect 17684 2508 17736 2514
rect 17684 2450 17736 2456
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 16764 2372 16816 2378
rect 16764 2314 16816 2320
rect 15108 2304 15160 2310
rect 15108 2246 15160 2252
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 15016 1964 15068 1970
rect 15016 1906 15068 1912
rect 15120 800 15148 2246
rect 15580 800 15608 2246
rect 16040 800 16068 2246
rect 16408 1170 16436 2246
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 16408 1142 16528 1170
rect 16500 800 16528 1142
rect 16960 800 16988 2246
rect 17420 800 17448 2246
rect 17788 2038 17816 5222
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17868 4208 17920 4214
rect 17868 4150 17920 4156
rect 17880 3738 17908 4150
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17880 2922 17908 3674
rect 17972 3194 18000 4490
rect 18524 4282 18552 7754
rect 19536 7274 19564 8774
rect 19628 8537 19656 11494
rect 19720 10538 19748 12406
rect 19812 11665 19840 14214
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 20168 13252 20220 13258
rect 20168 13194 20220 13200
rect 19892 13184 19944 13190
rect 19892 13126 19944 13132
rect 19904 12918 19932 13126
rect 19892 12912 19944 12918
rect 19892 12854 19944 12860
rect 20076 12912 20128 12918
rect 20076 12854 20128 12860
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 19798 11656 19854 11665
rect 19798 11591 19854 11600
rect 19800 11076 19852 11082
rect 19800 11018 19852 11024
rect 19708 10532 19760 10538
rect 19708 10474 19760 10480
rect 19812 10470 19840 11018
rect 19800 10464 19852 10470
rect 19800 10406 19852 10412
rect 19614 8528 19670 8537
rect 19614 8463 19670 8472
rect 19812 8022 19840 10406
rect 19904 9926 19932 11698
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19800 8016 19852 8022
rect 19800 7958 19852 7964
rect 19524 7268 19576 7274
rect 19524 7210 19576 7216
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 18788 5840 18840 5846
rect 18788 5782 18840 5788
rect 18800 4622 18828 5782
rect 20088 5778 20116 12854
rect 20180 8090 20208 13194
rect 20272 12170 20300 13874
rect 20260 12164 20312 12170
rect 20260 12106 20312 12112
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20456 7410 20484 8230
rect 20548 7818 20576 9862
rect 20640 8974 20668 15302
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20732 9382 20760 14962
rect 21088 14816 21140 14822
rect 21088 14758 21140 14764
rect 21100 14414 21128 14758
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 20904 14340 20956 14346
rect 20904 14282 20956 14288
rect 20916 13530 20944 14282
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 21100 13274 21128 14350
rect 21192 13410 21220 16050
rect 21468 15502 21496 16050
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 21284 14074 21312 15370
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 21192 13382 21312 13410
rect 21180 13320 21232 13326
rect 21100 13268 21180 13274
rect 21100 13262 21232 13268
rect 21100 13246 21220 13262
rect 21100 12986 21128 13246
rect 21284 13138 21312 13382
rect 21192 13110 21312 13138
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 21008 11830 21036 12038
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 20916 11098 20944 11494
rect 21008 11218 21036 11766
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 20916 11070 21036 11098
rect 20812 9920 20864 9926
rect 20812 9862 20864 9868
rect 20824 9722 20852 9862
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20720 9376 20772 9382
rect 20720 9318 20772 9324
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20640 8634 20668 8910
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20536 7812 20588 7818
rect 20536 7754 20588 7760
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20732 5914 20760 9318
rect 20824 8974 20852 9658
rect 21008 9586 21036 11070
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 20812 8968 20864 8974
rect 20812 8910 20864 8916
rect 20824 8566 20852 8910
rect 20812 8560 20864 8566
rect 20812 8502 20864 8508
rect 20824 8090 20852 8502
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 20824 7546 20852 8026
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 20076 5772 20128 5778
rect 20076 5714 20128 5720
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20812 5568 20864 5574
rect 20812 5510 20864 5516
rect 19522 5264 19578 5273
rect 19522 5199 19578 5208
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 18788 4616 18840 4622
rect 18788 4558 18840 4564
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18524 4078 18552 4218
rect 18512 4072 18564 4078
rect 18512 4014 18564 4020
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 19536 3738 19564 5199
rect 20272 4826 20300 5510
rect 20824 5234 20852 5510
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 19892 4480 19944 4486
rect 19892 4422 19944 4428
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 18880 3664 18932 3670
rect 18880 3606 18932 3612
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 18892 3058 18920 3606
rect 19156 3188 19208 3194
rect 19432 3188 19484 3194
rect 19208 3148 19432 3176
rect 19156 3130 19208 3136
rect 19432 3130 19484 3136
rect 19708 3188 19760 3194
rect 19708 3130 19760 3136
rect 19338 3088 19394 3097
rect 18880 3052 18932 3058
rect 18932 3012 19288 3040
rect 19338 3023 19340 3032
rect 18880 2994 18932 3000
rect 19260 2922 19288 3012
rect 19392 3023 19394 3032
rect 19340 2994 19392 3000
rect 19720 2990 19748 3130
rect 19904 3058 19932 4422
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20364 3058 20392 3674
rect 20732 3058 20760 4966
rect 21008 4010 21036 9522
rect 21192 6458 21220 13110
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21284 12238 21312 12922
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21364 10600 21416 10606
rect 21364 10542 21416 10548
rect 21376 9926 21404 10542
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21560 7886 21588 14010
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21548 7880 21600 7886
rect 21548 7822 21600 7828
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21180 6452 21232 6458
rect 21180 6394 21232 6400
rect 21548 6316 21600 6322
rect 21548 6258 21600 6264
rect 21560 5817 21588 6258
rect 21546 5808 21602 5817
rect 21546 5743 21602 5752
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 21362 4176 21418 4185
rect 21362 4111 21418 4120
rect 20996 4004 21048 4010
rect 20996 3946 21048 3952
rect 21376 3738 21404 4111
rect 21364 3732 21416 3738
rect 21364 3674 21416 3680
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 19892 3052 19944 3058
rect 19892 2994 19944 3000
rect 20352 3052 20404 3058
rect 20352 2994 20404 3000
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 21180 2984 21232 2990
rect 21180 2926 21232 2932
rect 17868 2916 17920 2922
rect 17868 2858 17920 2864
rect 18696 2916 18748 2922
rect 18696 2858 18748 2864
rect 19248 2916 19300 2922
rect 19248 2858 19300 2864
rect 19892 2916 19944 2922
rect 19892 2858 19944 2864
rect 20720 2916 20772 2922
rect 20720 2858 20772 2864
rect 18328 2848 18380 2854
rect 18328 2790 18380 2796
rect 18340 2446 18368 2790
rect 18708 2446 18736 2858
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 19248 2576 19300 2582
rect 19248 2518 19300 2524
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 18788 2304 18840 2310
rect 18788 2246 18840 2252
rect 17776 2032 17828 2038
rect 17776 1974 17828 1980
rect 17880 800 17908 2246
rect 18340 800 18368 2246
rect 18800 800 18828 2246
rect 19260 800 19288 2518
rect 19904 2446 19932 2858
rect 20444 2848 20496 2854
rect 20444 2790 20496 2796
rect 20456 2530 20484 2790
rect 20272 2514 20484 2530
rect 20260 2508 20484 2514
rect 20312 2502 20484 2508
rect 20260 2450 20312 2456
rect 20732 2446 20760 2858
rect 21192 2446 21220 2926
rect 22100 2916 22152 2922
rect 22100 2858 22152 2864
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 19892 2440 19944 2446
rect 19892 2382 19944 2388
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 21180 2440 21232 2446
rect 21180 2382 21232 2388
rect 19708 2304 19760 2310
rect 20260 2304 20312 2310
rect 19708 2246 19760 2252
rect 20180 2264 20260 2292
rect 19720 800 19748 2246
rect 20180 800 20208 2264
rect 20260 2246 20312 2252
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 21088 2304 21140 2310
rect 21088 2246 21140 2252
rect 20640 800 20668 2246
rect 21100 800 21128 2246
rect 21560 800 21588 2790
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 22112 1442 22140 2858
rect 22020 1414 22140 1442
rect 22020 800 22048 1414
rect 22480 800 22508 3470
rect 11992 734 12296 762
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13266 0 13322 800
rect 13726 0 13782 800
rect 14186 0 14242 800
rect 14646 0 14702 800
rect 15106 0 15162 800
rect 15566 0 15622 800
rect 16026 0 16082 800
rect 16486 0 16542 800
rect 16946 0 17002 800
rect 17406 0 17462 800
rect 17866 0 17922 800
rect 18326 0 18382 800
rect 18786 0 18842 800
rect 19246 0 19302 800
rect 19706 0 19762 800
rect 20166 0 20222 800
rect 20626 0 20682 800
rect 21086 0 21142 800
rect 21546 0 21602 800
rect 22006 0 22062 800
rect 22466 0 22522 800
<< via2 >>
rect 1490 20204 1492 20224
rect 1492 20204 1544 20224
rect 1544 20204 1546 20224
rect 1490 20168 1546 20204
rect 1858 20596 1914 20632
rect 1858 20576 1860 20596
rect 1860 20576 1912 20596
rect 1912 20576 1914 20596
rect 2226 20984 2282 21040
rect 1490 19352 1546 19408
rect 1490 18944 1546 19000
rect 1490 18572 1492 18592
rect 1492 18572 1544 18592
rect 1544 18572 1546 18592
rect 1490 18536 1546 18572
rect 1490 17720 1546 17776
rect 1490 17312 1546 17368
rect 1674 17992 1730 18048
rect 1858 19760 1914 19816
rect 1950 19352 2006 19408
rect 2318 19660 2320 19680
rect 2320 19660 2372 19680
rect 2372 19660 2374 19680
rect 2318 19624 2374 19660
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 1858 18148 1914 18184
rect 1858 18128 1860 18148
rect 1860 18128 1912 18148
rect 1912 18128 1914 18148
rect 1490 16940 1492 16960
rect 1492 16940 1544 16960
rect 1544 16940 1546 16960
rect 1490 16904 1546 16940
rect 1490 16088 1546 16144
rect 1490 15680 1546 15736
rect 1490 15308 1492 15328
rect 1492 15308 1544 15328
rect 1544 15308 1546 15328
rect 1490 15272 1546 15308
rect 1490 14456 1546 14512
rect 1490 14048 1546 14104
rect 1490 13676 1492 13696
rect 1492 13676 1544 13696
rect 1544 13676 1546 13696
rect 1490 13640 1546 13676
rect 1490 13232 1546 13288
rect 1398 12844 1454 12880
rect 1398 12824 1400 12844
rect 1400 12824 1452 12844
rect 1452 12824 1454 12844
rect 1398 12008 1454 12064
rect 1398 11600 1454 11656
rect 1398 10784 1454 10840
rect 1398 10376 1454 10432
rect 1398 10004 1400 10024
rect 1400 10004 1452 10024
rect 1452 10004 1454 10024
rect 1398 9968 1454 10004
rect 1858 16496 1914 16552
rect 1674 12416 1730 12472
rect 1858 14884 1914 14920
rect 1858 14864 1860 14884
rect 1860 14864 1912 14884
rect 1912 14864 1914 14884
rect 1674 11192 1730 11248
rect 1582 9968 1638 10024
rect 1674 9560 1730 9616
rect 1398 9152 1454 9208
rect 1674 8744 1730 8800
rect 1398 8336 1454 8392
rect 1398 7928 1454 7984
rect 1398 7520 1454 7576
rect 2686 19488 2742 19544
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 4342 19488 4398 19544
rect 4250 19352 4306 19408
rect 4986 19352 5042 19408
rect 4158 16532 4160 16552
rect 4160 16532 4212 16552
rect 4212 16532 4214 16552
rect 4158 16496 4214 16532
rect 1582 7268 1638 7304
rect 1582 7248 1584 7268
rect 1584 7248 1636 7268
rect 1636 7248 1638 7268
rect 1674 7112 1730 7168
rect 1398 6740 1400 6760
rect 1400 6740 1452 6760
rect 1452 6740 1454 6760
rect 1398 6704 1454 6740
rect 1674 6296 1730 6352
rect 1398 5908 1454 5944
rect 1398 5888 1400 5908
rect 1400 5888 1452 5908
rect 1452 5888 1454 5908
rect 1582 5788 1584 5808
rect 1584 5788 1636 5808
rect 1636 5788 1638 5808
rect 1582 5752 1638 5788
rect 1398 5480 1454 5536
rect 1674 5072 1730 5128
rect 1490 4664 1546 4720
rect 2226 6704 2282 6760
rect 1490 3476 1492 3496
rect 1492 3476 1544 3496
rect 1544 3476 1546 3496
rect 1490 3440 1546 3476
rect 1674 3440 1730 3496
rect 1858 3032 1914 3088
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 2870 10104 2926 10160
rect 2410 9444 2466 9480
rect 2410 9424 2412 9444
rect 2412 9424 2464 9444
rect 2464 9424 2466 9444
rect 2410 7384 2466 7440
rect 2226 4256 2282 4312
rect 2226 3848 2282 3904
rect 3146 10104 3202 10160
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3974 12824 4030 12880
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3790 10124 3846 10160
rect 3790 10104 3792 10124
rect 3792 10104 3844 10124
rect 3844 10104 3846 10124
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3238 8472 3294 8528
rect 2870 8336 2926 8392
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 4066 7792 4122 7848
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 2778 6296 2834 6352
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 2502 3576 2558 3632
rect 2318 3032 2374 3088
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 4618 14592 4674 14648
rect 5170 17584 5226 17640
rect 5262 16088 5318 16144
rect 5078 15544 5134 15600
rect 5078 14320 5134 14376
rect 5722 19352 5778 19408
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 6550 19352 6606 19408
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 6182 17040 6238 17096
rect 5906 16108 5962 16144
rect 5906 16088 5908 16108
rect 5908 16088 5960 16108
rect 5960 16088 5962 16108
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 4710 10376 4766 10432
rect 4710 10104 4766 10160
rect 4986 9424 5042 9480
rect 5262 13232 5318 13288
rect 2778 2624 2834 2680
rect 4710 5208 4766 5264
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 2226 2216 2282 2272
rect 2134 1808 2190 1864
rect 5170 8356 5226 8392
rect 5170 8336 5172 8356
rect 5172 8336 5224 8356
rect 5224 8336 5226 8356
rect 5722 11192 5778 11248
rect 5630 9832 5686 9888
rect 6366 15852 6368 15872
rect 6368 15852 6420 15872
rect 6420 15852 6422 15872
rect 6366 15816 6422 15852
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6274 14456 6330 14512
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6458 13912 6514 13968
rect 6182 13504 6238 13560
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 6550 12960 6606 13016
rect 6550 12280 6606 12336
rect 6734 16224 6790 16280
rect 7470 20304 7526 20360
rect 7010 19352 7066 19408
rect 6918 17720 6974 17776
rect 6918 16088 6974 16144
rect 6734 13504 6790 13560
rect 6826 12552 6882 12608
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6734 12008 6790 12064
rect 5906 9560 5962 9616
rect 5722 7948 5778 7984
rect 5722 7928 5724 7948
rect 5724 7928 5776 7948
rect 5776 7928 5778 7948
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6090 10124 6146 10160
rect 6090 10104 6092 10124
rect 6092 10104 6144 10124
rect 6144 10104 6146 10124
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 5998 9288 6054 9344
rect 6642 10648 6698 10704
rect 7378 12724 7380 12744
rect 7380 12724 7432 12744
rect 7432 12724 7434 12744
rect 7378 12688 7434 12724
rect 7194 11192 7250 11248
rect 7010 10240 7066 10296
rect 6826 9036 6882 9072
rect 6826 9016 6828 9036
rect 6828 9016 6880 9036
rect 6880 9016 6882 9036
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 5446 5752 5502 5808
rect 5262 3984 5318 4040
rect 5906 7384 5962 7440
rect 5814 5616 5870 5672
rect 6090 8336 6146 8392
rect 6366 7928 6422 7984
rect 6550 7928 6606 7984
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6550 6840 6606 6896
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6550 5888 6606 5944
rect 6826 6840 6882 6896
rect 6826 6740 6828 6760
rect 6828 6740 6880 6760
rect 6880 6740 6882 6760
rect 6826 6704 6882 6740
rect 7286 10376 7342 10432
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8574 19896 8630 19952
rect 7746 17176 7802 17232
rect 8298 18400 8354 18456
rect 8206 16224 8262 16280
rect 7746 15988 7748 16008
rect 7748 15988 7800 16008
rect 7800 15988 7802 16008
rect 7746 15952 7802 15988
rect 9218 20440 9274 20496
rect 9218 19352 9274 19408
rect 9034 19216 9090 19272
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 9310 19080 9366 19136
rect 8482 18672 8538 18728
rect 8390 16244 8446 16280
rect 8390 16224 8392 16244
rect 8392 16224 8444 16244
rect 8444 16224 8446 16244
rect 8114 15136 8170 15192
rect 8298 15136 8354 15192
rect 8114 15000 8170 15056
rect 7654 12960 7710 13016
rect 7930 11872 7986 11928
rect 7102 7656 7158 7712
rect 7102 7248 7158 7304
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 7010 6024 7066 6080
rect 6550 5108 6552 5128
rect 6552 5108 6604 5128
rect 6604 5108 6606 5128
rect 6550 5072 6606 5108
rect 7010 5344 7066 5400
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6550 4120 6606 4176
rect 6182 3576 6238 3632
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 7378 3304 7434 3360
rect 7562 6160 7618 6216
rect 7930 10548 7932 10568
rect 7932 10548 7984 10568
rect 7984 10548 7986 10568
rect 7930 10512 7986 10548
rect 9770 19760 9826 19816
rect 9586 19624 9642 19680
rect 9402 18536 9458 18592
rect 9770 18808 9826 18864
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 9402 18028 9404 18048
rect 9404 18028 9456 18048
rect 9456 18028 9458 18048
rect 9402 17992 9458 18028
rect 9586 17992 9642 18048
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 9678 17740 9734 17776
rect 9678 17720 9680 17740
rect 9680 17720 9732 17740
rect 9732 17720 9734 17740
rect 9586 17584 9642 17640
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 9034 15156 9090 15192
rect 9034 15136 9036 15156
rect 9036 15136 9088 15156
rect 9088 15136 9090 15156
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8758 14492 8760 14512
rect 8760 14492 8812 14512
rect 8812 14492 8814 14512
rect 8758 14456 8814 14492
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 9402 15952 9458 16008
rect 9402 15544 9458 15600
rect 9402 15444 9404 15464
rect 9404 15444 9456 15464
rect 9456 15444 9458 15464
rect 9402 15408 9458 15444
rect 9310 14864 9366 14920
rect 8666 13388 8722 13424
rect 8666 13368 8668 13388
rect 8668 13368 8720 13388
rect 8720 13368 8722 13388
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 8298 10104 8354 10160
rect 7746 6024 7802 6080
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 9126 10512 9182 10568
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 8482 9868 8484 9888
rect 8484 9868 8536 9888
rect 8536 9868 8538 9888
rect 8482 9832 8538 9868
rect 8482 9324 8484 9344
rect 8484 9324 8536 9344
rect 8536 9324 8538 9344
rect 8482 9288 8538 9324
rect 8666 9560 8722 9616
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8666 8880 8722 8936
rect 7930 6604 7932 6624
rect 7932 6604 7984 6624
rect 7984 6604 7986 6624
rect 7930 6568 7986 6604
rect 7930 5208 7986 5264
rect 8298 6316 8354 6352
rect 8298 6296 8300 6316
rect 8300 6296 8352 6316
rect 8352 6296 8354 6316
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8574 6296 8630 6352
rect 8390 6024 8446 6080
rect 8298 5616 8354 5672
rect 8022 4528 8078 4584
rect 8114 3984 8170 4040
rect 7746 3712 7802 3768
rect 7654 3032 7710 3088
rect 8298 4256 8354 4312
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 9126 6840 9182 6896
rect 10138 19488 10194 19544
rect 10230 19352 10286 19408
rect 9954 18572 9956 18592
rect 9956 18572 10008 18592
rect 10008 18572 10010 18592
rect 9954 18536 10010 18572
rect 9954 16904 10010 16960
rect 10046 16516 10102 16552
rect 10046 16496 10048 16516
rect 10048 16496 10100 16516
rect 10100 16496 10102 16516
rect 9586 12144 9642 12200
rect 9954 15988 9956 16008
rect 9956 15988 10008 16008
rect 10008 15988 10010 16008
rect 9954 15952 10010 15988
rect 9954 15408 10010 15464
rect 9862 13132 9864 13152
rect 9864 13132 9916 13152
rect 9916 13132 9918 13152
rect 9862 13096 9918 13132
rect 9402 11192 9458 11248
rect 9494 10804 9550 10840
rect 9494 10784 9496 10804
rect 9496 10784 9548 10804
rect 9548 10784 9550 10804
rect 9770 10784 9826 10840
rect 9494 10548 9496 10568
rect 9496 10548 9548 10568
rect 9548 10548 9550 10568
rect 9494 10512 9550 10548
rect 9402 9968 9458 10024
rect 9402 9560 9458 9616
rect 9586 9424 9642 9480
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 8850 5344 8906 5400
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 9034 4256 9090 4312
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 9126 3712 9182 3768
rect 8574 3168 8630 3224
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 9310 6568 9366 6624
rect 9310 5364 9366 5400
rect 9310 5344 9312 5364
rect 9312 5344 9364 5364
rect 9364 5344 9366 5364
rect 10230 18128 10286 18184
rect 10506 18536 10562 18592
rect 10506 16496 10562 16552
rect 10966 19116 10968 19136
rect 10968 19116 11020 19136
rect 11020 19116 11022 19136
rect 10966 19080 11022 19116
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 12622 20576 12678 20632
rect 10690 15952 10746 16008
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11794 18264 11850 18320
rect 11518 18028 11520 18048
rect 11520 18028 11572 18048
rect 11572 18028 11574 18048
rect 11518 17992 11574 18028
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 9954 12280 10010 12336
rect 9954 11328 10010 11384
rect 9770 9460 9772 9480
rect 9772 9460 9824 9480
rect 9824 9460 9826 9480
rect 9770 9424 9826 9460
rect 9770 9324 9772 9344
rect 9772 9324 9824 9344
rect 9824 9324 9826 9344
rect 9770 9288 9826 9324
rect 9678 8880 9734 8936
rect 9770 7792 9826 7848
rect 9586 6840 9642 6896
rect 9678 6740 9680 6760
rect 9680 6740 9732 6760
rect 9732 6740 9734 6760
rect 9678 6704 9734 6740
rect 9494 5208 9550 5264
rect 9310 4936 9366 4992
rect 9310 3576 9366 3632
rect 9678 4664 9734 4720
rect 9494 3576 9550 3632
rect 9218 2352 9274 2408
rect 9954 7112 10010 7168
rect 10506 13912 10562 13968
rect 10414 13776 10470 13832
rect 10506 12960 10562 13016
rect 10414 11192 10470 11248
rect 10414 10784 10470 10840
rect 10874 13132 10876 13152
rect 10876 13132 10928 13152
rect 10928 13132 10930 13152
rect 10874 13096 10930 13132
rect 10966 12960 11022 13016
rect 10782 11636 10784 11656
rect 10784 11636 10836 11656
rect 10836 11636 10838 11656
rect 10782 11600 10838 11636
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11242 14456 11298 14512
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11978 15000 12034 15056
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11702 12824 11758 12880
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11426 11736 11482 11792
rect 14278 20576 14334 20632
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 12162 17992 12218 18048
rect 12346 17584 12402 17640
rect 12438 16904 12494 16960
rect 12806 17992 12862 18048
rect 12714 17584 12770 17640
rect 13266 17856 13322 17912
rect 13174 16940 13176 16960
rect 13176 16940 13228 16960
rect 13228 16940 13230 16960
rect 13174 16904 13230 16940
rect 12438 13776 12494 13832
rect 12530 12416 12586 12472
rect 11978 11736 12034 11792
rect 11610 11328 11666 11384
rect 11610 11076 11666 11112
rect 11610 11056 11612 11076
rect 11612 11056 11664 11076
rect 11664 11056 11666 11076
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 10322 9424 10378 9480
rect 10506 8916 10508 8936
rect 10508 8916 10560 8936
rect 10560 8916 10562 8936
rect 10506 8880 10562 8916
rect 10414 7248 10470 7304
rect 10322 5888 10378 5944
rect 11150 9968 11206 10024
rect 10874 8880 10930 8936
rect 11058 8472 11114 8528
rect 10414 5616 10470 5672
rect 10322 5108 10324 5128
rect 10324 5108 10376 5128
rect 10376 5108 10378 5128
rect 10322 5072 10378 5108
rect 10322 3032 10378 3088
rect 10598 5072 10654 5128
rect 10506 3848 10562 3904
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11978 10920 12034 10976
rect 11978 10648 12034 10704
rect 12162 10648 12218 10704
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11334 7828 11336 7848
rect 11336 7828 11388 7848
rect 11388 7828 11390 7848
rect 11334 7792 11390 7828
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11702 6976 11758 7032
rect 10874 5752 10930 5808
rect 11058 5616 11114 5672
rect 10690 4120 10746 4176
rect 10598 3576 10654 3632
rect 11058 4256 11114 4312
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11334 6024 11390 6080
rect 11794 6296 11850 6352
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11426 5208 11482 5264
rect 11334 4800 11390 4856
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11334 3848 11390 3904
rect 11518 3712 11574 3768
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11886 5344 11942 5400
rect 12070 6160 12126 6216
rect 12070 5752 12126 5808
rect 11886 4936 11942 4992
rect 12070 3984 12126 4040
rect 11978 3712 12034 3768
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12622 11056 12678 11112
rect 12530 9288 12586 9344
rect 12530 8744 12586 8800
rect 12346 7792 12402 7848
rect 13818 19080 13874 19136
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13726 17992 13782 18048
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 14278 15952 14334 16008
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 14646 20304 14702 20360
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 16026 20460 16082 20496
rect 16026 20440 16028 20460
rect 16028 20440 16080 20460
rect 16080 20440 16082 20460
rect 14462 15408 14518 15464
rect 12898 9016 12954 9072
rect 12990 7112 13046 7168
rect 12530 5888 12586 5944
rect 12622 5752 12678 5808
rect 12438 5480 12494 5536
rect 12530 4936 12586 4992
rect 12622 4820 12678 4856
rect 12622 4800 12624 4820
rect 12624 4800 12676 4820
rect 12676 4800 12678 4820
rect 13358 11192 13414 11248
rect 12622 3440 12678 3496
rect 13266 9288 13322 9344
rect 13266 8744 13322 8800
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 14370 13096 14426 13152
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13542 10104 13598 10160
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13726 10512 13782 10568
rect 13634 8780 13636 8800
rect 13636 8780 13688 8800
rect 13688 8780 13690 8800
rect 13634 8744 13690 8780
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 13450 7928 13506 7984
rect 13542 7248 13598 7304
rect 13450 6024 13506 6080
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13358 4936 13414 4992
rect 13082 3168 13138 3224
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 14370 6704 14426 6760
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 13726 4528 13782 4584
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 13818 3732 13874 3768
rect 13818 3712 13820 3732
rect 13820 3712 13872 3732
rect 13872 3712 13874 3732
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 16118 17040 16174 17096
rect 14830 14456 14886 14512
rect 15014 14320 15070 14376
rect 14646 12144 14702 12200
rect 14830 10920 14886 10976
rect 14462 4120 14518 4176
rect 15014 7792 15070 7848
rect 15382 10668 15438 10704
rect 15382 10648 15384 10668
rect 15384 10648 15436 10668
rect 15436 10648 15438 10668
rect 15474 8744 15530 8800
rect 14738 5480 14794 5536
rect 15566 5616 15622 5672
rect 15750 5072 15806 5128
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 17774 17756 17776 17776
rect 17776 17756 17828 17776
rect 17828 17756 17830 17776
rect 17774 17720 17830 17756
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 18694 19896 18750 19952
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19522 18672 19578 18728
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16394 13776 16450 13832
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 17038 12688 17094 12744
rect 18050 16088 18106 16144
rect 17958 13232 18014 13288
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 20718 19372 20774 19408
rect 20718 19352 20720 19372
rect 20720 19352 20772 19372
rect 20772 19352 20774 19372
rect 21178 19760 21234 19816
rect 20994 18808 21050 18864
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 20718 17176 20774 17232
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19062 14864 19118 14920
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21270 17176 21326 17232
rect 21454 17176 21510 17232
rect 21178 16496 21234 16552
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16210 9424 16266 9480
rect 16210 9016 16266 9072
rect 16026 5344 16082 5400
rect 15842 4120 15898 4176
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16670 9560 16726 9616
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 18970 13404 18972 13424
rect 18972 13404 19024 13424
rect 19024 13404 19026 13424
rect 18970 13368 19026 13404
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 18326 12280 18382 12336
rect 17406 8880 17462 8936
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16486 6296 16542 6352
rect 16946 5616 17002 5672
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 16302 4256 16358 4312
rect 15290 3576 15346 3632
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 15934 3168 15990 3224
rect 15106 3052 15162 3088
rect 15106 3032 15108 3052
rect 15108 3032 15160 3052
rect 15160 3032 15162 3052
rect 17130 4528 17186 4584
rect 17406 5208 17462 5264
rect 17406 4664 17462 4720
rect 17866 9560 17922 9616
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19430 8492 19486 8528
rect 19430 8472 19432 8492
rect 19432 8472 19484 8492
rect 19484 8472 19486 8492
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 17406 3032 17462 3088
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 19798 11600 19854 11656
rect 19614 8472 19670 8528
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 19522 5208 19578 5264
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 19338 3052 19394 3088
rect 19338 3032 19340 3052
rect 19340 3032 19392 3052
rect 19392 3032 19394 3052
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21546 5752 21602 5808
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 21362 4120 21418 4176
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
<< metal3 >>
rect 0 21042 800 21072
rect 2221 21042 2287 21045
rect 0 21040 2287 21042
rect 0 20984 2226 21040
rect 2282 20984 2287 21040
rect 0 20982 2287 20984
rect 0 20952 800 20982
rect 2221 20979 2287 20982
rect 6144 20704 6460 20705
rect 0 20634 800 20664
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 1853 20634 1919 20637
rect 0 20632 1919 20634
rect 0 20576 1858 20632
rect 1914 20576 1919 20632
rect 0 20574 1919 20576
rect 0 20544 800 20574
rect 1853 20571 1919 20574
rect 12617 20634 12683 20637
rect 14273 20634 14339 20637
rect 12617 20632 14339 20634
rect 12617 20576 12622 20632
rect 12678 20576 14278 20632
rect 14334 20576 14339 20632
rect 12617 20574 14339 20576
rect 12617 20571 12683 20574
rect 14273 20571 14339 20574
rect 9213 20498 9279 20501
rect 16021 20498 16087 20501
rect 9213 20496 16087 20498
rect 9213 20440 9218 20496
rect 9274 20440 16026 20496
rect 16082 20440 16087 20496
rect 9213 20438 16087 20440
rect 9213 20435 9279 20438
rect 16021 20435 16087 20438
rect 7465 20362 7531 20365
rect 14641 20362 14707 20365
rect 7465 20360 14707 20362
rect 7465 20304 7470 20360
rect 7526 20304 14646 20360
rect 14702 20304 14707 20360
rect 7465 20302 14707 20304
rect 7465 20299 7531 20302
rect 14641 20299 14707 20302
rect 0 20226 800 20256
rect 1485 20226 1551 20229
rect 0 20224 1551 20226
rect 0 20168 1490 20224
rect 1546 20168 1551 20224
rect 0 20166 1551 20168
rect 0 20136 800 20166
rect 1485 20163 1551 20166
rect 3545 20160 3861 20161
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 19139 20095 19455 20096
rect 8569 19954 8635 19957
rect 18689 19954 18755 19957
rect 8569 19952 18755 19954
rect 8569 19896 8574 19952
rect 8630 19896 18694 19952
rect 18750 19896 18755 19952
rect 8569 19894 18755 19896
rect 8569 19891 8635 19894
rect 18689 19891 18755 19894
rect 0 19818 800 19848
rect 1853 19818 1919 19821
rect 0 19816 1919 19818
rect 0 19760 1858 19816
rect 1914 19760 1919 19816
rect 0 19758 1919 19760
rect 0 19728 800 19758
rect 1853 19755 1919 19758
rect 9765 19818 9831 19821
rect 21173 19818 21239 19821
rect 9765 19816 21239 19818
rect 9765 19760 9770 19816
rect 9826 19760 21178 19816
rect 21234 19760 21239 19816
rect 9765 19758 21239 19760
rect 9765 19755 9831 19758
rect 21173 19755 21239 19758
rect 2313 19682 2379 19685
rect 9581 19682 9647 19685
rect 2313 19680 5642 19682
rect 2313 19624 2318 19680
rect 2374 19624 5642 19680
rect 2313 19622 5642 19624
rect 2313 19619 2379 19622
rect 2681 19546 2747 19549
rect 4337 19546 4403 19549
rect 2681 19544 4403 19546
rect 2681 19488 2686 19544
rect 2742 19488 4342 19544
rect 4398 19488 4403 19544
rect 2681 19486 4403 19488
rect 2681 19483 2747 19486
rect 4337 19483 4403 19486
rect 0 19410 800 19440
rect 1485 19410 1551 19413
rect 0 19408 1551 19410
rect 0 19352 1490 19408
rect 1546 19352 1551 19408
rect 0 19350 1551 19352
rect 0 19320 800 19350
rect 1485 19347 1551 19350
rect 1945 19410 2011 19413
rect 4245 19410 4311 19413
rect 1945 19408 4311 19410
rect 1945 19352 1950 19408
rect 2006 19352 4250 19408
rect 4306 19352 4311 19408
rect 1945 19350 4311 19352
rect 1945 19347 2011 19350
rect 4245 19347 4311 19350
rect 4981 19410 5047 19413
rect 5390 19410 5396 19412
rect 4981 19408 5396 19410
rect 4981 19352 4986 19408
rect 5042 19352 5396 19408
rect 4981 19350 5396 19352
rect 4981 19347 5047 19350
rect 5390 19348 5396 19350
rect 5460 19348 5466 19412
rect 5582 19410 5642 19622
rect 9581 19680 10610 19682
rect 9581 19624 9586 19680
rect 9642 19624 10610 19680
rect 9581 19622 10610 19624
rect 9581 19619 9647 19622
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 9990 19484 9996 19548
rect 10060 19546 10066 19548
rect 10133 19546 10199 19549
rect 10060 19544 10199 19546
rect 10060 19488 10138 19544
rect 10194 19488 10199 19544
rect 10060 19486 10199 19488
rect 10060 19484 10066 19486
rect 10133 19483 10199 19486
rect 5717 19410 5783 19413
rect 5582 19408 5783 19410
rect 5582 19352 5722 19408
rect 5778 19352 5783 19408
rect 5582 19350 5783 19352
rect 5717 19347 5783 19350
rect 5942 19348 5948 19412
rect 6012 19410 6018 19412
rect 6545 19410 6611 19413
rect 6012 19408 6611 19410
rect 6012 19352 6550 19408
rect 6606 19352 6611 19408
rect 6012 19350 6611 19352
rect 6012 19348 6018 19350
rect 6545 19347 6611 19350
rect 7005 19410 7071 19413
rect 9213 19412 9279 19413
rect 7966 19410 7972 19412
rect 7005 19408 7972 19410
rect 7005 19352 7010 19408
rect 7066 19352 7972 19408
rect 7005 19350 7972 19352
rect 7005 19347 7071 19350
rect 7966 19348 7972 19350
rect 8036 19348 8042 19412
rect 9213 19408 9260 19412
rect 9324 19410 9330 19412
rect 10225 19410 10291 19413
rect 10358 19410 10364 19412
rect 9213 19352 9218 19408
rect 9213 19348 9260 19352
rect 9324 19350 9370 19410
rect 10225 19408 10364 19410
rect 10225 19352 10230 19408
rect 10286 19352 10364 19408
rect 10225 19350 10364 19352
rect 9324 19348 9330 19350
rect 9213 19347 9279 19348
rect 10225 19347 10291 19350
rect 10358 19348 10364 19350
rect 10428 19348 10434 19412
rect 10550 19410 10610 19622
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 21738 19551 22054 19552
rect 20713 19410 20779 19413
rect 10550 19408 20779 19410
rect 10550 19352 20718 19408
rect 20774 19352 20779 19408
rect 10550 19350 20779 19352
rect 20713 19347 20779 19350
rect 9029 19274 9095 19277
rect 11094 19274 11100 19276
rect 9029 19272 11100 19274
rect 9029 19216 9034 19272
rect 9090 19216 11100 19272
rect 9029 19214 11100 19216
rect 9029 19211 9095 19214
rect 11094 19212 11100 19214
rect 11164 19212 11170 19276
rect 9305 19138 9371 19141
rect 10961 19138 11027 19141
rect 13813 19138 13879 19141
rect 9305 19136 11027 19138
rect 9305 19080 9310 19136
rect 9366 19080 10966 19136
rect 11022 19080 11027 19136
rect 9305 19078 11027 19080
rect 9305 19075 9371 19078
rect 10961 19075 11027 19078
rect 12390 19136 13879 19138
rect 12390 19080 13818 19136
rect 13874 19080 13879 19136
rect 12390 19078 13879 19080
rect 3545 19072 3861 19073
rect 0 19002 800 19032
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 1485 19002 1551 19005
rect 12390 19002 12450 19078
rect 13813 19075 13879 19078
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 0 19000 1551 19002
rect 0 18944 1490 19000
rect 1546 18944 1551 19000
rect 0 18942 1551 18944
rect 0 18912 800 18942
rect 1485 18939 1551 18942
rect 9630 18942 12450 19002
rect 8150 18804 8156 18868
rect 8220 18866 8226 18868
rect 9630 18866 9690 18942
rect 8220 18806 9690 18866
rect 9765 18866 9831 18869
rect 20989 18866 21055 18869
rect 9765 18864 21055 18866
rect 9765 18808 9770 18864
rect 9826 18808 20994 18864
rect 21050 18808 21055 18864
rect 9765 18806 21055 18808
rect 8220 18804 8226 18806
rect 9765 18803 9831 18806
rect 20989 18803 21055 18806
rect 8477 18730 8543 18733
rect 19517 18730 19583 18733
rect 8477 18728 19583 18730
rect 8477 18672 8482 18728
rect 8538 18672 19522 18728
rect 19578 18672 19583 18728
rect 8477 18670 19583 18672
rect 8477 18667 8543 18670
rect 19517 18667 19583 18670
rect 0 18594 800 18624
rect 1485 18594 1551 18597
rect 0 18592 1551 18594
rect 0 18536 1490 18592
rect 1546 18536 1551 18592
rect 0 18534 1551 18536
rect 0 18504 800 18534
rect 1485 18531 1551 18534
rect 9397 18596 9463 18597
rect 9397 18592 9444 18596
rect 9508 18594 9514 18596
rect 9949 18594 10015 18597
rect 10501 18594 10567 18597
rect 9397 18536 9402 18592
rect 9397 18532 9444 18536
rect 9508 18534 9554 18594
rect 9949 18592 10567 18594
rect 9949 18536 9954 18592
rect 10010 18536 10506 18592
rect 10562 18536 10567 18592
rect 9949 18534 10567 18536
rect 9508 18532 9514 18534
rect 9397 18531 9463 18532
rect 9949 18531 10015 18534
rect 10501 18531 10567 18534
rect 6144 18528 6460 18529
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 21738 18463 22054 18464
rect 7598 18396 7604 18460
rect 7668 18458 7674 18460
rect 8293 18458 8359 18461
rect 7668 18456 8359 18458
rect 7668 18400 8298 18456
rect 8354 18400 8359 18456
rect 7668 18398 8359 18400
rect 7668 18396 7674 18398
rect 8293 18395 8359 18398
rect 6862 18260 6868 18324
rect 6932 18322 6938 18324
rect 11789 18322 11855 18325
rect 6932 18320 11855 18322
rect 6932 18264 11794 18320
rect 11850 18264 11855 18320
rect 6932 18262 11855 18264
rect 6932 18260 6938 18262
rect 11789 18259 11855 18262
rect 0 18186 800 18216
rect 1853 18186 1919 18189
rect 0 18184 1919 18186
rect 0 18128 1858 18184
rect 1914 18128 1919 18184
rect 0 18126 1919 18128
rect 0 18096 800 18126
rect 1853 18123 1919 18126
rect 8334 18124 8340 18188
rect 8404 18186 8410 18188
rect 10225 18186 10291 18189
rect 8404 18184 10291 18186
rect 8404 18128 10230 18184
rect 10286 18128 10291 18184
rect 8404 18126 10291 18128
rect 8404 18124 8410 18126
rect 10225 18123 10291 18126
rect 1669 18050 1735 18053
rect 9397 18052 9463 18053
rect 2446 18050 2452 18052
rect 1669 18048 2452 18050
rect 1669 17992 1674 18048
rect 1730 17992 2452 18048
rect 1669 17990 2452 17992
rect 1669 17987 1735 17990
rect 2446 17988 2452 17990
rect 2516 17988 2522 18052
rect 9397 18050 9444 18052
rect 9352 18048 9444 18050
rect 9352 17992 9402 18048
rect 9352 17990 9444 17992
rect 9397 17988 9444 17990
rect 9508 17988 9514 18052
rect 9581 18050 9647 18053
rect 11513 18050 11579 18053
rect 12157 18050 12223 18053
rect 9581 18048 12223 18050
rect 9581 17992 9586 18048
rect 9642 17992 11518 18048
rect 11574 17992 12162 18048
rect 12218 17992 12223 18048
rect 9581 17990 12223 17992
rect 9397 17987 9463 17988
rect 9581 17987 9647 17990
rect 11513 17987 11579 17990
rect 12157 17987 12223 17990
rect 12801 18050 12867 18053
rect 13721 18050 13787 18053
rect 12801 18048 13787 18050
rect 12801 17992 12806 18048
rect 12862 17992 13726 18048
rect 13782 17992 13787 18048
rect 12801 17990 13787 17992
rect 12801 17987 12867 17990
rect 13721 17987 13787 17990
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 19139 17919 19455 17920
rect 13261 17914 13327 17917
rect 9262 17912 13327 17914
rect 9262 17856 13266 17912
rect 13322 17856 13327 17912
rect 9262 17854 13327 17856
rect 0 17778 800 17808
rect 1485 17778 1551 17781
rect 0 17776 1551 17778
rect 0 17720 1490 17776
rect 1546 17720 1551 17776
rect 0 17718 1551 17720
rect 0 17688 800 17718
rect 1485 17715 1551 17718
rect 6913 17778 6979 17781
rect 9262 17778 9322 17854
rect 13261 17851 13327 17854
rect 6913 17776 9322 17778
rect 6913 17720 6918 17776
rect 6974 17720 9322 17776
rect 6913 17718 9322 17720
rect 9673 17778 9739 17781
rect 17769 17778 17835 17781
rect 9673 17776 17835 17778
rect 9673 17720 9678 17776
rect 9734 17720 17774 17776
rect 17830 17720 17835 17776
rect 9673 17718 17835 17720
rect 6913 17715 6979 17718
rect 9673 17715 9739 17718
rect 17769 17715 17835 17718
rect 5165 17642 5231 17645
rect 9581 17642 9647 17645
rect 5165 17640 9647 17642
rect 5165 17584 5170 17640
rect 5226 17584 9586 17640
rect 9642 17584 9647 17640
rect 5165 17582 9647 17584
rect 5165 17579 5231 17582
rect 9581 17579 9647 17582
rect 12341 17642 12407 17645
rect 12709 17642 12775 17645
rect 12341 17640 12775 17642
rect 12341 17584 12346 17640
rect 12402 17584 12714 17640
rect 12770 17584 12775 17640
rect 12341 17582 12775 17584
rect 12341 17579 12407 17582
rect 12709 17579 12775 17582
rect 6144 17440 6460 17441
rect 0 17370 800 17400
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 1485 17370 1551 17373
rect 0 17368 1551 17370
rect 0 17312 1490 17368
rect 1546 17312 1551 17368
rect 0 17310 1551 17312
rect 0 17280 800 17310
rect 1485 17307 1551 17310
rect 7741 17234 7807 17237
rect 20713 17234 20779 17237
rect 21265 17234 21331 17237
rect 7741 17232 21331 17234
rect 7741 17176 7746 17232
rect 7802 17176 20718 17232
rect 20774 17176 21270 17232
rect 21326 17176 21331 17232
rect 7741 17174 21331 17176
rect 7741 17171 7807 17174
rect 20713 17171 20779 17174
rect 21265 17171 21331 17174
rect 21449 17234 21515 17237
rect 22200 17234 23000 17264
rect 21449 17232 23000 17234
rect 21449 17176 21454 17232
rect 21510 17176 23000 17232
rect 21449 17174 23000 17176
rect 21449 17171 21515 17174
rect 22200 17144 23000 17174
rect 6177 17098 6243 17101
rect 16113 17098 16179 17101
rect 6177 17096 16179 17098
rect 6177 17040 6182 17096
rect 6238 17040 16118 17096
rect 16174 17040 16179 17096
rect 6177 17038 16179 17040
rect 6177 17035 6243 17038
rect 16113 17035 16179 17038
rect 0 16962 800 16992
rect 1485 16962 1551 16965
rect 0 16960 1551 16962
rect 0 16904 1490 16960
rect 1546 16904 1551 16960
rect 0 16902 1551 16904
rect 0 16872 800 16902
rect 1485 16899 1551 16902
rect 9806 16900 9812 16964
rect 9876 16962 9882 16964
rect 9949 16962 10015 16965
rect 9876 16960 10015 16962
rect 9876 16904 9954 16960
rect 10010 16904 10015 16960
rect 9876 16902 10015 16904
rect 9876 16900 9882 16902
rect 9949 16899 10015 16902
rect 12433 16962 12499 16965
rect 13169 16962 13235 16965
rect 12433 16960 13235 16962
rect 12433 16904 12438 16960
rect 12494 16904 13174 16960
rect 13230 16904 13235 16960
rect 12433 16902 13235 16904
rect 12433 16899 12499 16902
rect 13169 16899 13235 16902
rect 3545 16896 3861 16897
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 19139 16831 19455 16832
rect 0 16554 800 16584
rect 1853 16554 1919 16557
rect 0 16552 1919 16554
rect 0 16496 1858 16552
rect 1914 16496 1919 16552
rect 0 16494 1919 16496
rect 0 16464 800 16494
rect 1853 16491 1919 16494
rect 4153 16554 4219 16557
rect 10041 16554 10107 16557
rect 4153 16552 10107 16554
rect 4153 16496 4158 16552
rect 4214 16496 10046 16552
rect 10102 16496 10107 16552
rect 4153 16494 10107 16496
rect 4153 16491 4219 16494
rect 10041 16491 10107 16494
rect 10501 16554 10567 16557
rect 21173 16554 21239 16557
rect 10501 16552 21239 16554
rect 10501 16496 10506 16552
rect 10562 16496 21178 16552
rect 21234 16496 21239 16552
rect 10501 16494 21239 16496
rect 10501 16491 10567 16494
rect 21173 16491 21239 16494
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 21738 16287 22054 16288
rect 6729 16282 6795 16285
rect 6862 16282 6868 16284
rect 6729 16280 6868 16282
rect 6729 16224 6734 16280
rect 6790 16224 6868 16280
rect 6729 16222 6868 16224
rect 6729 16219 6795 16222
rect 6862 16220 6868 16222
rect 6932 16220 6938 16284
rect 7782 16220 7788 16284
rect 7852 16282 7858 16284
rect 8201 16282 8267 16285
rect 8385 16282 8451 16285
rect 7852 16280 8451 16282
rect 7852 16224 8206 16280
rect 8262 16224 8390 16280
rect 8446 16224 8451 16280
rect 7852 16222 8451 16224
rect 7852 16220 7858 16222
rect 8201 16219 8267 16222
rect 8385 16219 8451 16222
rect 0 16146 800 16176
rect 1485 16146 1551 16149
rect 0 16144 1551 16146
rect 0 16088 1490 16144
rect 1546 16088 1551 16144
rect 0 16086 1551 16088
rect 0 16056 800 16086
rect 1485 16083 1551 16086
rect 5257 16146 5323 16149
rect 5901 16146 5967 16149
rect 5257 16144 5967 16146
rect 5257 16088 5262 16144
rect 5318 16088 5906 16144
rect 5962 16088 5967 16144
rect 5257 16086 5967 16088
rect 5257 16083 5323 16086
rect 5901 16083 5967 16086
rect 6913 16146 6979 16149
rect 18045 16146 18111 16149
rect 6913 16144 18111 16146
rect 6913 16088 6918 16144
rect 6974 16088 18050 16144
rect 18106 16088 18111 16144
rect 6913 16086 18111 16088
rect 6913 16083 6979 16086
rect 18045 16083 18111 16086
rect 7741 16010 7807 16013
rect 9397 16012 9463 16013
rect 7741 16008 9322 16010
rect 7741 15952 7746 16008
rect 7802 15952 9322 16008
rect 7741 15950 9322 15952
rect 7741 15947 7807 15950
rect 5758 15812 5764 15876
rect 5828 15874 5834 15876
rect 6361 15874 6427 15877
rect 5828 15872 6427 15874
rect 5828 15816 6366 15872
rect 6422 15816 6427 15872
rect 5828 15814 6427 15816
rect 9262 15874 9322 15950
rect 9397 16008 9444 16012
rect 9508 16010 9514 16012
rect 9949 16010 10015 16013
rect 9508 16008 10015 16010
rect 9397 15952 9402 16008
rect 9508 15952 9954 16008
rect 10010 15952 10015 16008
rect 9397 15948 9444 15952
rect 9508 15950 10015 15952
rect 9508 15948 9514 15950
rect 9397 15947 9463 15948
rect 9949 15947 10015 15950
rect 10685 16010 10751 16013
rect 11830 16010 11836 16012
rect 10685 16008 11836 16010
rect 10685 15952 10690 16008
rect 10746 15952 11836 16008
rect 10685 15950 11836 15952
rect 10685 15947 10751 15950
rect 11830 15948 11836 15950
rect 11900 15948 11906 16012
rect 14273 16010 14339 16013
rect 12390 16008 14339 16010
rect 12390 15952 14278 16008
rect 14334 15952 14339 16008
rect 12390 15950 14339 15952
rect 12390 15874 12450 15950
rect 14273 15947 14339 15950
rect 9262 15814 12450 15874
rect 5828 15812 5834 15814
rect 6361 15811 6427 15814
rect 3545 15808 3861 15809
rect 0 15738 800 15768
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 1485 15738 1551 15741
rect 0 15736 1551 15738
rect 0 15680 1490 15736
rect 1546 15680 1551 15736
rect 0 15678 1551 15680
rect 0 15648 800 15678
rect 1485 15675 1551 15678
rect 5073 15602 5139 15605
rect 5073 15600 8448 15602
rect 5073 15544 5078 15600
rect 5134 15544 8448 15600
rect 5073 15542 8448 15544
rect 5073 15539 5139 15542
rect 8388 15466 8448 15542
rect 8518 15540 8524 15604
rect 8588 15602 8594 15604
rect 9397 15602 9463 15605
rect 8588 15600 9463 15602
rect 8588 15544 9402 15600
rect 9458 15544 9463 15600
rect 8588 15542 9463 15544
rect 8588 15540 8594 15542
rect 9397 15539 9463 15542
rect 9397 15466 9463 15469
rect 8388 15464 9463 15466
rect 8388 15408 9402 15464
rect 9458 15408 9463 15464
rect 8388 15406 9463 15408
rect 9397 15403 9463 15406
rect 9949 15466 10015 15469
rect 14457 15466 14523 15469
rect 9949 15464 14523 15466
rect 9949 15408 9954 15464
rect 10010 15408 14462 15464
rect 14518 15408 14523 15464
rect 9949 15406 14523 15408
rect 9949 15403 10015 15406
rect 14457 15403 14523 15406
rect 0 15330 800 15360
rect 1485 15330 1551 15333
rect 0 15328 1551 15330
rect 0 15272 1490 15328
rect 1546 15272 1551 15328
rect 0 15270 1551 15272
rect 0 15240 800 15270
rect 1485 15267 1551 15270
rect 6144 15264 6460 15265
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 21738 15199 22054 15200
rect 8109 15194 8175 15197
rect 8293 15194 8359 15197
rect 9029 15194 9095 15197
rect 8109 15192 9095 15194
rect 8109 15136 8114 15192
rect 8170 15136 8298 15192
rect 8354 15136 9034 15192
rect 9090 15136 9095 15192
rect 8109 15134 9095 15136
rect 8109 15131 8175 15134
rect 8293 15131 8359 15134
rect 9029 15131 9095 15134
rect 8109 15060 8175 15061
rect 8109 15058 8156 15060
rect 8064 15056 8156 15058
rect 8064 15000 8114 15056
rect 8064 14998 8156 15000
rect 8109 14996 8156 14998
rect 8220 14996 8226 15060
rect 11973 15058 12039 15061
rect 8572 15056 12039 15058
rect 8572 15000 11978 15056
rect 12034 15000 12039 15056
rect 8572 14998 12039 15000
rect 8109 14995 8175 14996
rect 0 14922 800 14952
rect 1853 14922 1919 14925
rect 0 14920 1919 14922
rect 0 14864 1858 14920
rect 1914 14864 1919 14920
rect 0 14862 1919 14864
rect 0 14832 800 14862
rect 1853 14859 1919 14862
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 4613 14650 4679 14653
rect 8572 14650 8632 14998
rect 11973 14995 12039 14998
rect 9305 14922 9371 14925
rect 19057 14922 19123 14925
rect 9305 14920 19123 14922
rect 9305 14864 9310 14920
rect 9366 14864 19062 14920
rect 19118 14864 19123 14920
rect 9305 14862 19123 14864
rect 9305 14859 9371 14862
rect 19057 14859 19123 14862
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 19139 14655 19455 14656
rect 4613 14648 8632 14650
rect 4613 14592 4618 14648
rect 4674 14592 8632 14648
rect 4613 14590 8632 14592
rect 4613 14587 4679 14590
rect 0 14514 800 14544
rect 1485 14514 1551 14517
rect 0 14512 1551 14514
rect 0 14456 1490 14512
rect 1546 14456 1551 14512
rect 0 14454 1551 14456
rect 0 14424 800 14454
rect 1485 14451 1551 14454
rect 6269 14514 6335 14517
rect 8150 14514 8156 14516
rect 6269 14512 8156 14514
rect 6269 14456 6274 14512
rect 6330 14456 8156 14512
rect 6269 14454 8156 14456
rect 6269 14451 6335 14454
rect 8150 14452 8156 14454
rect 8220 14514 8226 14516
rect 8753 14514 8819 14517
rect 8220 14512 8819 14514
rect 8220 14456 8758 14512
rect 8814 14456 8819 14512
rect 8220 14454 8819 14456
rect 8220 14452 8226 14454
rect 8753 14451 8819 14454
rect 11237 14514 11303 14517
rect 14825 14514 14891 14517
rect 11237 14512 14891 14514
rect 11237 14456 11242 14512
rect 11298 14456 14830 14512
rect 14886 14456 14891 14512
rect 11237 14454 14891 14456
rect 11237 14451 11303 14454
rect 14825 14451 14891 14454
rect 5073 14378 5139 14381
rect 5206 14378 5212 14380
rect 5073 14376 5212 14378
rect 5073 14320 5078 14376
rect 5134 14320 5212 14376
rect 5073 14318 5212 14320
rect 5073 14315 5139 14318
rect 5206 14316 5212 14318
rect 5276 14378 5282 14380
rect 15009 14378 15075 14381
rect 5276 14376 15075 14378
rect 5276 14320 15014 14376
rect 15070 14320 15075 14376
rect 5276 14318 15075 14320
rect 5276 14316 5282 14318
rect 15009 14315 15075 14318
rect 6144 14176 6460 14177
rect 0 14106 800 14136
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 1485 14106 1551 14109
rect 0 14104 1551 14106
rect 0 14048 1490 14104
rect 1546 14048 1551 14104
rect 0 14046 1551 14048
rect 0 14016 800 14046
rect 1485 14043 1551 14046
rect 6453 13970 6519 13973
rect 10501 13970 10567 13973
rect 6453 13968 10567 13970
rect 6453 13912 6458 13968
rect 6514 13912 10506 13968
rect 10562 13912 10567 13968
rect 6453 13910 10567 13912
rect 6453 13907 6519 13910
rect 10501 13907 10567 13910
rect 10409 13834 10475 13837
rect 8572 13832 10475 13834
rect 8572 13776 10414 13832
rect 10470 13776 10475 13832
rect 8572 13774 10475 13776
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 6862 13636 6868 13700
rect 6932 13698 6938 13700
rect 8572 13698 8632 13774
rect 10409 13771 10475 13774
rect 12433 13834 12499 13837
rect 16389 13834 16455 13837
rect 12433 13832 16455 13834
rect 12433 13776 12438 13832
rect 12494 13776 16394 13832
rect 16450 13776 16455 13832
rect 12433 13774 16455 13776
rect 12433 13771 12499 13774
rect 16389 13771 16455 13774
rect 6932 13638 8632 13698
rect 6932 13636 6938 13638
rect 3545 13632 3861 13633
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 19139 13567 19455 13568
rect 5390 13500 5396 13564
rect 5460 13562 5466 13564
rect 6177 13562 6243 13565
rect 6729 13562 6795 13565
rect 5460 13560 6795 13562
rect 5460 13504 6182 13560
rect 6238 13504 6734 13560
rect 6790 13504 6795 13560
rect 5460 13502 6795 13504
rect 5460 13500 5466 13502
rect 6177 13499 6243 13502
rect 6729 13499 6795 13502
rect 8661 13426 8727 13429
rect 18965 13426 19031 13429
rect 8661 13424 19031 13426
rect 8661 13368 8666 13424
rect 8722 13368 18970 13424
rect 19026 13368 19031 13424
rect 8661 13366 19031 13368
rect 8661 13363 8727 13366
rect 18965 13363 19031 13366
rect 0 13290 800 13320
rect 1485 13290 1551 13293
rect 0 13288 1551 13290
rect 0 13232 1490 13288
rect 1546 13232 1551 13288
rect 0 13230 1551 13232
rect 0 13200 800 13230
rect 1485 13227 1551 13230
rect 5257 13290 5323 13293
rect 17953 13290 18019 13293
rect 5257 13288 18019 13290
rect 5257 13232 5262 13288
rect 5318 13232 17958 13288
rect 18014 13232 18019 13288
rect 5257 13230 18019 13232
rect 5257 13227 5323 13230
rect 17953 13227 18019 13230
rect 9857 13154 9923 13157
rect 10869 13154 10935 13157
rect 9857 13152 10935 13154
rect 9857 13096 9862 13152
rect 9918 13096 10874 13152
rect 10930 13096 10935 13152
rect 9857 13094 10935 13096
rect 9857 13091 9923 13094
rect 10869 13091 10935 13094
rect 14365 13154 14431 13157
rect 14365 13152 14474 13154
rect 14365 13096 14370 13152
rect 14426 13096 14474 13152
rect 14365 13091 14474 13096
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 6545 13018 6611 13021
rect 7649 13018 7715 13021
rect 6545 13016 7715 13018
rect 6545 12960 6550 13016
rect 6606 12960 7654 13016
rect 7710 12960 7715 13016
rect 6545 12958 7715 12960
rect 6545 12955 6611 12958
rect 7649 12955 7715 12958
rect 10501 13018 10567 13021
rect 10961 13018 11027 13021
rect 10501 13016 11027 13018
rect 10501 12960 10506 13016
rect 10562 12960 10966 13016
rect 11022 12960 11027 13016
rect 10501 12958 11027 12960
rect 10501 12955 10567 12958
rect 10961 12955 11027 12958
rect 0 12882 800 12912
rect 1393 12882 1459 12885
rect 0 12880 1459 12882
rect 0 12824 1398 12880
rect 1454 12824 1459 12880
rect 0 12822 1459 12824
rect 0 12792 800 12822
rect 1393 12819 1459 12822
rect 3969 12882 4035 12885
rect 11697 12882 11763 12885
rect 3969 12880 11763 12882
rect 3969 12824 3974 12880
rect 4030 12824 11702 12880
rect 11758 12824 11763 12880
rect 3969 12822 11763 12824
rect 3969 12819 4035 12822
rect 11697 12819 11763 12822
rect 7373 12746 7439 12749
rect 14414 12746 14474 13091
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 21738 13023 22054 13024
rect 17033 12746 17099 12749
rect 7373 12744 17099 12746
rect 7373 12688 7378 12744
rect 7434 12688 17038 12744
rect 17094 12688 17099 12744
rect 7373 12686 17099 12688
rect 7373 12683 7439 12686
rect 17033 12683 17099 12686
rect 6821 12612 6887 12613
rect 6821 12608 6868 12612
rect 6932 12610 6938 12612
rect 6821 12552 6826 12608
rect 6821 12548 6868 12552
rect 6932 12550 6978 12610
rect 6932 12548 6938 12550
rect 6821 12547 6887 12548
rect 3545 12544 3861 12545
rect 0 12474 800 12504
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 1669 12474 1735 12477
rect 0 12472 1735 12474
rect 0 12416 1674 12472
rect 1730 12416 1735 12472
rect 0 12414 1735 12416
rect 0 12384 800 12414
rect 1669 12411 1735 12414
rect 6678 12412 6684 12476
rect 6748 12474 6754 12476
rect 12525 12474 12591 12477
rect 6748 12414 8632 12474
rect 6748 12412 6754 12414
rect 6545 12338 6611 12341
rect 6502 12336 6611 12338
rect 6502 12280 6550 12336
rect 6606 12280 6611 12336
rect 6502 12275 6611 12280
rect 8572 12338 8632 12414
rect 9262 12472 12591 12474
rect 9262 12416 12530 12472
rect 12586 12416 12591 12472
rect 9262 12414 12591 12416
rect 9262 12338 9322 12414
rect 12525 12411 12591 12414
rect 8572 12278 9322 12338
rect 9949 12338 10015 12341
rect 18321 12338 18387 12341
rect 9949 12336 18387 12338
rect 9949 12280 9954 12336
rect 10010 12280 18326 12336
rect 18382 12280 18387 12336
rect 9949 12278 18387 12280
rect 9949 12275 10015 12278
rect 18321 12275 18387 12278
rect 6502 12202 6562 12275
rect 9581 12202 9647 12205
rect 14641 12202 14707 12205
rect 6502 12142 9322 12202
rect 0 12066 800 12096
rect 1393 12066 1459 12069
rect 6729 12068 6795 12069
rect 0 12064 1459 12066
rect 0 12008 1398 12064
rect 1454 12008 1459 12064
rect 0 12006 1459 12008
rect 0 11976 800 12006
rect 1393 12003 1459 12006
rect 6678 12004 6684 12068
rect 6748 12066 6795 12068
rect 9262 12066 9322 12142
rect 9581 12200 14707 12202
rect 9581 12144 9586 12200
rect 9642 12144 14646 12200
rect 14702 12144 14707 12200
rect 9581 12142 14707 12144
rect 9581 12139 9647 12142
rect 14641 12139 14707 12142
rect 10910 12066 10916 12068
rect 6748 12064 6840 12066
rect 6790 12008 6840 12064
rect 6748 12006 6840 12008
rect 9262 12006 10916 12066
rect 6748 12004 6795 12006
rect 10910 12004 10916 12006
rect 10980 12004 10986 12068
rect 6729 12003 6795 12004
rect 6144 12000 6460 12001
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 21738 11935 22054 11936
rect 7925 11930 7991 11933
rect 8150 11930 8156 11932
rect 7925 11928 8156 11930
rect 7925 11872 7930 11928
rect 7986 11872 8156 11928
rect 7925 11870 8156 11872
rect 7925 11867 7991 11870
rect 8150 11868 8156 11870
rect 8220 11868 8226 11932
rect 11421 11794 11487 11797
rect 11830 11794 11836 11796
rect 11421 11792 11836 11794
rect 11421 11736 11426 11792
rect 11482 11736 11836 11792
rect 11421 11734 11836 11736
rect 11421 11731 11487 11734
rect 11830 11732 11836 11734
rect 11900 11794 11906 11796
rect 11973 11794 12039 11797
rect 11900 11792 12039 11794
rect 11900 11736 11978 11792
rect 12034 11736 12039 11792
rect 11900 11734 12039 11736
rect 11900 11732 11906 11734
rect 11973 11731 12039 11734
rect 0 11658 800 11688
rect 1393 11658 1459 11661
rect 0 11656 1459 11658
rect 0 11600 1398 11656
rect 1454 11600 1459 11656
rect 0 11598 1459 11600
rect 0 11568 800 11598
rect 1393 11595 1459 11598
rect 10777 11658 10843 11661
rect 19793 11658 19859 11661
rect 10777 11656 19859 11658
rect 10777 11600 10782 11656
rect 10838 11600 19798 11656
rect 19854 11600 19859 11656
rect 10777 11598 19859 11600
rect 10777 11595 10843 11598
rect 19793 11595 19859 11598
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 19139 11391 19455 11392
rect 9949 11388 10015 11389
rect 9949 11386 9996 11388
rect 9904 11384 9996 11386
rect 9904 11328 9954 11384
rect 9904 11326 9996 11328
rect 9949 11324 9996 11326
rect 10060 11324 10066 11388
rect 11605 11386 11671 11389
rect 12198 11386 12204 11388
rect 11605 11384 12204 11386
rect 11605 11328 11610 11384
rect 11666 11328 12204 11384
rect 11605 11326 12204 11328
rect 9949 11323 10015 11324
rect 11605 11323 11671 11326
rect 12198 11324 12204 11326
rect 12268 11324 12274 11388
rect 0 11250 800 11280
rect 1669 11250 1735 11253
rect 0 11248 1735 11250
rect 0 11192 1674 11248
rect 1730 11192 1735 11248
rect 0 11190 1735 11192
rect 0 11160 800 11190
rect 1669 11187 1735 11190
rect 5717 11252 5783 11253
rect 5717 11248 5764 11252
rect 5828 11250 5834 11252
rect 7189 11250 7255 11253
rect 9397 11250 9463 11253
rect 5717 11192 5722 11248
rect 5717 11188 5764 11192
rect 5828 11190 5874 11250
rect 7189 11248 9463 11250
rect 7189 11192 7194 11248
rect 7250 11192 9402 11248
rect 9458 11192 9463 11248
rect 7189 11190 9463 11192
rect 5828 11188 5834 11190
rect 5717 11187 5783 11188
rect 7189 11187 7255 11190
rect 9397 11187 9463 11190
rect 10409 11250 10475 11253
rect 13353 11250 13419 11253
rect 10409 11248 13419 11250
rect 10409 11192 10414 11248
rect 10470 11192 13358 11248
rect 13414 11192 13419 11248
rect 10409 11190 13419 11192
rect 10409 11187 10475 11190
rect 13353 11187 13419 11190
rect 11605 11114 11671 11117
rect 12617 11114 12683 11117
rect 11605 11112 12683 11114
rect 11605 11056 11610 11112
rect 11666 11056 12622 11112
rect 12678 11056 12683 11112
rect 11605 11054 12683 11056
rect 11605 11051 11671 11054
rect 12617 11051 12683 11054
rect 11973 10978 12039 10981
rect 14825 10978 14891 10981
rect 11973 10976 14891 10978
rect 11973 10920 11978 10976
rect 12034 10920 14830 10976
rect 14886 10920 14891 10976
rect 11973 10918 14891 10920
rect 11973 10915 12039 10918
rect 14825 10915 14891 10918
rect 6144 10912 6460 10913
rect 0 10842 800 10872
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 1393 10842 1459 10845
rect 0 10840 1459 10842
rect 0 10784 1398 10840
rect 1454 10784 1459 10840
rect 0 10782 1459 10784
rect 0 10752 800 10782
rect 1393 10779 1459 10782
rect 7598 10780 7604 10844
rect 7668 10842 7674 10844
rect 9489 10842 9555 10845
rect 7668 10840 9555 10842
rect 7668 10784 9494 10840
rect 9550 10784 9555 10840
rect 7668 10782 9555 10784
rect 7668 10780 7674 10782
rect 9489 10779 9555 10782
rect 9765 10842 9831 10845
rect 10409 10844 10475 10845
rect 10358 10842 10364 10844
rect 9765 10840 10364 10842
rect 10428 10842 10475 10844
rect 10428 10840 10556 10842
rect 9765 10784 9770 10840
rect 9826 10784 10364 10840
rect 10470 10784 10556 10840
rect 9765 10782 10364 10784
rect 9765 10779 9831 10782
rect 10358 10780 10364 10782
rect 10428 10782 10556 10784
rect 10428 10780 10475 10782
rect 10409 10779 10475 10780
rect 6637 10706 6703 10709
rect 11973 10706 12039 10709
rect 6637 10704 12039 10706
rect 6637 10648 6642 10704
rect 6698 10648 11978 10704
rect 12034 10648 12039 10704
rect 6637 10646 12039 10648
rect 6637 10643 6703 10646
rect 11973 10643 12039 10646
rect 12157 10706 12223 10709
rect 15377 10706 15443 10709
rect 12157 10704 15443 10706
rect 12157 10648 12162 10704
rect 12218 10648 15382 10704
rect 15438 10648 15443 10704
rect 12157 10646 15443 10648
rect 12157 10643 12223 10646
rect 15377 10643 15443 10646
rect 7598 10508 7604 10572
rect 7668 10570 7674 10572
rect 7925 10570 7991 10573
rect 7668 10568 7991 10570
rect 7668 10512 7930 10568
rect 7986 10512 7991 10568
rect 7668 10510 7991 10512
rect 7668 10508 7674 10510
rect 7925 10507 7991 10510
rect 8518 10508 8524 10572
rect 8588 10570 8594 10572
rect 9121 10570 9187 10573
rect 8588 10568 9187 10570
rect 8588 10512 9126 10568
rect 9182 10512 9187 10568
rect 8588 10510 9187 10512
rect 8588 10508 8594 10510
rect 9121 10507 9187 10510
rect 9489 10570 9555 10573
rect 13721 10570 13787 10573
rect 9489 10568 13787 10570
rect 9489 10512 9494 10568
rect 9550 10512 13726 10568
rect 13782 10512 13787 10568
rect 9489 10510 13787 10512
rect 9489 10507 9555 10510
rect 13721 10507 13787 10510
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 4705 10434 4771 10437
rect 7281 10434 7347 10437
rect 4705 10432 7347 10434
rect 4705 10376 4710 10432
rect 4766 10376 7286 10432
rect 7342 10376 7347 10432
rect 4705 10374 7347 10376
rect 4705 10371 4771 10374
rect 7281 10371 7347 10374
rect 3545 10368 3861 10369
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 19139 10303 19455 10304
rect 5206 10236 5212 10300
rect 5276 10298 5282 10300
rect 7005 10298 7071 10301
rect 5276 10296 7071 10298
rect 5276 10240 7010 10296
rect 7066 10240 7071 10296
rect 5276 10238 7071 10240
rect 5276 10236 5282 10238
rect 7005 10235 7071 10238
rect 2865 10162 2931 10165
rect 3141 10162 3207 10165
rect 3785 10162 3851 10165
rect 4705 10162 4771 10165
rect 2865 10160 4771 10162
rect 2865 10104 2870 10160
rect 2926 10104 3146 10160
rect 3202 10104 3790 10160
rect 3846 10104 4710 10160
rect 4766 10104 4771 10160
rect 2865 10102 4771 10104
rect 2865 10099 2931 10102
rect 3141 10099 3207 10102
rect 3785 10099 3851 10102
rect 4705 10099 4771 10102
rect 6085 10162 6151 10165
rect 7782 10162 7788 10164
rect 6085 10160 7788 10162
rect 6085 10104 6090 10160
rect 6146 10104 7788 10160
rect 6085 10102 7788 10104
rect 6085 10099 6151 10102
rect 7782 10100 7788 10102
rect 7852 10100 7858 10164
rect 8293 10162 8359 10165
rect 13537 10162 13603 10165
rect 8293 10160 13603 10162
rect 8293 10104 8298 10160
rect 8354 10104 13542 10160
rect 13598 10104 13603 10160
rect 8293 10102 13603 10104
rect 8293 10099 8359 10102
rect 13537 10099 13603 10102
rect 0 10026 800 10056
rect 1393 10026 1459 10029
rect 0 10024 1459 10026
rect 0 9968 1398 10024
rect 1454 9968 1459 10024
rect 0 9966 1459 9968
rect 0 9936 800 9966
rect 1393 9963 1459 9966
rect 1577 10026 1643 10029
rect 9397 10026 9463 10029
rect 11145 10026 11211 10029
rect 1577 10024 11211 10026
rect 1577 9968 1582 10024
rect 1638 9968 9402 10024
rect 9458 9968 11150 10024
rect 11206 9968 11211 10024
rect 1577 9966 11211 9968
rect 1577 9963 1643 9966
rect 9397 9963 9463 9966
rect 11145 9963 11211 9966
rect 5390 9828 5396 9892
rect 5460 9890 5466 9892
rect 5625 9890 5691 9893
rect 5460 9888 5691 9890
rect 5460 9832 5630 9888
rect 5686 9832 5691 9888
rect 5460 9830 5691 9832
rect 5460 9828 5466 9830
rect 5625 9827 5691 9830
rect 8334 9828 8340 9892
rect 8404 9890 8410 9892
rect 8477 9890 8543 9893
rect 8404 9888 8543 9890
rect 8404 9832 8482 9888
rect 8538 9832 8543 9888
rect 8404 9830 8543 9832
rect 8404 9828 8410 9830
rect 8477 9827 8543 9830
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 21738 9759 22054 9760
rect 0 9618 800 9648
rect 1669 9618 1735 9621
rect 0 9616 1735 9618
rect 0 9560 1674 9616
rect 1730 9560 1735 9616
rect 0 9558 1735 9560
rect 0 9528 800 9558
rect 1669 9555 1735 9558
rect 5901 9618 5967 9621
rect 8661 9618 8727 9621
rect 5901 9616 8727 9618
rect 5901 9560 5906 9616
rect 5962 9560 8666 9616
rect 8722 9560 8727 9616
rect 5901 9558 8727 9560
rect 5901 9555 5967 9558
rect 8661 9555 8727 9558
rect 9397 9618 9463 9621
rect 16665 9618 16731 9621
rect 17861 9618 17927 9621
rect 9397 9616 17927 9618
rect 9397 9560 9402 9616
rect 9458 9560 16670 9616
rect 16726 9560 17866 9616
rect 17922 9560 17927 9616
rect 9397 9558 17927 9560
rect 9397 9555 9463 9558
rect 16665 9555 16731 9558
rect 17861 9555 17927 9558
rect 2405 9484 2471 9485
rect 2405 9482 2452 9484
rect 2360 9480 2452 9482
rect 2360 9424 2410 9480
rect 2360 9422 2452 9424
rect 2405 9420 2452 9422
rect 2516 9420 2522 9484
rect 4981 9482 5047 9485
rect 9581 9482 9647 9485
rect 4981 9480 9647 9482
rect 4981 9424 4986 9480
rect 5042 9424 9586 9480
rect 9642 9424 9647 9480
rect 4981 9422 9647 9424
rect 2405 9419 2471 9420
rect 4981 9419 5047 9422
rect 9581 9419 9647 9422
rect 9765 9484 9831 9485
rect 9765 9480 9812 9484
rect 9876 9482 9882 9484
rect 10317 9482 10383 9485
rect 16205 9482 16271 9485
rect 9765 9424 9770 9480
rect 9765 9420 9812 9424
rect 9876 9422 9922 9482
rect 10317 9480 16271 9482
rect 10317 9424 10322 9480
rect 10378 9424 16210 9480
rect 16266 9424 16271 9480
rect 10317 9422 16271 9424
rect 9876 9420 9882 9422
rect 9765 9419 9831 9420
rect 10317 9419 10383 9422
rect 16205 9419 16271 9422
rect 5993 9346 6059 9349
rect 8477 9348 8543 9349
rect 9765 9348 9831 9349
rect 8477 9346 8524 9348
rect 5993 9344 8524 9346
rect 5993 9288 5998 9344
rect 6054 9288 8482 9344
rect 5993 9286 8524 9288
rect 5993 9283 6059 9286
rect 8477 9284 8524 9286
rect 8588 9284 8594 9348
rect 9765 9346 9812 9348
rect 9720 9344 9812 9346
rect 9720 9288 9770 9344
rect 9720 9286 9812 9288
rect 9765 9284 9812 9286
rect 9876 9284 9882 9348
rect 12525 9346 12591 9349
rect 13261 9346 13327 9349
rect 12525 9344 13327 9346
rect 12525 9288 12530 9344
rect 12586 9288 13266 9344
rect 13322 9288 13327 9344
rect 12525 9286 13327 9288
rect 8477 9283 8543 9284
rect 9765 9283 9831 9284
rect 12525 9283 12591 9286
rect 13261 9283 13327 9286
rect 3545 9280 3861 9281
rect 0 9210 800 9240
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 1393 9210 1459 9213
rect 0 9208 1459 9210
rect 0 9152 1398 9208
rect 1454 9152 1459 9208
rect 0 9150 1459 9152
rect 0 9120 800 9150
rect 1393 9147 1459 9150
rect 6821 9074 6887 9077
rect 12893 9074 12959 9077
rect 6821 9072 12959 9074
rect 6821 9016 6826 9072
rect 6882 9016 12898 9072
rect 12954 9016 12959 9072
rect 6821 9014 12959 9016
rect 13264 9074 13324 9283
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 16205 9074 16271 9077
rect 13264 9072 16271 9074
rect 13264 9016 16210 9072
rect 16266 9016 16271 9072
rect 13264 9014 16271 9016
rect 6821 9011 6887 9014
rect 12893 9011 12959 9014
rect 16205 9011 16271 9014
rect 8661 8938 8727 8941
rect 9673 8938 9739 8941
rect 10501 8938 10567 8941
rect 8661 8936 10567 8938
rect 8661 8880 8666 8936
rect 8722 8880 9678 8936
rect 9734 8880 10506 8936
rect 10562 8880 10567 8936
rect 8661 8878 10567 8880
rect 8661 8875 8727 8878
rect 9673 8875 9739 8878
rect 10501 8875 10567 8878
rect 10869 8938 10935 8941
rect 17401 8938 17467 8941
rect 10869 8936 17467 8938
rect 10869 8880 10874 8936
rect 10930 8880 17406 8936
rect 17462 8880 17467 8936
rect 10869 8878 17467 8880
rect 10869 8875 10935 8878
rect 17401 8875 17467 8878
rect 0 8802 800 8832
rect 1669 8802 1735 8805
rect 0 8800 1735 8802
rect 0 8744 1674 8800
rect 1730 8744 1735 8800
rect 0 8742 1735 8744
rect 0 8712 800 8742
rect 1669 8739 1735 8742
rect 12525 8802 12591 8805
rect 13261 8802 13327 8805
rect 13629 8802 13695 8805
rect 15469 8802 15535 8805
rect 12525 8800 15535 8802
rect 12525 8744 12530 8800
rect 12586 8744 13266 8800
rect 13322 8744 13634 8800
rect 13690 8744 15474 8800
rect 15530 8744 15535 8800
rect 12525 8742 15535 8744
rect 12525 8739 12591 8742
rect 13261 8739 13327 8742
rect 13629 8739 13695 8742
rect 15469 8739 15535 8742
rect 6144 8736 6460 8737
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 21738 8671 22054 8672
rect 3233 8530 3299 8533
rect 11053 8530 11119 8533
rect 19425 8530 19491 8533
rect 19609 8530 19675 8533
rect 3233 8528 6194 8530
rect 3233 8472 3238 8528
rect 3294 8472 6194 8528
rect 3233 8470 6194 8472
rect 3233 8467 3299 8470
rect 0 8394 800 8424
rect 6134 8397 6194 8470
rect 11053 8528 19675 8530
rect 11053 8472 11058 8528
rect 11114 8472 19430 8528
rect 19486 8472 19614 8528
rect 19670 8472 19675 8528
rect 11053 8470 19675 8472
rect 11053 8467 11119 8470
rect 19425 8467 19491 8470
rect 19609 8467 19675 8470
rect 1393 8394 1459 8397
rect 0 8392 1459 8394
rect 0 8336 1398 8392
rect 1454 8336 1459 8392
rect 0 8334 1459 8336
rect 0 8304 800 8334
rect 1393 8331 1459 8334
rect 2865 8394 2931 8397
rect 5165 8394 5231 8397
rect 2865 8392 5231 8394
rect 2865 8336 2870 8392
rect 2926 8336 5170 8392
rect 5226 8336 5231 8392
rect 2865 8334 5231 8336
rect 2865 8331 2931 8334
rect 5165 8331 5231 8334
rect 6085 8392 6194 8397
rect 6085 8336 6090 8392
rect 6146 8336 6194 8392
rect 6085 8334 6194 8336
rect 6085 8331 6151 8334
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 0 7986 800 8016
rect 1393 7986 1459 7989
rect 0 7984 1459 7986
rect 0 7928 1398 7984
rect 1454 7928 1459 7984
rect 0 7926 1459 7928
rect 0 7896 800 7926
rect 1393 7923 1459 7926
rect 5717 7986 5783 7989
rect 6361 7986 6427 7989
rect 5717 7984 6427 7986
rect 5717 7928 5722 7984
rect 5778 7928 6366 7984
rect 6422 7928 6427 7984
rect 5717 7926 6427 7928
rect 5717 7923 5783 7926
rect 6361 7923 6427 7926
rect 6545 7986 6611 7989
rect 13445 7986 13511 7989
rect 6545 7984 13511 7986
rect 6545 7928 6550 7984
rect 6606 7928 13450 7984
rect 13506 7928 13511 7984
rect 6545 7926 13511 7928
rect 6545 7923 6611 7926
rect 13445 7923 13511 7926
rect 4061 7850 4127 7853
rect 9765 7850 9831 7853
rect 11329 7850 11395 7853
rect 4061 7848 9831 7850
rect 4061 7792 4066 7848
rect 4122 7792 9770 7848
rect 9826 7792 9831 7848
rect 4061 7790 9831 7792
rect 4061 7787 4127 7790
rect 9765 7787 9831 7790
rect 9998 7848 11395 7850
rect 9998 7792 11334 7848
rect 11390 7792 11395 7848
rect 9998 7790 11395 7792
rect 7097 7714 7163 7717
rect 9998 7714 10058 7790
rect 11329 7787 11395 7790
rect 12341 7850 12407 7853
rect 15009 7850 15075 7853
rect 12341 7848 15075 7850
rect 12341 7792 12346 7848
rect 12402 7792 15014 7848
rect 15070 7792 15075 7848
rect 12341 7790 15075 7792
rect 12341 7787 12407 7790
rect 15009 7787 15075 7790
rect 7097 7712 10058 7714
rect 7097 7656 7102 7712
rect 7158 7656 10058 7712
rect 7097 7654 10058 7656
rect 7097 7651 7163 7654
rect 6144 7648 6460 7649
rect 0 7578 800 7608
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 1393 7578 1459 7581
rect 0 7576 1459 7578
rect 0 7520 1398 7576
rect 1454 7520 1459 7576
rect 0 7518 1459 7520
rect 0 7488 800 7518
rect 1393 7515 1459 7518
rect 2405 7442 2471 7445
rect 5901 7442 5967 7445
rect 2405 7440 5967 7442
rect 2405 7384 2410 7440
rect 2466 7384 5906 7440
rect 5962 7384 5967 7440
rect 2405 7382 5967 7384
rect 2405 7379 2471 7382
rect 5901 7379 5967 7382
rect 1577 7306 1643 7309
rect 7097 7306 7163 7309
rect 1577 7304 7163 7306
rect 1577 7248 1582 7304
rect 1638 7248 7102 7304
rect 7158 7248 7163 7304
rect 1577 7246 7163 7248
rect 1577 7243 1643 7246
rect 7097 7243 7163 7246
rect 10409 7306 10475 7309
rect 13537 7306 13603 7309
rect 10409 7304 13603 7306
rect 10409 7248 10414 7304
rect 10470 7248 13542 7304
rect 13598 7248 13603 7304
rect 10409 7246 13603 7248
rect 10409 7243 10475 7246
rect 13537 7243 13603 7246
rect 0 7170 800 7200
rect 1669 7170 1735 7173
rect 0 7168 1735 7170
rect 0 7112 1674 7168
rect 1730 7112 1735 7168
rect 0 7110 1735 7112
rect 0 7080 800 7110
rect 1669 7107 1735 7110
rect 9949 7170 10015 7173
rect 12985 7170 13051 7173
rect 9949 7168 13051 7170
rect 9949 7112 9954 7168
rect 10010 7112 12990 7168
rect 13046 7112 13051 7168
rect 9949 7110 13051 7112
rect 9949 7107 10015 7110
rect 12985 7107 13051 7110
rect 3545 7104 3861 7105
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 19139 7039 19455 7040
rect 11697 7034 11763 7037
rect 11654 7032 11763 7034
rect 11654 6976 11702 7032
rect 11758 6976 11763 7032
rect 11654 6971 11763 6976
rect 6545 6898 6611 6901
rect 6821 6898 6887 6901
rect 6545 6896 6887 6898
rect 6545 6840 6550 6896
rect 6606 6840 6826 6896
rect 6882 6840 6887 6896
rect 6545 6838 6887 6840
rect 6545 6835 6611 6838
rect 6821 6835 6887 6838
rect 8518 6836 8524 6900
rect 8588 6898 8594 6900
rect 9121 6898 9187 6901
rect 8588 6896 9187 6898
rect 8588 6840 9126 6896
rect 9182 6840 9187 6896
rect 8588 6838 9187 6840
rect 8588 6836 8594 6838
rect 9121 6835 9187 6838
rect 9581 6898 9647 6901
rect 11654 6898 11714 6971
rect 9581 6896 11714 6898
rect 9581 6840 9586 6896
rect 9642 6840 11714 6896
rect 9581 6838 11714 6840
rect 9581 6835 9647 6838
rect 0 6762 800 6792
rect 1393 6762 1459 6765
rect 0 6760 1459 6762
rect 0 6704 1398 6760
rect 1454 6704 1459 6760
rect 0 6702 1459 6704
rect 0 6672 800 6702
rect 1393 6699 1459 6702
rect 2221 6762 2287 6765
rect 6821 6762 6887 6765
rect 9673 6762 9739 6765
rect 14365 6762 14431 6765
rect 2221 6760 9739 6762
rect 2221 6704 2226 6760
rect 2282 6704 6826 6760
rect 6882 6704 9678 6760
rect 9734 6704 9739 6760
rect 2221 6702 9739 6704
rect 2221 6699 2287 6702
rect 6821 6699 6887 6702
rect 9673 6699 9739 6702
rect 9814 6760 14431 6762
rect 9814 6704 14370 6760
rect 14426 6704 14431 6760
rect 9814 6702 14431 6704
rect 7925 6628 7991 6629
rect 7925 6624 7972 6628
rect 8036 6626 8042 6628
rect 9305 6626 9371 6629
rect 9814 6626 9874 6702
rect 14365 6699 14431 6702
rect 7925 6568 7930 6624
rect 7925 6564 7972 6568
rect 8036 6566 8082 6626
rect 9305 6624 9874 6626
rect 9305 6568 9310 6624
rect 9366 6568 9874 6624
rect 9305 6566 9874 6568
rect 8036 6564 8042 6566
rect 7925 6563 7991 6564
rect 9305 6563 9371 6566
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 21738 6495 22054 6496
rect 0 6354 800 6384
rect 1669 6354 1735 6357
rect 0 6352 1735 6354
rect 0 6296 1674 6352
rect 1730 6296 1735 6352
rect 0 6294 1735 6296
rect 0 6264 800 6294
rect 1669 6291 1735 6294
rect 2773 6354 2839 6357
rect 8293 6354 8359 6357
rect 8569 6354 8635 6357
rect 2773 6352 8635 6354
rect 2773 6296 2778 6352
rect 2834 6296 8298 6352
rect 8354 6296 8574 6352
rect 8630 6296 8635 6352
rect 2773 6294 8635 6296
rect 2773 6291 2839 6294
rect 8293 6291 8359 6294
rect 8569 6291 8635 6294
rect 11789 6354 11855 6357
rect 16481 6354 16547 6357
rect 11789 6352 16547 6354
rect 11789 6296 11794 6352
rect 11850 6296 16486 6352
rect 16542 6296 16547 6352
rect 11789 6294 16547 6296
rect 11789 6291 11855 6294
rect 16481 6291 16547 6294
rect 7557 6218 7623 6221
rect 12065 6218 12131 6221
rect 7557 6216 12131 6218
rect 7557 6160 7562 6216
rect 7618 6160 12070 6216
rect 12126 6160 12131 6216
rect 7557 6158 12131 6160
rect 7557 6155 7623 6158
rect 12065 6155 12131 6158
rect 5942 6020 5948 6084
rect 6012 6082 6018 6084
rect 7005 6082 7071 6085
rect 6012 6080 7071 6082
rect 6012 6024 7010 6080
rect 7066 6024 7071 6080
rect 6012 6022 7071 6024
rect 6012 6020 6018 6022
rect 7005 6019 7071 6022
rect 7741 6082 7807 6085
rect 8385 6082 8451 6085
rect 7741 6080 8451 6082
rect 7741 6024 7746 6080
rect 7802 6024 8390 6080
rect 8446 6024 8451 6080
rect 7741 6022 8451 6024
rect 7741 6019 7807 6022
rect 8385 6019 8451 6022
rect 11329 6082 11395 6085
rect 13445 6082 13511 6085
rect 11329 6080 13511 6082
rect 11329 6024 11334 6080
rect 11390 6024 13450 6080
rect 13506 6024 13511 6080
rect 11329 6022 13511 6024
rect 11329 6019 11395 6022
rect 13445 6019 13511 6022
rect 3545 6016 3861 6017
rect 0 5946 800 5976
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 1393 5946 1459 5949
rect 6545 5946 6611 5949
rect 0 5944 1459 5946
rect 0 5888 1398 5944
rect 1454 5888 1459 5944
rect 0 5886 1459 5888
rect 0 5856 800 5886
rect 1393 5883 1459 5886
rect 5214 5944 6611 5946
rect 5214 5888 6550 5944
rect 6606 5888 6611 5944
rect 5214 5886 6611 5888
rect 1577 5810 1643 5813
rect 5214 5810 5274 5886
rect 6545 5883 6611 5886
rect 10317 5946 10383 5949
rect 12525 5946 12591 5949
rect 10317 5944 12591 5946
rect 10317 5888 10322 5944
rect 10378 5888 12530 5944
rect 12586 5888 12591 5944
rect 10317 5886 12591 5888
rect 10317 5883 10383 5886
rect 12525 5883 12591 5886
rect 1577 5808 5274 5810
rect 1577 5752 1582 5808
rect 1638 5752 5274 5808
rect 1577 5750 5274 5752
rect 5441 5810 5507 5813
rect 10869 5810 10935 5813
rect 5441 5808 10935 5810
rect 5441 5752 5446 5808
rect 5502 5752 10874 5808
rect 10930 5752 10935 5808
rect 5441 5750 10935 5752
rect 1577 5747 1643 5750
rect 5441 5747 5507 5750
rect 10869 5747 10935 5750
rect 12065 5810 12131 5813
rect 12617 5810 12683 5813
rect 12065 5808 12683 5810
rect 12065 5752 12070 5808
rect 12126 5752 12622 5808
rect 12678 5752 12683 5808
rect 12065 5750 12683 5752
rect 12065 5747 12131 5750
rect 12617 5747 12683 5750
rect 21541 5810 21607 5813
rect 22200 5810 23000 5840
rect 21541 5808 23000 5810
rect 21541 5752 21546 5808
rect 21602 5752 23000 5808
rect 21541 5750 23000 5752
rect 21541 5747 21607 5750
rect 22200 5720 23000 5750
rect 5809 5674 5875 5677
rect 8293 5674 8359 5677
rect 5809 5672 8359 5674
rect 5809 5616 5814 5672
rect 5870 5616 8298 5672
rect 8354 5616 8359 5672
rect 5809 5614 8359 5616
rect 5809 5611 5875 5614
rect 8293 5611 8359 5614
rect 9806 5612 9812 5676
rect 9876 5674 9882 5676
rect 10409 5674 10475 5677
rect 9876 5672 10475 5674
rect 9876 5616 10414 5672
rect 10470 5616 10475 5672
rect 9876 5614 10475 5616
rect 9876 5612 9882 5614
rect 10409 5611 10475 5614
rect 11053 5674 11119 5677
rect 15561 5674 15627 5677
rect 16941 5674 17007 5677
rect 11053 5672 17007 5674
rect 11053 5616 11058 5672
rect 11114 5616 15566 5672
rect 15622 5616 16946 5672
rect 17002 5616 17007 5672
rect 11053 5614 17007 5616
rect 11053 5611 11119 5614
rect 15561 5611 15627 5614
rect 16941 5611 17007 5614
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 12433 5538 12499 5541
rect 14733 5538 14799 5541
rect 12433 5536 14799 5538
rect 12433 5480 12438 5536
rect 12494 5480 14738 5536
rect 14794 5480 14799 5536
rect 12433 5478 14799 5480
rect 12433 5475 12499 5478
rect 14733 5475 14799 5478
rect 6144 5472 6460 5473
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 21738 5407 22054 5408
rect 7005 5402 7071 5405
rect 8845 5402 8911 5405
rect 9305 5404 9371 5405
rect 7005 5400 8911 5402
rect 7005 5344 7010 5400
rect 7066 5344 8850 5400
rect 8906 5344 8911 5400
rect 7005 5342 8911 5344
rect 7005 5339 7071 5342
rect 8845 5339 8911 5342
rect 9254 5340 9260 5404
rect 9324 5402 9371 5404
rect 11881 5402 11947 5405
rect 16021 5402 16087 5405
rect 9324 5400 9416 5402
rect 9366 5344 9416 5400
rect 9324 5342 9416 5344
rect 11881 5400 16087 5402
rect 11881 5344 11886 5400
rect 11942 5344 16026 5400
rect 16082 5344 16087 5400
rect 11881 5342 16087 5344
rect 9324 5340 9371 5342
rect 9305 5339 9371 5340
rect 11881 5339 11947 5342
rect 16021 5339 16087 5342
rect 4705 5266 4771 5269
rect 7925 5266 7991 5269
rect 4705 5264 7991 5266
rect 4705 5208 4710 5264
rect 4766 5208 7930 5264
rect 7986 5208 7991 5264
rect 4705 5206 7991 5208
rect 4705 5203 4771 5206
rect 7925 5203 7991 5206
rect 9489 5266 9555 5269
rect 9489 5264 10610 5266
rect 9489 5208 9494 5264
rect 9550 5208 10610 5264
rect 9489 5206 10610 5208
rect 9489 5203 9555 5206
rect 0 5130 800 5160
rect 10550 5133 10610 5206
rect 11094 5204 11100 5268
rect 11164 5266 11170 5268
rect 11421 5266 11487 5269
rect 17401 5266 17467 5269
rect 19517 5266 19583 5269
rect 11164 5264 19583 5266
rect 11164 5208 11426 5264
rect 11482 5208 17406 5264
rect 17462 5208 19522 5264
rect 19578 5208 19583 5264
rect 11164 5206 19583 5208
rect 11164 5204 11170 5206
rect 11421 5203 11487 5206
rect 17401 5203 17467 5206
rect 19517 5203 19583 5206
rect 1669 5130 1735 5133
rect 0 5128 1735 5130
rect 0 5072 1674 5128
rect 1730 5072 1735 5128
rect 0 5070 1735 5072
rect 0 5040 800 5070
rect 1669 5067 1735 5070
rect 6545 5130 6611 5133
rect 10317 5130 10383 5133
rect 6545 5128 10383 5130
rect 6545 5072 6550 5128
rect 6606 5072 10322 5128
rect 10378 5072 10383 5128
rect 6545 5070 10383 5072
rect 10550 5130 10659 5133
rect 15745 5130 15811 5133
rect 10550 5128 15811 5130
rect 10550 5072 10598 5128
rect 10654 5072 15750 5128
rect 15806 5072 15811 5128
rect 10550 5070 15811 5072
rect 6545 5067 6611 5070
rect 10317 5067 10383 5070
rect 10593 5067 10659 5070
rect 15745 5067 15811 5070
rect 9305 4994 9371 4997
rect 11881 4994 11947 4997
rect 9305 4992 11947 4994
rect 9305 4936 9310 4992
rect 9366 4936 11886 4992
rect 11942 4936 11947 4992
rect 9305 4934 11947 4936
rect 9305 4931 9371 4934
rect 11881 4931 11947 4934
rect 12525 4994 12591 4997
rect 13353 4994 13419 4997
rect 12525 4992 13419 4994
rect 12525 4936 12530 4992
rect 12586 4936 13358 4992
rect 13414 4936 13419 4992
rect 12525 4934 13419 4936
rect 12525 4931 12591 4934
rect 13353 4931 13419 4934
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 19139 4863 19455 4864
rect 10910 4796 10916 4860
rect 10980 4858 10986 4860
rect 11329 4858 11395 4861
rect 10980 4856 11395 4858
rect 10980 4800 11334 4856
rect 11390 4800 11395 4856
rect 10980 4798 11395 4800
rect 10980 4796 10986 4798
rect 11329 4795 11395 4798
rect 12198 4796 12204 4860
rect 12268 4858 12274 4860
rect 12617 4858 12683 4861
rect 12268 4856 12683 4858
rect 12268 4800 12622 4856
rect 12678 4800 12683 4856
rect 12268 4798 12683 4800
rect 12268 4796 12274 4798
rect 12617 4795 12683 4798
rect 0 4722 800 4752
rect 1485 4722 1551 4725
rect 0 4720 1551 4722
rect 0 4664 1490 4720
rect 1546 4664 1551 4720
rect 0 4662 1551 4664
rect 0 4632 800 4662
rect 1485 4659 1551 4662
rect 9673 4722 9739 4725
rect 17401 4722 17467 4725
rect 9673 4720 17467 4722
rect 9673 4664 9678 4720
rect 9734 4664 17406 4720
rect 17462 4664 17467 4720
rect 9673 4662 17467 4664
rect 9673 4659 9739 4662
rect 17401 4659 17467 4662
rect 8017 4586 8083 4589
rect 13721 4586 13787 4589
rect 17125 4586 17191 4589
rect 8017 4584 12450 4586
rect 8017 4528 8022 4584
rect 8078 4528 12450 4584
rect 8017 4526 12450 4528
rect 8017 4523 8083 4526
rect 6144 4384 6460 4385
rect 0 4314 800 4344
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 2221 4314 2287 4317
rect 0 4312 2287 4314
rect 0 4256 2226 4312
rect 2282 4256 2287 4312
rect 0 4254 2287 4256
rect 0 4224 800 4254
rect 2221 4251 2287 4254
rect 8293 4314 8359 4317
rect 9029 4314 9095 4317
rect 11053 4314 11119 4317
rect 8293 4312 11119 4314
rect 8293 4256 8298 4312
rect 8354 4256 9034 4312
rect 9090 4256 11058 4312
rect 11114 4256 11119 4312
rect 8293 4254 11119 4256
rect 12390 4314 12450 4526
rect 13721 4584 17191 4586
rect 13721 4528 13726 4584
rect 13782 4528 17130 4584
rect 17186 4528 17191 4584
rect 13721 4526 17191 4528
rect 13721 4523 13787 4526
rect 17125 4523 17191 4526
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 16297 4314 16363 4317
rect 12390 4312 16363 4314
rect 12390 4256 16302 4312
rect 16358 4256 16363 4312
rect 12390 4254 16363 4256
rect 8293 4251 8359 4254
rect 9029 4251 9095 4254
rect 11053 4251 11119 4254
rect 16297 4251 16363 4254
rect 6545 4178 6611 4181
rect 10685 4178 10751 4181
rect 14457 4178 14523 4181
rect 6545 4176 14523 4178
rect 6545 4120 6550 4176
rect 6606 4120 10690 4176
rect 10746 4120 14462 4176
rect 14518 4120 14523 4176
rect 6545 4118 14523 4120
rect 6545 4115 6611 4118
rect 10685 4115 10751 4118
rect 14457 4115 14523 4118
rect 15837 4178 15903 4181
rect 21357 4178 21423 4181
rect 15837 4176 21423 4178
rect 15837 4120 15842 4176
rect 15898 4120 21362 4176
rect 21418 4120 21423 4176
rect 15837 4118 21423 4120
rect 15837 4115 15903 4118
rect 21357 4115 21423 4118
rect 5257 4042 5323 4045
rect 5390 4042 5396 4044
rect 5257 4040 5396 4042
rect 5257 3984 5262 4040
rect 5318 3984 5396 4040
rect 5257 3982 5396 3984
rect 5257 3979 5323 3982
rect 5390 3980 5396 3982
rect 5460 3980 5466 4044
rect 8109 4042 8175 4045
rect 12065 4042 12131 4045
rect 8109 4040 12131 4042
rect 8109 3984 8114 4040
rect 8170 3984 12070 4040
rect 12126 3984 12131 4040
rect 8109 3982 12131 3984
rect 8109 3979 8175 3982
rect 12065 3979 12131 3982
rect 0 3906 800 3936
rect 2221 3906 2287 3909
rect 0 3904 2287 3906
rect 0 3848 2226 3904
rect 2282 3848 2287 3904
rect 0 3846 2287 3848
rect 0 3816 800 3846
rect 2221 3843 2287 3846
rect 10501 3906 10567 3909
rect 11329 3906 11395 3909
rect 10501 3904 11395 3906
rect 10501 3848 10506 3904
rect 10562 3848 11334 3904
rect 11390 3848 11395 3904
rect 10501 3846 11395 3848
rect 10501 3843 10567 3846
rect 11329 3843 11395 3846
rect 3545 3840 3861 3841
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 19139 3775 19455 3776
rect 7741 3770 7807 3773
rect 5950 3768 7807 3770
rect 5950 3712 7746 3768
rect 7802 3712 7807 3768
rect 5950 3710 7807 3712
rect 2497 3634 2563 3637
rect 5950 3634 6010 3710
rect 7741 3707 7807 3710
rect 9121 3770 9187 3773
rect 11513 3770 11579 3773
rect 11973 3770 12039 3773
rect 13813 3770 13879 3773
rect 9121 3768 11898 3770
rect 9121 3712 9126 3768
rect 9182 3712 11518 3768
rect 11574 3712 11898 3768
rect 9121 3710 11898 3712
rect 9121 3707 9187 3710
rect 11513 3707 11579 3710
rect 2497 3632 6010 3634
rect 2497 3576 2502 3632
rect 2558 3576 6010 3632
rect 2497 3574 6010 3576
rect 6177 3634 6243 3637
rect 9305 3634 9371 3637
rect 6177 3632 9371 3634
rect 6177 3576 6182 3632
rect 6238 3576 9310 3632
rect 9366 3576 9371 3632
rect 6177 3574 9371 3576
rect 2497 3571 2563 3574
rect 6177 3571 6243 3574
rect 9305 3571 9371 3574
rect 9489 3634 9555 3637
rect 10593 3634 10659 3637
rect 9489 3632 10659 3634
rect 9489 3576 9494 3632
rect 9550 3576 10598 3632
rect 10654 3576 10659 3632
rect 9489 3574 10659 3576
rect 11838 3634 11898 3710
rect 11973 3768 13879 3770
rect 11973 3712 11978 3768
rect 12034 3712 13818 3768
rect 13874 3712 13879 3768
rect 11973 3710 13879 3712
rect 11973 3707 12039 3710
rect 13813 3707 13879 3710
rect 15285 3634 15351 3637
rect 11838 3632 15351 3634
rect 11838 3576 15290 3632
rect 15346 3576 15351 3632
rect 11838 3574 15351 3576
rect 9489 3571 9555 3574
rect 10593 3571 10659 3574
rect 15285 3571 15351 3574
rect 0 3498 800 3528
rect 1485 3498 1551 3501
rect 0 3496 1551 3498
rect 0 3440 1490 3496
rect 1546 3440 1551 3496
rect 0 3438 1551 3440
rect 0 3408 800 3438
rect 1485 3435 1551 3438
rect 1669 3498 1735 3501
rect 12617 3498 12683 3501
rect 1669 3496 7298 3498
rect 1669 3440 1674 3496
rect 1730 3440 7298 3496
rect 1669 3438 7298 3440
rect 1669 3435 1735 3438
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 7238 3226 7298 3438
rect 8526 3496 12683 3498
rect 8526 3440 12622 3496
rect 12678 3440 12683 3496
rect 8526 3438 12683 3440
rect 7373 3362 7439 3365
rect 8526 3362 8586 3438
rect 12617 3435 12683 3438
rect 7373 3360 8586 3362
rect 7373 3304 7378 3360
rect 7434 3304 8586 3360
rect 7373 3302 8586 3304
rect 7373 3299 7439 3302
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 21738 3231 22054 3232
rect 8569 3226 8635 3229
rect 7238 3224 8635 3226
rect 7238 3168 8574 3224
rect 8630 3168 8635 3224
rect 7238 3166 8635 3168
rect 8569 3163 8635 3166
rect 13077 3226 13143 3229
rect 15929 3226 15995 3229
rect 13077 3224 15995 3226
rect 13077 3168 13082 3224
rect 13138 3168 15934 3224
rect 15990 3168 15995 3224
rect 13077 3166 15995 3168
rect 13077 3163 13143 3166
rect 15929 3163 15995 3166
rect 0 3090 800 3120
rect 1853 3090 1919 3093
rect 0 3088 1919 3090
rect 0 3032 1858 3088
rect 1914 3032 1919 3088
rect 0 3030 1919 3032
rect 0 3000 800 3030
rect 1853 3027 1919 3030
rect 2313 3090 2379 3093
rect 7649 3090 7715 3093
rect 2313 3088 7715 3090
rect 2313 3032 2318 3088
rect 2374 3032 7654 3088
rect 7710 3032 7715 3088
rect 2313 3030 7715 3032
rect 2313 3027 2379 3030
rect 7649 3027 7715 3030
rect 10317 3090 10383 3093
rect 15101 3090 15167 3093
rect 10317 3088 15167 3090
rect 10317 3032 10322 3088
rect 10378 3032 15106 3088
rect 15162 3032 15167 3088
rect 10317 3030 15167 3032
rect 10317 3027 10383 3030
rect 15101 3027 15167 3030
rect 17401 3090 17467 3093
rect 19333 3090 19399 3093
rect 17401 3088 19399 3090
rect 17401 3032 17406 3088
rect 17462 3032 19338 3088
rect 19394 3032 19399 3088
rect 17401 3030 19399 3032
rect 17401 3027 17467 3030
rect 19333 3027 19399 3030
rect 3545 2752 3861 2753
rect 0 2682 800 2712
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 2773 2682 2839 2685
rect 0 2680 2839 2682
rect 0 2624 2778 2680
rect 2834 2624 2839 2680
rect 0 2622 2839 2624
rect 0 2592 800 2622
rect 2773 2619 2839 2622
rect 9213 2410 9279 2413
rect 9438 2410 9444 2412
rect 9213 2408 9444 2410
rect 9213 2352 9218 2408
rect 9274 2352 9444 2408
rect 9213 2350 9444 2352
rect 9213 2347 9279 2350
rect 9438 2348 9444 2350
rect 9508 2348 9514 2412
rect 0 2274 800 2304
rect 2221 2274 2287 2277
rect 0 2272 2287 2274
rect 0 2216 2226 2272
rect 2282 2216 2287 2272
rect 0 2214 2287 2216
rect 0 2184 800 2214
rect 2221 2211 2287 2214
rect 6144 2208 6460 2209
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 21738 2143 22054 2144
rect 0 1866 800 1896
rect 2129 1866 2195 1869
rect 0 1864 2195 1866
rect 0 1808 2134 1864
rect 2190 1808 2195 1864
rect 0 1806 2195 1808
rect 0 1776 800 1806
rect 2129 1803 2195 1806
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 5396 19348 5460 19412
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 9996 19484 10060 19548
rect 5948 19348 6012 19412
rect 7972 19348 8036 19412
rect 9260 19408 9324 19412
rect 9260 19352 9274 19408
rect 9274 19352 9324 19408
rect 9260 19348 9324 19352
rect 10364 19348 10428 19412
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 11100 19212 11164 19276
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 8156 18804 8220 18868
rect 9444 18592 9508 18596
rect 9444 18536 9458 18592
rect 9458 18536 9508 18592
rect 9444 18532 9508 18536
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 7604 18396 7668 18460
rect 6868 18260 6932 18324
rect 8340 18124 8404 18188
rect 2452 17988 2516 18052
rect 9444 18048 9508 18052
rect 9444 17992 9458 18048
rect 9458 17992 9508 18048
rect 9444 17988 9508 17992
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 9812 16900 9876 16964
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 6868 16220 6932 16284
rect 7788 16220 7852 16284
rect 5764 15812 5828 15876
rect 9444 16008 9508 16012
rect 9444 15952 9458 16008
rect 9458 15952 9508 16008
rect 9444 15948 9508 15952
rect 11836 15948 11900 16012
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 8524 15540 8588 15604
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 8156 15056 8220 15060
rect 8156 15000 8170 15056
rect 8170 15000 8220 15056
rect 8156 14996 8220 15000
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 8156 14452 8220 14516
rect 5212 14316 5276 14380
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 6868 13636 6932 13700
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 5396 13500 5460 13564
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 6868 12608 6932 12612
rect 6868 12552 6882 12608
rect 6882 12552 6932 12608
rect 6868 12548 6932 12552
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 6684 12412 6748 12476
rect 6684 12064 6748 12068
rect 6684 12008 6734 12064
rect 6734 12008 6748 12064
rect 6684 12004 6748 12008
rect 10916 12004 10980 12068
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 8156 11868 8220 11932
rect 11836 11732 11900 11796
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 9996 11384 10060 11388
rect 9996 11328 10010 11384
rect 10010 11328 10060 11384
rect 9996 11324 10060 11328
rect 12204 11324 12268 11388
rect 5764 11248 5828 11252
rect 5764 11192 5778 11248
rect 5778 11192 5828 11248
rect 5764 11188 5828 11192
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 7604 10780 7668 10844
rect 10364 10840 10428 10844
rect 10364 10784 10414 10840
rect 10414 10784 10428 10840
rect 10364 10780 10428 10784
rect 7604 10508 7668 10572
rect 8524 10508 8588 10572
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 5212 10236 5276 10300
rect 7788 10100 7852 10164
rect 5396 9828 5460 9892
rect 8340 9828 8404 9892
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 2452 9480 2516 9484
rect 2452 9424 2466 9480
rect 2466 9424 2516 9480
rect 2452 9420 2516 9424
rect 9812 9480 9876 9484
rect 9812 9424 9826 9480
rect 9826 9424 9876 9480
rect 9812 9420 9876 9424
rect 8524 9344 8588 9348
rect 8524 9288 8538 9344
rect 8538 9288 8588 9344
rect 8524 9284 8588 9288
rect 9812 9344 9876 9348
rect 9812 9288 9826 9344
rect 9826 9288 9876 9344
rect 9812 9284 9876 9288
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 8524 6836 8588 6900
rect 7972 6624 8036 6628
rect 7972 6568 7986 6624
rect 7986 6568 8036 6624
rect 7972 6564 8036 6568
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 5948 6020 6012 6084
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 9812 5612 9876 5676
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 9260 5400 9324 5404
rect 9260 5344 9310 5400
rect 9310 5344 9324 5400
rect 9260 5340 9324 5344
rect 11100 5204 11164 5268
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 10916 4796 10980 4860
rect 12204 4796 12268 4860
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 5396 3980 5460 4044
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 9444 2348 9508 2412
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 5395 19412 5461 19413
rect 5395 19348 5396 19412
rect 5460 19348 5461 19412
rect 5395 19347 5461 19348
rect 5947 19412 6013 19413
rect 5947 19348 5948 19412
rect 6012 19348 6013 19412
rect 5947 19347 6013 19348
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 2451 18052 2517 18053
rect 2451 17988 2452 18052
rect 2516 17988 2517 18052
rect 2451 17987 2517 17988
rect 2454 9485 2514 17987
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 5211 14380 5277 14381
rect 5211 14316 5212 14380
rect 5276 14316 5277 14380
rect 5211 14315 5277 14316
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 2451 9484 2517 9485
rect 2451 9420 2452 9484
rect 2516 9420 2517 9484
rect 2451 9419 2517 9420
rect 3543 9280 3863 10304
rect 5214 10301 5274 14315
rect 5398 13565 5458 19347
rect 5763 15876 5829 15877
rect 5763 15812 5764 15876
rect 5828 15812 5829 15876
rect 5763 15811 5829 15812
rect 5395 13564 5461 13565
rect 5395 13500 5396 13564
rect 5460 13500 5461 13564
rect 5395 13499 5461 13500
rect 5766 11253 5826 15811
rect 5763 11252 5829 11253
rect 5763 11188 5764 11252
rect 5828 11188 5829 11252
rect 5763 11187 5829 11188
rect 5211 10300 5277 10301
rect 5211 10236 5212 10300
rect 5276 10236 5277 10300
rect 5211 10235 5277 10236
rect 5395 9892 5461 9893
rect 5395 9828 5396 9892
rect 5460 9828 5461 9892
rect 5395 9827 5461 9828
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 5398 4045 5458 9827
rect 5950 6085 6010 19347
rect 6142 18528 6462 19552
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 7971 19412 8037 19413
rect 7971 19348 7972 19412
rect 8036 19348 8037 19412
rect 7971 19347 8037 19348
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 7603 18460 7669 18461
rect 7603 18396 7604 18460
rect 7668 18396 7669 18460
rect 7603 18395 7669 18396
rect 6867 18324 6933 18325
rect 6867 18260 6868 18324
rect 6932 18260 6933 18324
rect 6867 18259 6933 18260
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6870 16285 6930 18259
rect 6867 16284 6933 16285
rect 6867 16220 6868 16284
rect 6932 16220 6933 16284
rect 6867 16219 6933 16220
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6867 13700 6933 13701
rect 6867 13636 6868 13700
rect 6932 13636 6933 13700
rect 6867 13635 6933 13636
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6870 12613 6930 13635
rect 6867 12612 6933 12613
rect 6867 12548 6868 12612
rect 6932 12548 6933 12612
rect 6867 12547 6933 12548
rect 6683 12476 6749 12477
rect 6683 12412 6684 12476
rect 6748 12412 6749 12476
rect 6683 12411 6749 12412
rect 6686 12069 6746 12411
rect 6683 12068 6749 12069
rect 6683 12004 6684 12068
rect 6748 12004 6749 12068
rect 6683 12003 6749 12004
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 7606 10845 7666 18395
rect 7787 16284 7853 16285
rect 7787 16220 7788 16284
rect 7852 16220 7853 16284
rect 7787 16219 7853 16220
rect 7603 10844 7669 10845
rect 7603 10780 7604 10844
rect 7668 10780 7669 10844
rect 7603 10779 7669 10780
rect 7606 10573 7666 10779
rect 7603 10572 7669 10573
rect 7603 10508 7604 10572
rect 7668 10508 7669 10572
rect 7603 10507 7669 10508
rect 7790 10165 7850 16219
rect 7787 10164 7853 10165
rect 7787 10100 7788 10164
rect 7852 10100 7853 10164
rect 7787 10099 7853 10100
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 7974 6629 8034 19347
rect 8741 19072 9061 20096
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 9995 19548 10061 19549
rect 9995 19484 9996 19548
rect 10060 19484 10061 19548
rect 9995 19483 10061 19484
rect 9259 19412 9325 19413
rect 9259 19348 9260 19412
rect 9324 19348 9325 19412
rect 9259 19347 9325 19348
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8155 18868 8221 18869
rect 8155 18804 8156 18868
rect 8220 18804 8221 18868
rect 8155 18803 8221 18804
rect 8158 15061 8218 18803
rect 8339 18188 8405 18189
rect 8339 18124 8340 18188
rect 8404 18124 8405 18188
rect 8339 18123 8405 18124
rect 8155 15060 8221 15061
rect 8155 14996 8156 15060
rect 8220 14996 8221 15060
rect 8155 14995 8221 14996
rect 8155 14516 8221 14517
rect 8155 14452 8156 14516
rect 8220 14452 8221 14516
rect 8155 14451 8221 14452
rect 8158 11933 8218 14451
rect 8155 11932 8221 11933
rect 8155 11868 8156 11932
rect 8220 11868 8221 11932
rect 8155 11867 8221 11868
rect 8342 9893 8402 18123
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8523 15604 8589 15605
rect 8523 15540 8524 15604
rect 8588 15540 8589 15604
rect 8523 15539 8589 15540
rect 8526 10573 8586 15539
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8523 10572 8589 10573
rect 8523 10508 8524 10572
rect 8588 10508 8589 10572
rect 8523 10507 8589 10508
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8339 9892 8405 9893
rect 8339 9828 8340 9892
rect 8404 9828 8405 9892
rect 8339 9827 8405 9828
rect 8523 9348 8589 9349
rect 8523 9284 8524 9348
rect 8588 9284 8589 9348
rect 8523 9283 8589 9284
rect 8526 6901 8586 9283
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8523 6900 8589 6901
rect 8523 6836 8524 6900
rect 8588 6836 8589 6900
rect 8523 6835 8589 6836
rect 7971 6628 8037 6629
rect 7971 6564 7972 6628
rect 8036 6564 8037 6628
rect 7971 6563 8037 6564
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 5947 6084 6013 6085
rect 5947 6020 5948 6084
rect 6012 6020 6013 6084
rect 5947 6019 6013 6020
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 5395 4044 5461 4045
rect 5395 3980 5396 4044
rect 5460 3980 5461 4044
rect 5395 3979 5461 3980
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 9262 5405 9322 19347
rect 9443 18596 9509 18597
rect 9443 18532 9444 18596
rect 9508 18532 9509 18596
rect 9443 18531 9509 18532
rect 9446 18053 9506 18531
rect 9443 18052 9509 18053
rect 9443 17988 9444 18052
rect 9508 17988 9509 18052
rect 9443 17987 9509 17988
rect 9811 16964 9877 16965
rect 9811 16900 9812 16964
rect 9876 16900 9877 16964
rect 9811 16899 9877 16900
rect 9443 16012 9509 16013
rect 9443 15948 9444 16012
rect 9508 15948 9509 16012
rect 9443 15947 9509 15948
rect 9259 5404 9325 5405
rect 9259 5340 9260 5404
rect 9324 5340 9325 5404
rect 9259 5339 9325 5340
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 9446 2413 9506 15947
rect 9814 9485 9874 16899
rect 9998 11389 10058 19483
rect 10363 19412 10429 19413
rect 10363 19348 10364 19412
rect 10428 19348 10429 19412
rect 10363 19347 10429 19348
rect 9995 11388 10061 11389
rect 9995 11324 9996 11388
rect 10060 11324 10061 11388
rect 9995 11323 10061 11324
rect 10366 10845 10426 19347
rect 11099 19276 11165 19277
rect 11099 19212 11100 19276
rect 11164 19212 11165 19276
rect 11099 19211 11165 19212
rect 10915 12068 10981 12069
rect 10915 12004 10916 12068
rect 10980 12004 10981 12068
rect 10915 12003 10981 12004
rect 10363 10844 10429 10845
rect 10363 10780 10364 10844
rect 10428 10780 10429 10844
rect 10363 10779 10429 10780
rect 9811 9484 9877 9485
rect 9811 9420 9812 9484
rect 9876 9420 9877 9484
rect 9811 9419 9877 9420
rect 9811 9348 9877 9349
rect 9811 9284 9812 9348
rect 9876 9284 9877 9348
rect 9811 9283 9877 9284
rect 9814 5677 9874 9283
rect 9811 5676 9877 5677
rect 9811 5612 9812 5676
rect 9876 5612 9877 5676
rect 9811 5611 9877 5612
rect 10918 4861 10978 12003
rect 11102 5269 11162 19211
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 11835 16012 11901 16013
rect 11835 15948 11836 16012
rect 11900 15948 11901 16012
rect 11835 15947 11901 15948
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11838 11797 11898 15947
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 11835 11796 11901 11797
rect 11835 11732 11836 11796
rect 11900 11732 11901 11796
rect 11835 11731 11901 11732
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 12203 11388 12269 11389
rect 12203 11324 12204 11388
rect 12268 11324 12269 11388
rect 12203 11323 12269 11324
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11099 5268 11165 5269
rect 11099 5204 11100 5268
rect 11164 5204 11165 5268
rect 11099 5203 11165 5204
rect 10915 4860 10981 4861
rect 10915 4796 10916 4860
rect 10980 4796 10981 4860
rect 10915 4795 10981 4796
rect 11340 4384 11660 5408
rect 12206 4861 12266 11323
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 12203 4860 12269 4861
rect 12203 4796 12204 4860
rect 12268 4796 12269 4860
rect 12203 4795 12269 4796
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 9443 2412 9509 2413
rect 9443 2348 9444 2412
rect 9508 2348 9509 2412
rect 9443 2347 9509 2348
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1649977179
transform -1 0 12696 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1649977179
transform -1 0 15364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1649977179
transform 1 0 16836 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1649977179
transform -1 0 17388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1649977179
transform -1 0 17848 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1649977179
transform -1 0 19780 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1649977179
transform 1 0 19964 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1649977179
transform -1 0 15640 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1649977179
transform -1 0 16100 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1649977179
transform 1 0 18400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1649977179
transform -1 0 18032 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1649977179
transform -1 0 19596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1649977179
transform 1 0 7360 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1649977179
transform 1 0 6808 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1649977179
transform -1 0 6808 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1649977179
transform 1 0 7912 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1649977179
transform -1 0 9476 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1649977179
transform 1 0 8832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1649977179
transform 1 0 10028 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1649977179
transform -1 0 14996 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1649977179
transform -1 0 8740 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1649977179
transform -1 0 7912 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1649977179
transform -1 0 8832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1649977179
transform -1 0 14812 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1649977179
transform -1 0 16284 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 2852 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 3404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 2484 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 3036 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 3956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 3404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 2760 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 3772 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 21344 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 21344 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 2668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 2852 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 2116 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 1564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 1840 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 1840 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 2116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 2300 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 1840 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 2116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 2300 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 2116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 2300 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 2484 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 2484 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 2116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 2300 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 1840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 3220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 8464 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 8096 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 8280 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 9292 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 12052 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 11132 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 11868 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 12880 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 13064 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 14444 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 3680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 4232 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 5888 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 4600 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 6256 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 7360 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 7820 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 4324 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 8280 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 7728 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 8096 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 10672 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 10856 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 11408 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 8832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 13984 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 13708 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 4600 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 5152 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 5336 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 6532 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 6072 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 5888 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 6256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 7728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1649977179
transform -1 0 7176 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1649977179
transform -1 0 3036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1649977179
transform -1 0 3588 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1649977179
transform -1 0 3588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1649977179
transform -1 0 3220 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1649977179
transform -1 0 2852 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1649977179
transform -1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1649977179
transform -1 0 2484 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1649977179
transform -1 0 2852 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1649977179
transform -1 0 2484 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1649977179
transform -1 0 2208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1649977179
transform -1 0 2668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1649977179
transform -1 0 3128 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1649977179
transform -1 0 3312 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1649977179
transform -1 0 2852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1649977179
transform -1 0 3036 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1649977179
transform -1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1649977179
transform -1 0 19504 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 13524 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16008 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13892 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 11592 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13156 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20792 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21344 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18124 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform -1 0 18492 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 17756 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13340 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 13524 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20792 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20884 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 21252 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 21344 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20792 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18584 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 21160 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21344 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15916 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 16100 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18124 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18400 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 13708 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13524 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14168 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14352 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15640 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13984 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12512 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17112 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20608 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 20792 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18124 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21068 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16928 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19964 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 20976 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16744 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18124 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21160 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19780 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19596 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17664 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 20424 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 21344 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21252 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18124 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18124 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14536 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12972 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16192 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 19964 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17756 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15824 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform -1 0 16192 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13248 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13616 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13524 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13064 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13340 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 17940 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19596 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 18308 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13156 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 20700 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 19412 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15548 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 15732 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15916 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15272 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 15456 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18124 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18216 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11316 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 10764 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 9292 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10580 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12696 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12512 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 13984 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 9292 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_6__S
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16100 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 16468 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 4692 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12052 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 13524 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 8740 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 5520 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 5152 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17204 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 18400 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 9752 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 12696 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9200 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 5152 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 5428 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 5428 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 7360 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5888 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 4416 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 7360 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7268 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 7268 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6072 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5704 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 5888 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 7268 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 6256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 7268 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7268 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6900 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8556 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 7728 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7452 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 9108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 7544 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11684 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 9936 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14904 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14720 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15824 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 11868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17664 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17480 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 14352 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9752 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8740 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 13524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9844 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8096 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11040 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8372 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10948 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 11132 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11776 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11132 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9384 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9936 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7636 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5888 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7728 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 8464 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 9936 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 10120 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1649977179
transform -1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 7176 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8280 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 7360 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 8372 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A1
timestamp 1649977179
transform 1 0 8556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 9752 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 9936 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 9200 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 10396 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 5336 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 5428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 4692 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 11132 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 9108 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 10948 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__S
timestamp 1649977179
transform -1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 3220 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 12328 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 2944 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 4600 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 18768 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater151_A
timestamp 1649977179
transform 1 0 11500 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1649977179
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_157
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_162
timestamp 1649977179
transform 1 0 16008 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1649977179
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_182
timestamp 1649977179
transform 1 0 17848 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_187
timestamp 1649977179
transform 1 0 18308 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_217
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222
timestamp 1649977179
transform 1 0 21528 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_31
timestamp 1649977179
transform 1 0 3956 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_53
timestamp 1649977179
transform 1 0 5980 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_155
timestamp 1649977179
transform 1 0 15364 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_177 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_203
timestamp 1649977179
transform 1 0 19780 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_210
timestamp 1649977179
transform 1 0 20424 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_214
timestamp 1649977179
transform 1 0 20792 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_52
timestamp 1649977179
transform 1 0 5888 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_56
timestamp 1649977179
transform 1 0 6256 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_73
timestamp 1649977179
transform 1 0 7820 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_128
timestamp 1649977179
transform 1 0 12880 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_145 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_157
timestamp 1649977179
transform 1 0 15548 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_169 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16652 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_179 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17572 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_187
timestamp 1649977179
transform 1 0 18308 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_190
timestamp 1649977179
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_207
timestamp 1649977179
transform 1 0 20148 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_215
timestamp 1649977179
transform 1 0 20884 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_21
timestamp 1649977179
transform 1 0 3036 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_33
timestamp 1649977179
transform 1 0 4140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_45
timestamp 1649977179
transform 1 0 5244 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_66
timestamp 1649977179
transform 1 0 7176 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_86
timestamp 1649977179
transform 1 0 9016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_130
timestamp 1649977179
transform 1 0 13064 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_142
timestamp 1649977179
transform 1 0 14168 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_147
timestamp 1649977179
transform 1 0 14628 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_159
timestamp 1649977179
transform 1 0 15732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_178
timestamp 1649977179
transform 1 0 17480 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_190
timestamp 1649977179
transform 1 0 18584 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_202
timestamp 1649977179
transform 1 0 19688 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_214
timestamp 1649977179
transform 1 0 20792 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_222
timestamp 1649977179
transform 1 0 21528 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_55
timestamp 1649977179
transform 1 0 6164 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_69
timestamp 1649977179
transform 1 0 7452 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_87
timestamp 1649977179
transform 1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1649977179
transform 1 0 9476 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_123
timestamp 1649977179
transform 1 0 12420 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 1649977179
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_167
timestamp 1649977179
transform 1 0 16468 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_173
timestamp 1649977179
transform 1 0 17020 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_185
timestamp 1649977179
transform 1 0 18124 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_191
timestamp 1649977179
transform 1 0 18676 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_19
timestamp 1649977179
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_31
timestamp 1649977179
transform 1 0 3956 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_66
timestamp 1649977179
transform 1 0 7176 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_83
timestamp 1649977179
transform 1 0 8740 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_87
timestamp 1649977179
transform 1 0 9108 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_163
timestamp 1649977179
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_176
timestamp 1649977179
transform 1 0 17296 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_188
timestamp 1649977179
transform 1 0 18400 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_200
timestamp 1649977179
transform 1 0 19504 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_215
timestamp 1649977179
transform 1 0 20884 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_11
timestamp 1649977179
transform 1 0 2116 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_19
timestamp 1649977179
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_43
timestamp 1649977179
transform 1 0 5060 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_46
timestamp 1649977179
transform 1 0 5336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_69
timestamp 1649977179
transform 1 0 7452 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_96
timestamp 1649977179
transform 1 0 9936 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_100
timestamp 1649977179
transform 1 0 10304 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_110
timestamp 1649977179
transform 1 0 11224 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1649977179
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_186
timestamp 1649977179
transform 1 0 18216 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_214
timestamp 1649977179
transform 1 0 20792 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_222
timestamp 1649977179
transform 1 0 21528 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_31
timestamp 1649977179
transform 1 0 3956 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1649977179
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_92
timestamp 1649977179
transform 1 0 9568 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_102
timestamp 1649977179
transform 1 0 10488 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_120
timestamp 1649977179
transform 1 0 12144 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_130
timestamp 1649977179
transform 1 0 13064 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_138
timestamp 1649977179
transform 1 0 13800 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_148
timestamp 1649977179
transform 1 0 14720 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_160
timestamp 1649977179
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_49
timestamp 1649977179
transform 1 0 5612 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_80
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_107
timestamp 1649977179
transform 1 0 10948 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_115
timestamp 1649977179
transform 1 0 11684 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_125
timestamp 1649977179
transform 1 0 12604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_137
timestamp 1649977179
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_152
timestamp 1649977179
transform 1 0 15088 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_164
timestamp 1649977179
transform 1 0 16192 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_176
timestamp 1649977179
transform 1 0 17296 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_188
timestamp 1649977179
transform 1 0 18400 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_35
timestamp 1649977179
transform 1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_98
timestamp 1649977179
transform 1 0 10120 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_116
timestamp 1649977179
transform 1 0 11776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_131
timestamp 1649977179
transform 1 0 13156 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_197
timestamp 1649977179
transform 1 0 19228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_216
timestamp 1649977179
transform 1 0 20976 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_222
timestamp 1649977179
transform 1 0 21528 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_6
timestamp 1649977179
transform 1 0 1656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_21
timestamp 1649977179
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_57
timestamp 1649977179
transform 1 0 6348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_72
timestamp 1649977179
transform 1 0 7728 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1649977179
transform 1 0 9660 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_103
timestamp 1649977179
transform 1 0 10580 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_107
timestamp 1649977179
transform 1 0 10948 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_128
timestamp 1649977179
transform 1 0 12880 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_146
timestamp 1649977179
transform 1 0 14536 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_150
timestamp 1649977179
transform 1 0 14904 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_171
timestamp 1649977179
transform 1 0 16836 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_191
timestamp 1649977179
transform 1 0 18676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_219
timestamp 1649977179
transform 1 0 21252 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_22
timestamp 1649977179
transform 1 0 3128 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_30
timestamp 1649977179
transform 1 0 3864 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_46
timestamp 1649977179
transform 1 0 5336 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_59
timestamp 1649977179
transform 1 0 6532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_116
timestamp 1649977179
transform 1 0 11776 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_120
timestamp 1649977179
transform 1 0 12144 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_141
timestamp 1649977179
transform 1 0 14076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_160
timestamp 1649977179
transform 1 0 15824 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_214
timestamp 1649977179
transform 1 0 20792 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_222
timestamp 1649977179
transform 1 0 21528 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1649977179
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_33
timestamp 1649977179
transform 1 0 4140 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_114
timestamp 1649977179
transform 1 0 11592 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_118
timestamp 1649977179
transform 1 0 11960 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_137
timestamp 1649977179
transform 1 0 13708 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_159
timestamp 1649977179
transform 1 0 15732 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_183
timestamp 1649977179
transform 1 0 17940 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_187
timestamp 1649977179
transform 1 0 18308 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_218
timestamp 1649977179
transform 1 0 21160 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_222
timestamp 1649977179
transform 1 0 21528 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_22
timestamp 1649977179
transform 1 0 3128 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_34
timestamp 1649977179
transform 1 0 4232 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 1649977179
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_68
timestamp 1649977179
transform 1 0 7360 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_80
timestamp 1649977179
transform 1 0 8464 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_118
timestamp 1649977179
transform 1 0 11960 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1649977179
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_222
timestamp 1649977179
transform 1 0 21528 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_43
timestamp 1649977179
transform 1 0 5060 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1649977179
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_216
timestamp 1649977179
transform 1 0 20976 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_220
timestamp 1649977179
transform 1 0 21344 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_8
timestamp 1649977179
transform 1 0 1840 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_20
timestamp 1649977179
transform 1 0 2944 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_32
timestamp 1649977179
transform 1 0 4048 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_68
timestamp 1649977179
transform 1 0 7360 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_99
timestamp 1649977179
transform 1 0 10212 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1649977179
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_187
timestamp 1649977179
transform 1 0 18308 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_14
timestamp 1649977179
transform 1 0 2392 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1649977179
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_35
timestamp 1649977179
transform 1 0 4324 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_70
timestamp 1649977179
transform 1 0 7544 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_78
timestamp 1649977179
transform 1 0 8280 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_94
timestamp 1649977179
transform 1 0 9752 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_106
timestamp 1649977179
transform 1 0 10856 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1649977179
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1649977179
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1649977179
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_13
timestamp 1649977179
transform 1 0 2300 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_25
timestamp 1649977179
transform 1 0 3404 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_34
timestamp 1649977179
transform 1 0 4232 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_42
timestamp 1649977179
transform 1 0 4968 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_46
timestamp 1649977179
transform 1 0 5336 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_49
timestamp 1649977179
transform 1 0 5612 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_68
timestamp 1649977179
transform 1 0 7360 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_80
timestamp 1649977179
transform 1 0 8464 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_88
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_107
timestamp 1649977179
transform 1 0 10948 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_142
timestamp 1649977179
transform 1 0 14168 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_150
timestamp 1649977179
transform 1 0 14904 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_176
timestamp 1649977179
transform 1 0 17296 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_196
timestamp 1649977179
transform 1 0 19136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_216
timestamp 1649977179
transform 1 0 20976 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_222
timestamp 1649977179
transform 1 0 21528 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_11
timestamp 1649977179
transform 1 0 2116 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1649977179
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_44
timestamp 1649977179
transform 1 0 5152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_48
timestamp 1649977179
transform 1 0 5520 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_58
timestamp 1649977179
transform 1 0 6440 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_66
timestamp 1649977179
transform 1 0 7176 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_78
timestamp 1649977179
transform 1 0 8280 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_146
timestamp 1649977179
transform 1 0 14536 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_188
timestamp 1649977179
transform 1 0 18400 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_13
timestamp 1649977179
transform 1 0 2300 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_21
timestamp 1649977179
transform 1 0 3036 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_25
timestamp 1649977179
transform 1 0 3404 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_33
timestamp 1649977179
transform 1 0 4140 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_37
timestamp 1649977179
transform 1 0 4508 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_80
timestamp 1649977179
transform 1 0 8464 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_90
timestamp 1649977179
transform 1 0 9384 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_121
timestamp 1649977179
transform 1 0 12236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_160
timestamp 1649977179
transform 1 0 15824 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_216
timestamp 1649977179
transform 1 0 20976 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_222
timestamp 1649977179
transform 1 0 21528 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1649977179
transform 1 0 1748 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_11
timestamp 1649977179
transform 1 0 2116 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_23
timestamp 1649977179
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_40
timestamp 1649977179
transform 1 0 4784 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_52
timestamp 1649977179
transform 1 0 5888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_89
timestamp 1649977179
transform 1 0 9292 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_117
timestamp 1649977179
transform 1 0 11868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_123
timestamp 1649977179
transform 1 0 12420 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_143
timestamp 1649977179
transform 1 0 14260 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_155
timestamp 1649977179
transform 1 0 15364 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_199
timestamp 1649977179
transform 1 0 19412 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_203
timestamp 1649977179
transform 1 0 19780 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_220
timestamp 1649977179
transform 1 0 21344 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_7
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_19
timestamp 1649977179
transform 1 0 2852 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_31
timestamp 1649977179
transform 1 0 3956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_66
timestamp 1649977179
transform 1 0 7176 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_76
timestamp 1649977179
transform 1 0 8096 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_84
timestamp 1649977179
transform 1 0 8832 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_139
timestamp 1649977179
transform 1 0 13892 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_203
timestamp 1649977179
transform 1 0 19780 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_19
timestamp 1649977179
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_50
timestamp 1649977179
transform 1 0 5704 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_61
timestamp 1649977179
transform 1 0 6716 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_67
timestamp 1649977179
transform 1 0 7268 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1649977179
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_105
timestamp 1649977179
transform 1 0 10764 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_117
timestamp 1649977179
transform 1 0 11868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1649977179
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_163
timestamp 1649977179
transform 1 0 16100 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_182
timestamp 1649977179
transform 1 0 17848 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_187
timestamp 1649977179
transform 1 0 18308 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_201
timestamp 1649977179
transform 1 0 19596 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_220
timestamp 1649977179
transform 1 0 21344 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_14
timestamp 1649977179
transform 1 0 2392 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_19
timestamp 1649977179
transform 1 0 2852 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_50
timestamp 1649977179
transform 1 0 5704 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_70
timestamp 1649977179
transform 1 0 7544 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_100
timestamp 1649977179
transform 1 0 10304 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_157
timestamp 1649977179
transform 1 0 15548 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1649977179
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_222
timestamp 1649977179
transform 1 0 21528 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_11
timestamp 1649977179
transform 1 0 2116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_18
timestamp 1649977179
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1649977179
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_31
timestamp 1649977179
transform 1 0 3956 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_35
timestamp 1649977179
transform 1 0 4324 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_63
timestamp 1649977179
transform 1 0 6900 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1649977179
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_98
timestamp 1649977179
transform 1 0 10120 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_108
timestamp 1649977179
transform 1 0 11040 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_116
timestamp 1649977179
transform 1 0 11776 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_161
timestamp 1649977179
transform 1 0 15916 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_183
timestamp 1649977179
transform 1 0 17940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_7
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_19
timestamp 1649977179
transform 1 0 2852 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_23
timestamp 1649977179
transform 1 0 3220 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_28
timestamp 1649977179
transform 1 0 3680 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_40
timestamp 1649977179
transform 1 0 4784 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_68
timestamp 1649977179
transform 1 0 7360 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_80
timestamp 1649977179
transform 1 0 8464 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_85
timestamp 1649977179
transform 1 0 8924 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_95
timestamp 1649977179
transform 1 0 9844 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_116
timestamp 1649977179
transform 1 0 11776 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_158
timestamp 1649977179
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_201
timestamp 1649977179
transform 1 0 19596 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_222
timestamp 1649977179
transform 1 0 21528 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_11
timestamp 1649977179
transform 1 0 2116 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_19
timestamp 1649977179
transform 1 0 2852 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1649977179
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_40
timestamp 1649977179
transform 1 0 4784 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_57
timestamp 1649977179
transform 1 0 6348 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_61
timestamp 1649977179
transform 1 0 6716 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_112
timestamp 1649977179
transform 1 0 11408 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_116
timestamp 1649977179
transform 1 0 11776 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1649977179
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_164
timestamp 1649977179
transform 1 0 16192 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_170
timestamp 1649977179
transform 1 0 16744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_190
timestamp 1649977179
transform 1 0 18584 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_215
timestamp 1649977179
transform 1 0 20884 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_7
timestamp 1649977179
transform 1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_14
timestamp 1649977179
transform 1 0 2392 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_22
timestamp 1649977179
transform 1 0 3128 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_29
timestamp 1649977179
transform 1 0 3772 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_42
timestamp 1649977179
transform 1 0 4968 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1649977179
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_79
timestamp 1649977179
transform 1 0 8372 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_103
timestamp 1649977179
transform 1 0 10580 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_147
timestamp 1649977179
transform 1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_151
timestamp 1649977179
transform 1 0 14996 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_187
timestamp 1649977179
transform 1 0 18308 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_212
timestamp 1649977179
transform 1 0 20608 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_218
timestamp 1649977179
transform 1 0 21160 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1649977179
transform 1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1649977179
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_61
timestamp 1649977179
transform 1 0 6716 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1649977179
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_96
timestamp 1649977179
transform 1 0 9936 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_108
timestamp 1649977179
transform 1 0 11040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_114
timestamp 1649977179
transform 1 0 11592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1649977179
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_187
timestamp 1649977179
transform 1 0 18308 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_14
timestamp 1649977179
transform 1 0 2392 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_26
timestamp 1649977179
transform 1 0 3496 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_38
timestamp 1649977179
transform 1 0 4600 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1649977179
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_61
timestamp 1649977179
transform 1 0 6716 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_86
timestamp 1649977179
transform 1 0 9016 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_99
timestamp 1649977179
transform 1 0 10212 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_108
timestamp 1649977179
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_129
timestamp 1649977179
transform 1 0 12972 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_148
timestamp 1649977179
transform 1 0 14720 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_12
timestamp 1649977179
transform 1 0 2208 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1649977179
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_72
timestamp 1649977179
transform 1 0 7728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_88
timestamp 1649977179
transform 1 0 9200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_134
timestamp 1649977179
transform 1 0 13432 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_147
timestamp 1649977179
transform 1 0 14628 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_166
timestamp 1649977179
transform 1 0 16376 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_222
timestamp 1649977179
transform 1 0 21528 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_19
timestamp 1649977179
transform 1 0 2852 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_31
timestamp 1649977179
transform 1 0 3956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_43
timestamp 1649977179
transform 1 0 5060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_59
timestamp 1649977179
transform 1 0 6532 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_98
timestamp 1649977179
transform 1 0 10120 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_109
timestamp 1649977179
transform 1 0 11132 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_139
timestamp 1649977179
transform 1 0 13892 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_151
timestamp 1649977179
transform 1 0 14996 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1649977179
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_222
timestamp 1649977179
transform 1 0 21528 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1649977179
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_31
timestamp 1649977179
transform 1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_35
timestamp 1649977179
transform 1 0 4324 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_38
timestamp 1649977179
transform 1 0 4600 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_49
timestamp 1649977179
transform 1 0 5612 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_66
timestamp 1649977179
transform 1 0 7176 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_80
timestamp 1649977179
transform 1 0 8464 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_89
timestamp 1649977179
transform 1 0 9292 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_151
timestamp 1649977179
transform 1 0 14996 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_168
timestamp 1649977179
transform 1 0 16560 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_180
timestamp 1649977179
transform 1 0 17664 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_188
timestamp 1649977179
transform 1 0 18400 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_24
timestamp 1649977179
transform 1 0 3312 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_29
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_139
timestamp 1649977179
transform 1 0 13892 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1649977179
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_185
timestamp 1649977179
transform 1 0 18124 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_190
timestamp 1649977179
transform 1 0 18584 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_195
timestamp 1649977179
transform 1 0 19044 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_197
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1649977179
transform 1 0 21528 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _066_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1649977179
transform 1 0 2116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1649977179
transform 1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1649977179
transform 1 0 1840 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1649977179
transform 1 0 1564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1649977179
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1649977179
transform 1 0 1840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1649977179
transform 1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1649977179
transform 1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1649977179
transform 1 0 2208 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1649977179
transform 1 0 2576 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1649977179
transform 1 0 2392 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1649977179
transform 1 0 2852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1649977179
transform 1 0 3496 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1649977179
transform 1 0 2576 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform 1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1649977179
transform 1 0 2116 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1649977179
transform 1 0 2668 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1649977179
transform 1 0 13248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1649977179
transform -1 0 13800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1649977179
transform -1 0 14628 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1649977179
transform -1 0 14352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1649977179
transform -1 0 15180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1649977179
transform -1 0 12512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1649977179
transform -1 0 14904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1649977179
transform -1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1649977179
transform -1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1649977179
transform -1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform 1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1649977179
transform 1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1649977179
transform 1 0 20516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1649977179
transform 1 0 20148 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1649977179
transform -1 0 15916 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1649977179
transform -1 0 16376 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1649977179
transform -1 0 20148 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1649977179
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1649977179
transform -1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1649977179
transform -1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1649977179
transform -1 0 10764 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1649977179
transform -1 0 9660 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1649977179
transform -1 0 9568 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1649977179
transform -1 0 7820 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1649977179
transform -1 0 10028 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1649977179
transform -1 0 7452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1649977179
transform -1 0 7544 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1649977179
transform -1 0 8832 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1649977179
transform -1 0 9200 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1649977179
transform -1 0 9752 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1649977179
transform -1 0 10120 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1649977179
transform -1 0 10488 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1649977179
transform -1 0 8648 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1649977179
transform -1 0 14628 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1649977179
transform -1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1649977179
transform -1 0 8372 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1649977179
transform -1 0 9844 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1649977179
transform -1 0 9292 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1649977179
transform -1 0 14352 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1649977179
transform -1 0 16560 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 16008 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 3220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 2392 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 2944 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 3496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform 1 0 21344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 21344 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 1932 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 1932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 1932 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 1932 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform -1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform -1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform -1 0 1932 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform -1 0 4416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input32 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform -1 0 8464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1649977179
transform 1 0 9016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10120 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1649977179
transform -1 0 11408 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 10488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1649977179
transform -1 0 12420 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1649977179
transform 1 0 12420 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform -1 0 13984 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform -1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1649977179
transform 1 0 5060 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform -1 0 5336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1649977179
transform -1 0 6256 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1649977179
transform 1 0 6440 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1649977179
transform 1 0 6900 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1649977179
transform -1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1649977179
transform 1 0 7820 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1649977179
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform -1 0 4140 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform -1 0 9200 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1649977179
transform 1 0 9200 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1649977179
transform -1 0 10580 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1649977179
transform -1 0 10488 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform 1 0 10856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1649977179
transform -1 0 11500 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1649977179
transform -1 0 11408 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp 1649977179
transform -1 0 13892 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1649977179
transform 1 0 13524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1649977179
transform -1 0 4416 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 1649977179
transform -1 0 5336 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1649977179
transform -1 0 5612 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1649977179
transform -1 0 6256 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1649977179
transform 1 0 6256 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1649977179
transform 1 0 6716 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1649977179
transform -1 0 6716 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1649977179
transform 1 0 7636 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1649977179
transform 1 0 8096 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1649977179
transform -1 0 2300 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input72
timestamp 1649977179
transform -1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1649977179
transform 1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1649977179
transform -1 0 2300 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1649977179
transform -1 0 2300 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1649977179
transform -1 0 2300 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1649977179
transform -1 0 2024 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1649977179
transform -1 0 2024 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1649977179
transform -1 0 2668 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1649977179
transform -1 0 2392 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1649977179
transform -1 0 2852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1649977179
transform -1 0 3312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1649977179
transform -1 0 3680 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input87
timestamp 1649977179
transform 1 0 19504 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21252 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12052 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15272 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11500 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15732 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13800 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13708 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 10120 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14168 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13156 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 17112 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19320 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21160 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18124 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 -1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20884 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21344 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20792 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17112 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 18124 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21344 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15916 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18400 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13340 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12236 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13524 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14168 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12512 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15640 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13984 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12512 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14168 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17480 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19136 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20792 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18124 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18400 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21068 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16560 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 20148 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21620 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 20976 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16744 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13432 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12512 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12972 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17572 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21160 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19780 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19596 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17664 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18952 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20976 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19780 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21620 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16560 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14536 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14720 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21068 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19320 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21528 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17756 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15824 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 12972 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13616 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13156 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16560 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11868 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 16468 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19596 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18308 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 20700 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19412 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13616 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14996 0 -1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15272 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17572 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15364 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16744 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10580 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8464 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10488 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 9016 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1649977179
transform -1 0 6440 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_1.mux_l2_in_3__175 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1649977179
transform -1 0 5888 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform -1 0 11040 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1649977179
transform -1 0 7176 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1649977179
transform -1 0 12420 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13524 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9108 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5980 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1649977179
transform -1 0 2484 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_3.mux_l2_in_3__178
timestamp 1649977179
transform 1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1649977179
transform -1 0 2668 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1649977179
transform -1 0 5704 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1649977179
transform -1 0 11408 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12420 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10120 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 7360 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_4_
timestamp 1649977179
transform 1 0 4232 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_5_
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_6_
timestamp 1649977179
transform -1 0 2576 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11408 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7176 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1649977179
transform -1 0 4876 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_5.mux_l2_in_3__180
timestamp 1649977179
transform 1 0 5888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1649977179
transform -1 0 6256 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 12236 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1649977179
transform -1 0 9752 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1649977179
transform -1 0 13800 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 14076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15456 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8188 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1649977179
transform -1 0 4692 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_9.mux_l2_in_3__181
timestamp 1649977179
transform 1 0 5704 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1649977179
transform -1 0 4876 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14996 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1649977179
transform -1 0 10488 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 14352 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 14628 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13248 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1649977179
transform -1 0 8556 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1649977179
transform -1 0 5336 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_17.mux_l1_in_3__176
timestamp 1649977179
transform 1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_3_
timestamp 1649977179
transform -1 0 4876 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13340 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1649977179
transform -1 0 10488 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1649977179
transform -1 0 14720 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16100 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17572 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10212 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1649977179
transform -1 0 11868 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18124 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1649977179
transform -1 0 18216 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_25.mux_l2_in_1__177
timestamp 1649977179
transform -1 0 17296 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1649977179
transform -1 0 20792 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20608 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10212 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1649977179
transform -1 0 5152 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1649977179
transform -1 0 5428 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11224 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12236 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_33.mux_l2_in_1__179
timestamp 1649977179
transform 1 0 11868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1649977179
transform -1 0 17388 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19044 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5612 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_1.mux_l1_in_3__182
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1649977179
transform -1 0 6256 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5428 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5612 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6256 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6440 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6440 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_3.mux_l1_in_3__159
timestamp 1649977179
transform 1 0 7268 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1649977179
transform 1 0 6440 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 6256 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6164 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7268 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7912 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8740 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_5.mux_l1_in_3__165
timestamp 1649977179
transform -1 0 8004 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1649977179
transform 1 0 7912 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7084 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6900 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2668 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8464 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9292 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_7.mux_l1_in_3__166
timestamp 1649977179
transform 1 0 9384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_3_
timestamp 1649977179
transform -1 0 8556 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7820 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7820 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6992 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3036 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12236 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10120 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_9.mux_l2_in_1__167
timestamp 1649977179
transform 1 0 11316 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10488 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9752 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15088 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9108 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_11.mux_l2_in_1__183
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10488 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9108 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16008 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1649977179
transform -1 0 12604 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_13.mux_l2_in_1__184
timestamp 1649977179
transform 1 0 12880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12052 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11868 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 5428 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17848 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_15.mux_l2_in_1__185
timestamp 1649977179
transform -1 0 14352 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14260 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l3_in_0_
timestamp 1649977179
transform 1 0 13432 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6072 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9108 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_17.mux_l1_in_1__153
timestamp 1649977179
transform 1 0 9752 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1649977179
transform -1 0 9752 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_19.mux_l1_in_1__154
timestamp 1649977179
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_1_
timestamp 1649977179
transform -1 0 9108 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4232 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10212 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_21.mux_l1_in_1__155
timestamp 1649977179
transform 1 0 9752 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4508 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10120 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_23.mux_l1_in_1__156
timestamp 1649977179
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10304 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9292 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9936 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_25.mux_l1_in_1__157
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10488 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9660 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4784 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10580 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_29.mux_l2_in_0__158
timestamp 1649977179
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10212 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3404 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11132 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10396 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_31.mux_l2_in_0__160
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3496 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9568 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_33.mux_l2_in_0__161
timestamp 1649977179
transform 1 0 9476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8740 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7820 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_35.mux_l2_in_0__162
timestamp 1649977179
transform -1 0 7084 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2944 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6072 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5520 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_37.mux_l2_in_0__163
timestamp 1649977179
transform -1 0 5336 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2944 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8188 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_39.mux_l2_in_0__164
timestamp 1649977179
transform 1 0 7912 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8372 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7820 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6072 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1649977179
transform -1 0 5244 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1649977179
transform -1 0 8740 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6164 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1649977179
transform -1 0 6164 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_0.mux_l2_in_3__168
timestamp 1649977179
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1649977179
transform -1 0 5980 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8280 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 7084 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 8464 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9752 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4692 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5428 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1649977179
transform -1 0 8280 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_2.mux_l2_in_3__170
timestamp 1649977179
transform 1 0 9936 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6716 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1649977179
transform -1 0 8464 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1649977179
transform 1 0 9476 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9476 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5888 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1649977179
transform -1 0 4784 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5152 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1649977179
transform -1 0 4968 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_4_
timestamp 1649977179
transform 1 0 7544 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_5_
timestamp 1649977179
transform 1 0 7452 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_6_
timestamp 1649977179
transform -1 0 5152 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5980 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5888 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 7268 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_4.mux_l2_in_3__173
timestamp 1649977179
transform 1 0 5428 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1649977179
transform -1 0 5796 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 7452 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1649977179
transform -1 0 7544 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9752 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7360 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9476 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 10396 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1649977179
transform -1 0 5336 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_8.mux_l2_in_3__174
timestamp 1649977179
transform 1 0 5060 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1649977179
transform -1 0 5428 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9936 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1649977179
transform -1 0 7176 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1649977179
transform -1 0 9936 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9844 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4600 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10948 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1649977179
transform -1 0 3036 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_16.mux_l1_in_3__169
timestamp 1649977179
transform 1 0 2852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_3_
timestamp 1649977179
transform -1 0 3220 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10212 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7176 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9936 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9292 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3772 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1649977179
transform -1 0 2668 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_24.mux_l1_in_3__171
timestamp 1649977179
transform -1 0 3680 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_3_
timestamp 1649977179
transform -1 0 4600 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11040 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7268 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9384 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9016 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5704 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7268 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1649977179
transform -1 0 7176 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8004 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_32.mux_l2_in_1__172
timestamp 1649977179
transform -1 0 7636 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8464 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9292 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output88 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform -1 0 2116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform -1 0 2116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform -1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform -1 0 2116 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 2484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform -1 0 2116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform -1 0 2116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1649977179
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform 1 0 13340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1649977179
transform -1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1649977179
transform -1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1649977179
transform -1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1649977179
transform -1 0 19964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1649977179
transform 1 0 19964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1649977179
transform 1 0 21160 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1649977179
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1649977179
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform 1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1649977179
transform 1 0 15640 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1649977179
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1649977179
transform -1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1649977179
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1649977179
transform 1 0 13156 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1649977179
transform 1 0 18216 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1649977179
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1649977179
transform 1 0 19596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1649977179
transform 1 0 20792 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1649977179
transform 1 0 21160 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1649977179
transform 1 0 20976 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1649977179
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1649977179
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1649977179
transform 1 0 14444 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1649977179
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1649977179
transform 1 0 17020 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1649977179
transform 1 0 17388 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20424 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  repeater149
timestamp 1649977179
transform -1 0 6716 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater150
timestamp 1649977179
transform -1 0 11868 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater151
timestamp 1649977179
transform -1 0 11408 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater152
timestamp 1649977179
transform -1 0 13340 0 -1 10880
box -38 -48 406 592
<< labels >>
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 386 0 442 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_42_
port 2 nsew signal input
flabel metal2 s 846 0 902 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_43_
port 3 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_44_
port 4 nsew signal input
flabel metal2 s 1766 0 1822 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_45_
port 5 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_46_
port 6 nsew signal input
flabel metal2 s 2686 0 2742 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_47_
port 7 nsew signal input
flabel metal2 s 3146 0 3202 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_48_
port 8 nsew signal input
flabel metal2 s 3606 0 3662 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_49_
port 9 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 bottom_right_grid_pin_1_
port 10 nsew signal input
flabel metal3 s 22200 5720 23000 5840 0 FreeSans 480 0 0 0 ccff_head
port 11 nsew signal input
flabel metal3 s 22200 17144 23000 17264 0 FreeSans 480 0 0 0 ccff_tail
port 12 nsew signal tristate
flabel metal3 s 0 5040 800 5160 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 13 nsew signal input
flabel metal3 s 0 9120 800 9240 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 14 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 15 nsew signal input
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 16 nsew signal input
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 17 nsew signal input
flabel metal3 s 0 10752 800 10872 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 18 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 19 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 20 nsew signal input
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 21 nsew signal input
flabel metal3 s 0 12384 800 12504 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 22 nsew signal input
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 23 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 24 nsew signal input
flabel metal3 s 0 5856 800 5976 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 25 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 26 nsew signal input
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 27 nsew signal input
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 28 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 29 nsew signal input
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 30 nsew signal input
flabel metal3 s 0 8304 800 8424 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 31 nsew signal input
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 32 nsew signal input
flabel metal3 s 0 13200 800 13320 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 33 nsew signal tristate
flabel metal3 s 0 17280 800 17400 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 34 nsew signal tristate
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 35 nsew signal tristate
flabel metal3 s 0 18096 800 18216 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 36 nsew signal tristate
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 37 nsew signal tristate
flabel metal3 s 0 18912 800 19032 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 38 nsew signal tristate
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 39 nsew signal tristate
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 40 nsew signal tristate
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 41 nsew signal tristate
flabel metal3 s 0 20544 800 20664 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 42 nsew signal tristate
flabel metal3 s 0 20952 800 21072 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 43 nsew signal tristate
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 44 nsew signal tristate
flabel metal3 s 0 14016 800 14136 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 45 nsew signal tristate
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 46 nsew signal tristate
flabel metal3 s 0 14832 800 14952 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 47 nsew signal tristate
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 48 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 49 nsew signal tristate
flabel metal3 s 0 16056 800 16176 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 50 nsew signal tristate
flabel metal3 s 0 16464 800 16584 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 51 nsew signal tristate
flabel metal3 s 0 16872 800 16992 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 52 nsew signal tristate
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 53 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 54 nsew signal input
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 55 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 56 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 57 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 58 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 59 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 60 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 61 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 62 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 63 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 64 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 65 nsew signal input
flabel metal2 s 5446 0 5502 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 66 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 67 nsew signal input
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 68 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 69 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 70 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 71 nsew signal input
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 72 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 73 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 74 nsew signal tristate
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 75 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 76 nsew signal tristate
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 77 nsew signal tristate
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 78 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 79 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 80 nsew signal tristate
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 81 nsew signal tristate
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 82 nsew signal tristate
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 83 nsew signal tristate
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 84 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 85 nsew signal tristate
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 86 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 87 nsew signal tristate
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 88 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 89 nsew signal tristate
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 90 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 91 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 92 nsew signal tristate
flabel metal2 s 3882 22200 3938 23000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 93 nsew signal input
flabel metal2 s 8482 22200 8538 23000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 94 nsew signal input
flabel metal2 s 8942 22200 8998 23000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 95 nsew signal input
flabel metal2 s 9402 22200 9458 23000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 96 nsew signal input
flabel metal2 s 9862 22200 9918 23000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 97 nsew signal input
flabel metal2 s 10322 22200 10378 23000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 98 nsew signal input
flabel metal2 s 10782 22200 10838 23000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 99 nsew signal input
flabel metal2 s 11242 22200 11298 23000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 100 nsew signal input
flabel metal2 s 11702 22200 11758 23000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 101 nsew signal input
flabel metal2 s 12162 22200 12218 23000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 102 nsew signal input
flabel metal2 s 12622 22200 12678 23000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 103 nsew signal input
flabel metal2 s 4342 22200 4398 23000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 104 nsew signal input
flabel metal2 s 4802 22200 4858 23000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 105 nsew signal input
flabel metal2 s 5262 22200 5318 23000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 106 nsew signal input
flabel metal2 s 5722 22200 5778 23000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 107 nsew signal input
flabel metal2 s 6182 22200 6238 23000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 108 nsew signal input
flabel metal2 s 6642 22200 6698 23000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 109 nsew signal input
flabel metal2 s 7102 22200 7158 23000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 110 nsew signal input
flabel metal2 s 7562 22200 7618 23000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 111 nsew signal input
flabel metal2 s 8022 22200 8078 23000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 112 nsew signal input
flabel metal2 s 13082 22200 13138 23000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 113 nsew signal tristate
flabel metal2 s 17682 22200 17738 23000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 114 nsew signal tristate
flabel metal2 s 18142 22200 18198 23000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 115 nsew signal tristate
flabel metal2 s 18602 22200 18658 23000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 116 nsew signal tristate
flabel metal2 s 19062 22200 19118 23000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 117 nsew signal tristate
flabel metal2 s 19522 22200 19578 23000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 118 nsew signal tristate
flabel metal2 s 19982 22200 20038 23000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 119 nsew signal tristate
flabel metal2 s 20442 22200 20498 23000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 120 nsew signal tristate
flabel metal2 s 20902 22200 20958 23000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 121 nsew signal tristate
flabel metal2 s 21362 22200 21418 23000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 122 nsew signal tristate
flabel metal2 s 21822 22200 21878 23000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 123 nsew signal tristate
flabel metal2 s 13542 22200 13598 23000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 124 nsew signal tristate
flabel metal2 s 14002 22200 14058 23000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 125 nsew signal tristate
flabel metal2 s 14462 22200 14518 23000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 126 nsew signal tristate
flabel metal2 s 14922 22200 14978 23000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 127 nsew signal tristate
flabel metal2 s 15382 22200 15438 23000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 128 nsew signal tristate
flabel metal2 s 15842 22200 15898 23000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 129 nsew signal tristate
flabel metal2 s 16302 22200 16358 23000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 130 nsew signal tristate
flabel metal2 s 16762 22200 16818 23000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 131 nsew signal tristate
flabel metal2 s 17222 22200 17278 23000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 132 nsew signal tristate
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 left_bottom_grid_pin_34_
port 133 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 left_bottom_grid_pin_35_
port 134 nsew signal input
flabel metal3 s 0 2592 800 2712 0 FreeSans 480 0 0 0 left_bottom_grid_pin_36_
port 135 nsew signal input
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 left_bottom_grid_pin_37_
port 136 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 left_bottom_grid_pin_38_
port 137 nsew signal input
flabel metal3 s 0 3816 800 3936 0 FreeSans 480 0 0 0 left_bottom_grid_pin_39_
port 138 nsew signal input
flabel metal3 s 0 4224 800 4344 0 FreeSans 480 0 0 0 left_bottom_grid_pin_40_
port 139 nsew signal input
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 left_bottom_grid_pin_41_
port 140 nsew signal input
flabel metal2 s 22282 22200 22338 23000 0 FreeSans 224 90 0 0 prog_clk_0_N_in
port 141 nsew signal input
flabel metal2 s 202 22200 258 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_42_
port 142 nsew signal input
flabel metal2 s 662 22200 718 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_43_
port 143 nsew signal input
flabel metal2 s 1122 22200 1178 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_44_
port 144 nsew signal input
flabel metal2 s 1582 22200 1638 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_45_
port 145 nsew signal input
flabel metal2 s 2042 22200 2098 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_46_
port 146 nsew signal input
flabel metal2 s 2502 22200 2558 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_47_
port 147 nsew signal input
flabel metal2 s 2962 22200 3018 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_48_
port 148 nsew signal input
flabel metal2 s 3422 22200 3478 23000 0 FreeSans 224 90 0 0 top_left_grid_pin_49_
port 149 nsew signal input
flabel metal2 s 22742 22200 22798 23000 0 FreeSans 224 90 0 0 top_right_grid_pin_1_
port 150 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
