magic
tech sky130A
magscale 1 2
timestamp 1656241527
<< viali >>
rect 1593 17289 1627 17323
rect 1961 17289 1995 17323
rect 2329 17289 2363 17323
rect 2697 17289 2731 17323
rect 3065 17289 3099 17323
rect 3525 17289 3559 17323
rect 3985 17289 4019 17323
rect 4261 17289 4295 17323
rect 4537 17289 4571 17323
rect 4905 17289 4939 17323
rect 5641 17289 5675 17323
rect 6101 17289 6135 17323
rect 7297 17289 7331 17323
rect 7573 17289 7607 17323
rect 8033 17289 8067 17323
rect 8585 17289 8619 17323
rect 13461 17289 13495 17323
rect 13737 17289 13771 17323
rect 1777 17153 1811 17187
rect 2145 17153 2179 17187
rect 2513 17153 2547 17187
rect 2881 17153 2915 17187
rect 3249 17153 3283 17187
rect 3341 17153 3375 17187
rect 3801 17153 3835 17187
rect 4077 17153 4111 17187
rect 4721 17153 4755 17187
rect 5089 17153 5123 17187
rect 5457 17153 5491 17187
rect 5825 17153 5859 17187
rect 5917 17153 5951 17187
rect 6745 17153 6779 17187
rect 7113 17153 7147 17187
rect 7474 17153 7508 17187
rect 7941 17153 7975 17187
rect 8769 17153 8803 17187
rect 9321 17153 9355 17187
rect 9873 17153 9907 17187
rect 10609 17153 10643 17187
rect 11529 17153 11563 17187
rect 12449 17153 12483 17187
rect 13553 17153 13587 17187
rect 13921 17153 13955 17187
rect 14105 17153 14139 17187
rect 15117 17153 15151 17187
rect 8217 17085 8251 17119
rect 9597 17085 9631 17119
rect 9781 17085 9815 17119
rect 10333 17085 10367 17119
rect 11805 17085 11839 17119
rect 12725 17085 12759 17119
rect 14381 17085 14415 17119
rect 15301 17085 15335 17119
rect 5273 17017 5307 17051
rect 6561 17017 6595 17051
rect 6929 17017 6963 17051
rect 9045 16949 9079 16983
rect 9229 16949 9263 16983
rect 10241 16949 10275 16983
rect 11253 16949 11287 16983
rect 2605 16745 2639 16779
rect 2881 16745 2915 16779
rect 3341 16745 3375 16779
rect 5089 16745 5123 16779
rect 15301 16745 15335 16779
rect 1961 16677 1995 16711
rect 2421 16677 2455 16711
rect 3433 16677 3467 16711
rect 3985 16677 4019 16711
rect 4445 16677 4479 16711
rect 7757 16677 7791 16711
rect 8953 16677 8987 16711
rect 9229 16677 9263 16711
rect 11299 16677 11333 16711
rect 11989 16677 12023 16711
rect 6561 16609 6595 16643
rect 7297 16609 7331 16643
rect 8309 16609 8343 16643
rect 10149 16609 10183 16643
rect 10241 16609 10275 16643
rect 10701 16609 10735 16643
rect 11069 16609 11103 16643
rect 12725 16609 12759 16643
rect 13001 16609 13035 16643
rect 14657 16609 14691 16643
rect 1777 16541 1811 16575
rect 2145 16541 2179 16575
rect 2237 16541 2271 16575
rect 2789 16541 2823 16575
rect 3065 16541 3099 16575
rect 3157 16541 3191 16575
rect 3617 16541 3651 16575
rect 3801 16541 3835 16575
rect 4077 16541 4111 16575
rect 4629 16541 4663 16575
rect 4905 16541 4939 16575
rect 5181 16541 5215 16575
rect 5549 16541 5583 16575
rect 7113 16541 7147 16575
rect 7573 16541 7607 16575
rect 8585 16541 8619 16575
rect 9137 16541 9171 16575
rect 9413 16541 9447 16575
rect 13645 16541 13679 16575
rect 13921 16541 13955 16575
rect 14933 16541 14967 16575
rect 15025 16541 15059 16575
rect 6285 16473 6319 16507
rect 7205 16473 7239 16507
rect 10885 16473 10919 16507
rect 1593 16405 1627 16439
rect 4261 16405 4295 16439
rect 4813 16405 4847 16439
rect 5365 16405 5399 16439
rect 5733 16405 5767 16439
rect 5917 16405 5951 16439
rect 6377 16405 6411 16439
rect 6745 16405 6779 16439
rect 8125 16405 8159 16439
rect 8217 16405 8251 16439
rect 8769 16405 8803 16439
rect 9689 16405 9723 16439
rect 10057 16405 10091 16439
rect 10609 16405 10643 16439
rect 15485 16405 15519 16439
rect 2145 16201 2179 16235
rect 2421 16201 2455 16235
rect 2973 16201 3007 16235
rect 3709 16201 3743 16235
rect 4261 16201 4295 16235
rect 4905 16201 4939 16235
rect 5365 16201 5399 16235
rect 6837 16201 6871 16235
rect 7757 16201 7791 16235
rect 9045 16201 9079 16235
rect 9413 16201 9447 16235
rect 9505 16201 9539 16235
rect 9965 16201 9999 16235
rect 11529 16201 11563 16235
rect 11989 16201 12023 16235
rect 13553 16201 13587 16235
rect 4169 16133 4203 16167
rect 6745 16133 6779 16167
rect 10977 16133 11011 16167
rect 11897 16133 11931 16167
rect 13369 16133 13403 16167
rect 15669 16133 15703 16167
rect 1685 16065 1719 16099
rect 2053 16065 2087 16099
rect 2329 16065 2363 16099
rect 2605 16065 2639 16099
rect 2789 16065 2823 16099
rect 3525 16065 3559 16099
rect 4445 16065 4479 16099
rect 5733 16065 5767 16099
rect 5825 16065 5859 16099
rect 7205 16065 7239 16099
rect 7849 16065 7883 16099
rect 8677 16065 8711 16099
rect 10333 16065 10367 16099
rect 11069 16065 11103 16099
rect 12725 16065 12759 16099
rect 13737 16065 13771 16099
rect 3985 15997 4019 16031
rect 4997 15997 5031 16031
rect 5181 15997 5215 16031
rect 6009 15997 6043 16031
rect 6929 15997 6963 16031
rect 7665 15997 7699 16031
rect 8493 15997 8527 16031
rect 8585 15997 8619 16031
rect 9321 15997 9355 16031
rect 10425 15997 10459 16031
rect 10609 15997 10643 16031
rect 12081 15997 12115 16031
rect 12817 15997 12851 16031
rect 12909 15997 12943 16031
rect 13829 15997 13863 16031
rect 14013 15997 14047 16031
rect 1869 15929 1903 15963
rect 3341 15929 3375 15963
rect 6377 15929 6411 15963
rect 8217 15929 8251 15963
rect 13185 15929 13219 15963
rect 1501 15861 1535 15895
rect 3249 15861 3283 15895
rect 4537 15861 4571 15895
rect 7389 15861 7423 15895
rect 9873 15861 9907 15895
rect 11253 15861 11287 15895
rect 12357 15861 12391 15895
rect 1409 15657 1443 15691
rect 1777 15657 1811 15691
rect 2513 15657 2547 15691
rect 3433 15657 3467 15691
rect 4997 15657 5031 15691
rect 5457 15657 5491 15691
rect 5825 15657 5859 15691
rect 6377 15657 6411 15691
rect 8953 15657 8987 15691
rect 10241 15657 10275 15691
rect 12633 15657 12667 15691
rect 4169 15589 4203 15623
rect 7941 15589 7975 15623
rect 8033 15589 8067 15623
rect 13737 15589 13771 15623
rect 4813 15521 4847 15555
rect 5733 15521 5767 15555
rect 6285 15521 6319 15555
rect 6929 15521 6963 15555
rect 7389 15521 7423 15555
rect 8493 15521 8527 15555
rect 8585 15521 8619 15555
rect 9505 15521 9539 15555
rect 10793 15521 10827 15555
rect 11529 15521 11563 15555
rect 11621 15521 11655 15555
rect 11989 15521 12023 15555
rect 13001 15521 13035 15555
rect 14841 15521 14875 15555
rect 1593 15453 1627 15487
rect 1869 15453 1903 15487
rect 2697 15453 2731 15487
rect 2973 15453 3007 15487
rect 3617 15453 3651 15487
rect 4537 15453 4571 15487
rect 5181 15453 5215 15487
rect 6009 15453 6043 15487
rect 6745 15453 6779 15487
rect 9321 15453 9355 15487
rect 9781 15453 9815 15487
rect 10057 15453 10091 15487
rect 10701 15453 10735 15487
rect 12265 15453 12299 15487
rect 13921 15453 13955 15487
rect 14657 15453 14691 15487
rect 15117 15453 15151 15487
rect 7573 15385 7607 15419
rect 13185 15385 13219 15419
rect 13277 15385 13311 15419
rect 14289 15385 14323 15419
rect 2053 15317 2087 15351
rect 2145 15317 2179 15351
rect 2421 15317 2455 15351
rect 3065 15317 3099 15351
rect 3341 15317 3375 15351
rect 3801 15317 3835 15351
rect 4629 15317 4663 15351
rect 6837 15317 6871 15351
rect 7481 15317 7515 15351
rect 8401 15317 8435 15351
rect 9413 15317 9447 15351
rect 9965 15317 9999 15351
rect 10609 15317 10643 15351
rect 11069 15317 11103 15351
rect 11437 15317 11471 15351
rect 12173 15317 12207 15351
rect 12817 15317 12851 15351
rect 13645 15317 13679 15351
rect 14197 15317 14231 15351
rect 14565 15317 14599 15351
rect 3065 15113 3099 15147
rect 3525 15113 3559 15147
rect 4169 15113 4203 15147
rect 4445 15113 4479 15147
rect 4905 15113 4939 15147
rect 5273 15113 5307 15147
rect 6377 15113 6411 15147
rect 6561 15113 6595 15147
rect 7021 15113 7055 15147
rect 7389 15113 7423 15147
rect 7757 15113 7791 15147
rect 8677 15113 8711 15147
rect 9873 15113 9907 15147
rect 9965 15113 9999 15147
rect 11345 15113 11379 15147
rect 11897 15113 11931 15147
rect 12357 15113 12391 15147
rect 13737 15113 13771 15147
rect 14105 15113 14139 15147
rect 15577 15113 15611 15147
rect 2513 15045 2547 15079
rect 5641 15045 5675 15079
rect 6193 15045 6227 15079
rect 10977 15045 11011 15079
rect 13185 15045 13219 15079
rect 14473 15045 14507 15079
rect 1685 14977 1719 15011
rect 1961 14977 1995 15011
rect 4077 14977 4111 15011
rect 4353 14977 4387 15011
rect 4813 14977 4847 15011
rect 6929 14977 6963 15011
rect 8401 14977 8435 15011
rect 9045 14977 9079 15011
rect 10885 14977 10919 15011
rect 12725 14977 12759 15011
rect 12817 14977 12851 15011
rect 14289 14977 14323 15011
rect 3617 14909 3651 14943
rect 3801 14909 3835 14943
rect 4997 14909 5031 14943
rect 5733 14909 5767 14943
rect 5917 14909 5951 14943
rect 7113 14909 7147 14943
rect 7849 14909 7883 14943
rect 8033 14909 8067 14943
rect 9137 14909 9171 14943
rect 9321 14909 9355 14943
rect 10149 14909 10183 14943
rect 10701 14909 10735 14943
rect 11621 14909 11655 14943
rect 11805 14909 11839 14943
rect 12909 14909 12943 14943
rect 13461 14909 13495 14943
rect 13645 14909 13679 14943
rect 14657 14909 14691 14943
rect 14933 14909 14967 14943
rect 2881 14841 2915 14875
rect 9505 14841 9539 14875
rect 12265 14841 12299 14875
rect 1501 14773 1535 14807
rect 1777 14773 1811 14807
rect 2605 14773 2639 14807
rect 3157 14773 3191 14807
rect 8217 14773 8251 14807
rect 8493 14773 8527 14807
rect 10425 14773 10459 14807
rect 1501 14569 1535 14603
rect 5089 14569 5123 14603
rect 5917 14569 5951 14603
rect 7021 14569 7055 14603
rect 7297 14569 7331 14603
rect 8401 14569 8435 14603
rect 9413 14569 9447 14603
rect 11713 14569 11747 14603
rect 13553 14569 13587 14603
rect 8125 14501 8159 14535
rect 8953 14501 8987 14535
rect 2973 14433 3007 14467
rect 4353 14433 4387 14467
rect 5549 14433 5583 14467
rect 5733 14433 5767 14467
rect 6469 14433 6503 14467
rect 7849 14433 7883 14467
rect 9229 14433 9263 14467
rect 9689 14433 9723 14467
rect 10241 14433 10275 14467
rect 11161 14433 11195 14467
rect 13277 14433 13311 14467
rect 14565 14433 14599 14467
rect 1685 14365 1719 14399
rect 3157 14365 3191 14399
rect 4629 14365 4663 14399
rect 5457 14365 5491 14399
rect 6285 14365 6319 14399
rect 7665 14365 7699 14399
rect 8309 14365 8343 14399
rect 8585 14365 8619 14399
rect 8769 14365 8803 14399
rect 9137 14341 9171 14375
rect 13185 14365 13219 14399
rect 13737 14365 13771 14399
rect 14841 14365 14875 14399
rect 15634 14365 15668 14399
rect 3065 14297 3099 14331
rect 4997 14297 5031 14331
rect 11345 14297 11379 14331
rect 12918 14297 12952 14331
rect 14381 14297 14415 14331
rect 3525 14229 3559 14263
rect 3801 14229 3835 14263
rect 4169 14229 4203 14263
rect 4261 14229 4295 14263
rect 4813 14229 4847 14263
rect 6377 14229 6411 14263
rect 6745 14229 6779 14263
rect 7205 14229 7239 14263
rect 7757 14229 7791 14263
rect 9781 14229 9815 14263
rect 9965 14229 9999 14263
rect 10425 14229 10459 14263
rect 10517 14229 10551 14263
rect 10885 14229 10919 14263
rect 11253 14229 11287 14263
rect 11805 14229 11839 14263
rect 13921 14229 13955 14263
rect 14289 14229 14323 14263
rect 15531 14229 15565 14263
rect 3617 14025 3651 14059
rect 4721 14025 4755 14059
rect 7757 14025 7791 14059
rect 8033 14025 8067 14059
rect 8493 14025 8527 14059
rect 8861 14025 8895 14059
rect 9321 14025 9355 14059
rect 9689 14025 9723 14059
rect 10149 14025 10183 14059
rect 10517 14025 10551 14059
rect 13737 14025 13771 14059
rect 3433 13957 3467 13991
rect 4261 13957 4295 13991
rect 6622 13957 6656 13991
rect 8401 13957 8435 13991
rect 10057 13957 10091 13991
rect 10977 13957 11011 13991
rect 13829 13957 13863 13991
rect 15485 13957 15519 13991
rect 1685 13889 1719 13923
rect 2697 13889 2731 13923
rect 3157 13889 3191 13923
rect 5834 13889 5868 13923
rect 6101 13889 6135 13923
rect 6377 13889 6411 13923
rect 9229 13889 9263 13923
rect 11529 13889 11563 13923
rect 11796 13889 11830 13923
rect 13369 13889 13403 13923
rect 2789 13821 2823 13855
rect 2973 13821 3007 13855
rect 4353 13821 4387 13855
rect 8309 13821 8343 13855
rect 9137 13821 9171 13855
rect 9873 13821 9907 13855
rect 10701 13821 10735 13855
rect 10885 13821 10919 13855
rect 13185 13821 13219 13855
rect 13277 13821 13311 13855
rect 15669 13821 15703 13855
rect 1501 13753 1535 13787
rect 2329 13685 2363 13719
rect 4537 13685 4571 13719
rect 11345 13685 11379 13719
rect 12909 13685 12943 13719
rect 5273 13481 5307 13515
rect 5641 13481 5675 13515
rect 8953 13481 8987 13515
rect 9137 13481 9171 13515
rect 9781 13481 9815 13515
rect 11253 13481 11287 13515
rect 12909 13481 12943 13515
rect 13093 13481 13127 13515
rect 13185 13481 13219 13515
rect 14933 13481 14967 13515
rect 1777 13413 1811 13447
rect 2881 13413 2915 13447
rect 9597 13413 9631 13447
rect 11345 13413 11379 13447
rect 2237 13345 2271 13379
rect 3433 13345 3467 13379
rect 9873 13345 9907 13379
rect 12725 13345 12759 13379
rect 13737 13345 13771 13379
rect 14657 13345 14691 13379
rect 15485 13345 15519 13379
rect 1685 13277 1719 13311
rect 1961 13277 1995 13311
rect 2421 13277 2455 13311
rect 3249 13277 3283 13311
rect 3893 13277 3927 13311
rect 5457 13277 5491 13311
rect 7021 13277 7055 13311
rect 7205 13277 7239 13311
rect 7389 13277 7423 13311
rect 7656 13277 7690 13311
rect 10140 13277 10174 13311
rect 14565 13277 14599 13311
rect 15393 13277 15427 13311
rect 3341 13209 3375 13243
rect 4138 13209 4172 13243
rect 6754 13209 6788 13243
rect 12480 13209 12514 13243
rect 13645 13209 13679 13243
rect 15301 13209 15335 13243
rect 1501 13141 1535 13175
rect 2329 13141 2363 13175
rect 2789 13141 2823 13175
rect 8769 13141 8803 13175
rect 9413 13141 9447 13175
rect 13553 13141 13587 13175
rect 14105 13141 14139 13175
rect 14473 13141 14507 13175
rect 2421 12937 2455 12971
rect 3341 12937 3375 12971
rect 6193 12937 6227 12971
rect 7205 12937 7239 12971
rect 8769 12937 8803 12971
rect 10517 12937 10551 12971
rect 10701 12937 10735 12971
rect 10885 12937 10919 12971
rect 13001 12937 13035 12971
rect 13277 12937 13311 12971
rect 13737 12937 13771 12971
rect 14289 12937 14323 12971
rect 14749 12937 14783 12971
rect 15393 12937 15427 12971
rect 5058 12869 5092 12903
rect 8953 12869 8987 12903
rect 11253 12869 11287 12903
rect 14657 12869 14691 12903
rect 2329 12801 2363 12835
rect 2789 12801 2823 12835
rect 2881 12801 2915 12835
rect 4454 12801 4488 12835
rect 7389 12801 7423 12835
rect 7645 12801 7679 12835
rect 10158 12801 10192 12835
rect 10425 12801 10459 12835
rect 11529 12801 11563 12835
rect 11785 12801 11819 12835
rect 13829 12801 13863 12835
rect 15209 12801 15243 12835
rect 15485 12801 15519 12835
rect 3065 12733 3099 12767
rect 4721 12733 4755 12767
rect 4813 12733 4847 12767
rect 11161 12733 11195 12767
rect 13553 12733 13587 12767
rect 14841 12733 14875 12767
rect 14197 12665 14231 12699
rect 15669 12665 15703 12699
rect 9045 12597 9079 12631
rect 12909 12597 12943 12631
rect 2881 12393 2915 12427
rect 6745 12393 6779 12427
rect 8953 12393 8987 12427
rect 10885 12393 10919 12427
rect 14105 12393 14139 12427
rect 15577 12393 15611 12427
rect 15485 12325 15519 12359
rect 1777 12257 1811 12291
rect 2789 12257 2823 12291
rect 3341 12257 3375 12291
rect 3525 12257 3559 12291
rect 12633 12257 12667 12291
rect 13369 12257 13403 12291
rect 13829 12257 13863 12291
rect 14565 12257 14599 12291
rect 14749 12257 14783 12291
rect 15301 12257 15335 12291
rect 2605 12189 2639 12223
rect 3893 12189 3927 12223
rect 4629 12189 4663 12223
rect 4997 12189 5031 12223
rect 5181 12189 5215 12223
rect 5457 12189 5491 12223
rect 6653 12189 6687 12223
rect 8125 12189 8159 12223
rect 10077 12189 10111 12223
rect 10333 12189 10367 12223
rect 11069 12189 11103 12223
rect 13277 12189 13311 12223
rect 7880 12121 7914 12155
rect 8769 12121 8803 12155
rect 12366 12121 12400 12155
rect 14473 12121 14507 12155
rect 14933 12121 14967 12155
rect 1869 12053 1903 12087
rect 1961 12053 1995 12087
rect 2329 12053 2363 12087
rect 3249 12053 3283 12087
rect 11253 12053 11287 12087
rect 12817 12053 12851 12087
rect 13185 12053 13219 12087
rect 13737 12053 13771 12087
rect 1501 11849 1535 11883
rect 2605 11849 2639 11883
rect 4077 11849 4111 11883
rect 9505 11849 9539 11883
rect 12725 11849 12759 11883
rect 13001 11849 13035 11883
rect 13185 11849 13219 11883
rect 13829 11849 13863 11883
rect 14381 11849 14415 11883
rect 14565 11849 14599 11883
rect 14749 11849 14783 11883
rect 15577 11849 15611 11883
rect 2513 11781 2547 11815
rect 5190 11781 5224 11815
rect 10640 11781 10674 11815
rect 12265 11781 12299 11815
rect 14933 11781 14967 11815
rect 15393 11781 15427 11815
rect 1685 11713 1719 11747
rect 1961 11713 1995 11747
rect 3341 11713 3375 11747
rect 3433 11713 3467 11747
rect 12357 11713 12391 11747
rect 13737 11713 13771 11747
rect 15209 11713 15243 11747
rect 2789 11645 2823 11679
rect 3525 11645 3559 11679
rect 5457 11645 5491 11679
rect 10885 11645 10919 11679
rect 12449 11645 12483 11679
rect 14013 11645 14047 11679
rect 1777 11577 1811 11611
rect 2145 11509 2179 11543
rect 2973 11509 3007 11543
rect 3893 11509 3927 11543
rect 5641 11509 5675 11543
rect 5825 11509 5859 11543
rect 6009 11509 6043 11543
rect 7297 11509 7331 11543
rect 9321 11509 9355 11543
rect 11897 11509 11931 11543
rect 13369 11509 13403 11543
rect 14289 11509 14323 11543
rect 2053 11305 2087 11339
rect 5825 11305 5859 11339
rect 7297 11305 7331 11339
rect 8769 11305 8803 11339
rect 10517 11305 10551 11339
rect 15209 11305 15243 11339
rect 2881 11237 2915 11271
rect 4261 11237 4295 11271
rect 2513 11169 2547 11203
rect 2697 11169 2731 11203
rect 3341 11169 3375 11203
rect 3525 11169 3559 11203
rect 13461 11169 13495 11203
rect 14657 11169 14691 11203
rect 1685 11101 1719 11135
rect 2421 11101 2455 11135
rect 4077 11101 4111 11135
rect 4445 11101 4479 11135
rect 5917 11101 5951 11135
rect 6184 11101 6218 11135
rect 7389 11101 7423 11135
rect 9137 11101 9171 11135
rect 10609 11101 10643 11135
rect 3249 11033 3283 11067
rect 3801 11033 3835 11067
rect 4690 11033 4724 11067
rect 7656 11033 7690 11067
rect 9404 11033 9438 11067
rect 10865 11033 10899 11067
rect 13194 11033 13228 11067
rect 13921 11033 13955 11067
rect 14473 11033 14507 11067
rect 14565 11033 14599 11067
rect 14933 11033 14967 11067
rect 15301 11033 15335 11067
rect 1501 10965 1535 10999
rect 8953 10965 8987 10999
rect 11989 10965 12023 10999
rect 12081 10965 12115 10999
rect 14105 10965 14139 10999
rect 1869 10761 1903 10795
rect 2237 10761 2271 10795
rect 2329 10761 2363 10795
rect 2697 10761 2731 10795
rect 3157 10761 3191 10795
rect 3525 10761 3559 10795
rect 4353 10761 4387 10795
rect 4721 10761 4755 10795
rect 6469 10761 6503 10795
rect 10333 10761 10367 10795
rect 11989 10761 12023 10795
rect 12541 10761 12575 10795
rect 13277 10761 13311 10795
rect 3893 10693 3927 10727
rect 5834 10693 5868 10727
rect 12081 10693 12115 10727
rect 13185 10693 13219 10727
rect 1685 10625 1719 10659
rect 3065 10625 3099 10659
rect 7582 10625 7616 10659
rect 9220 10625 9254 10659
rect 2513 10557 2547 10591
rect 3341 10557 3375 10591
rect 3985 10557 4019 10591
rect 4169 10557 4203 10591
rect 6101 10557 6135 10591
rect 7849 10557 7883 10591
rect 8953 10557 8987 10591
rect 11897 10557 11931 10591
rect 13369 10557 13403 10591
rect 12449 10489 12483 10523
rect 12817 10489 12851 10523
rect 1501 10421 1535 10455
rect 4537 10421 4571 10455
rect 8033 10421 8067 10455
rect 8769 10421 8803 10455
rect 10517 10421 10551 10455
rect 1777 10217 1811 10251
rect 8769 10217 8803 10251
rect 2973 10149 3007 10183
rect 3893 10149 3927 10183
rect 2697 10081 2731 10115
rect 13185 10081 13219 10115
rect 15117 10081 15151 10115
rect 1685 10013 1719 10047
rect 1961 10013 1995 10047
rect 5006 10013 5040 10047
rect 5273 10013 5307 10047
rect 5457 10013 5491 10047
rect 5641 10013 5675 10047
rect 5825 10013 5859 10047
rect 7030 10013 7064 10047
rect 7297 10013 7331 10047
rect 7389 10013 7423 10047
rect 10149 10013 10183 10047
rect 15025 10013 15059 10047
rect 15393 10013 15427 10047
rect 7634 9945 7668 9979
rect 9965 9945 9999 9979
rect 10416 9945 10450 9979
rect 13001 9945 13035 9979
rect 14933 9945 14967 9979
rect 1501 9877 1535 9911
rect 2053 9877 2087 9911
rect 2421 9877 2455 9911
rect 2513 9877 2547 9911
rect 5917 9877 5951 9911
rect 11529 9877 11563 9911
rect 12633 9877 12667 9911
rect 13093 9877 13127 9911
rect 14565 9877 14599 9911
rect 15577 9877 15611 9911
rect 2329 9673 2363 9707
rect 9597 9673 9631 9707
rect 13185 9673 13219 9707
rect 14289 9673 14323 9707
rect 14749 9673 14783 9707
rect 5374 9605 5408 9639
rect 7604 9605 7638 9639
rect 8370 9605 8404 9639
rect 11345 9605 11379 9639
rect 15209 9605 15243 9639
rect 1685 9537 1719 9571
rect 1961 9537 1995 9571
rect 2697 9537 2731 9571
rect 4169 9537 4203 9571
rect 5641 9537 5675 9571
rect 10721 9537 10755 9571
rect 10977 9537 11011 9571
rect 12653 9537 12687 9571
rect 12909 9537 12943 9571
rect 13553 9537 13587 9571
rect 14657 9537 14691 9571
rect 2789 9469 2823 9503
rect 2973 9469 3007 9503
rect 3893 9469 3927 9503
rect 7849 9469 7883 9503
rect 8125 9469 8159 9503
rect 13645 9469 13679 9503
rect 13737 9469 13771 9503
rect 14841 9469 14875 9503
rect 15301 9469 15335 9503
rect 11529 9401 11563 9435
rect 1501 9333 1535 9367
rect 1777 9333 1811 9367
rect 4261 9333 4295 9367
rect 5825 9333 5859 9367
rect 6101 9333 6135 9367
rect 6469 9333 6503 9367
rect 8033 9333 8067 9367
rect 9505 9333 9539 9367
rect 2421 9129 2455 9163
rect 10057 9129 10091 9163
rect 14105 9129 14139 9163
rect 14933 9129 14967 9163
rect 12909 9061 12943 9095
rect 1869 8993 1903 9027
rect 3341 8993 3375 9027
rect 3525 8993 3559 9027
rect 13093 8993 13127 9027
rect 14749 8993 14783 9027
rect 15485 8993 15519 9027
rect 1961 8925 1995 8959
rect 3065 8925 3099 8959
rect 4445 8925 4479 8959
rect 5917 8925 5951 8959
rect 11437 8925 11471 8959
rect 11529 8925 11563 8959
rect 11785 8925 11819 8959
rect 15301 8925 15335 8959
rect 15393 8925 15427 8959
rect 2053 8857 2087 8891
rect 4690 8857 4724 8891
rect 6162 8857 6196 8891
rect 11192 8857 11226 8891
rect 13369 8857 13403 8891
rect 5825 8789 5859 8823
rect 7297 8789 7331 8823
rect 9413 8789 9447 8823
rect 9873 8789 9907 8823
rect 13277 8789 13311 8823
rect 13737 8789 13771 8823
rect 14473 8789 14507 8823
rect 14565 8789 14599 8823
rect 2421 8585 2455 8619
rect 2513 8585 2547 8619
rect 2881 8585 2915 8619
rect 2973 8585 3007 8619
rect 3341 8585 3375 8619
rect 3709 8585 3743 8619
rect 5549 8585 5583 8619
rect 5825 8585 5859 8619
rect 6009 8585 6043 8619
rect 6193 8585 6227 8619
rect 7205 8585 7239 8619
rect 7389 8585 7423 8619
rect 13369 8585 13403 8619
rect 13829 8585 13863 8619
rect 14381 8585 14415 8619
rect 14749 8585 14783 8619
rect 15393 8585 15427 8619
rect 1961 8517 1995 8551
rect 9198 8517 9232 8551
rect 14841 8517 14875 8551
rect 2053 8449 2087 8483
rect 4169 8449 4203 8483
rect 4425 8449 4459 8483
rect 8594 8449 8628 8483
rect 13461 8449 13495 8483
rect 1869 8381 1903 8415
rect 3157 8381 3191 8415
rect 3801 8381 3835 8415
rect 3985 8381 4019 8415
rect 8861 8381 8895 8415
rect 8953 8381 8987 8415
rect 13277 8381 13311 8415
rect 14933 8381 14967 8415
rect 7481 8313 7515 8347
rect 10333 8313 10367 8347
rect 12909 8313 12943 8347
rect 15485 8313 15519 8347
rect 10701 8245 10735 8279
rect 11529 8245 11563 8279
rect 12081 8245 12115 8279
rect 12725 8245 12759 8279
rect 1501 8041 1535 8075
rect 2881 8041 2915 8075
rect 3893 8041 3927 8075
rect 12265 8041 12299 8075
rect 14473 8041 14507 8075
rect 1777 7973 1811 8007
rect 12173 7973 12207 8007
rect 3525 7905 3559 7939
rect 15025 7905 15059 7939
rect 1685 7837 1719 7871
rect 1961 7837 1995 7871
rect 5017 7837 5051 7871
rect 5273 7837 5307 7871
rect 5457 7837 5491 7871
rect 6929 7837 6963 7871
rect 7205 7837 7239 7871
rect 8677 7837 8711 7871
rect 9045 7837 9079 7871
rect 9229 7837 9263 7871
rect 9321 7837 9355 7871
rect 10793 7837 10827 7871
rect 13645 7837 13679 7871
rect 2789 7769 2823 7803
rect 3341 7769 3375 7803
rect 6684 7769 6718 7803
rect 8410 7769 8444 7803
rect 9588 7769 9622 7803
rect 11060 7769 11094 7803
rect 13378 7769 13412 7803
rect 14933 7769 14967 7803
rect 3249 7701 3283 7735
rect 5549 7701 5583 7735
rect 7297 7701 7331 7735
rect 10701 7701 10735 7735
rect 14105 7701 14139 7735
rect 14289 7701 14323 7735
rect 14841 7701 14875 7735
rect 15485 7701 15519 7735
rect 15669 7701 15703 7735
rect 1777 7497 1811 7531
rect 2605 7497 2639 7531
rect 13001 7497 13035 7531
rect 15209 7497 15243 7531
rect 15577 7497 15611 7531
rect 3157 7429 3191 7463
rect 3801 7429 3835 7463
rect 9873 7429 9907 7463
rect 11774 7429 11808 7463
rect 14197 7429 14231 7463
rect 1685 7361 1719 7395
rect 1961 7361 1995 7395
rect 2145 7361 2179 7395
rect 5466 7361 5500 7395
rect 7001 7361 7035 7395
rect 9330 7361 9364 7395
rect 9597 7361 9631 7395
rect 9965 7361 9999 7395
rect 10232 7361 10266 7395
rect 13369 7361 13403 7395
rect 15117 7361 15151 7395
rect 3249 7293 3283 7327
rect 3433 7293 3467 7327
rect 5733 7293 5767 7327
rect 6745 7293 6779 7327
rect 11529 7293 11563 7327
rect 13461 7293 13495 7327
rect 13553 7293 13587 7327
rect 14289 7293 14323 7327
rect 14381 7293 14415 7327
rect 15301 7293 15335 7327
rect 2329 7225 2363 7259
rect 4077 7225 4111 7259
rect 8217 7225 8251 7259
rect 1501 7157 1535 7191
rect 2513 7157 2547 7191
rect 2789 7157 2823 7191
rect 3893 7157 3927 7191
rect 4353 7157 4387 7191
rect 5825 7157 5859 7191
rect 6101 7157 6135 7191
rect 6561 7157 6595 7191
rect 8125 7157 8159 7191
rect 11345 7157 11379 7191
rect 12909 7157 12943 7191
rect 13829 7157 13863 7191
rect 14749 7157 14783 7191
rect 1961 6953 1995 6987
rect 7297 6953 7331 6987
rect 9045 6953 9079 6987
rect 13921 6953 13955 6987
rect 1593 6817 1627 6851
rect 1777 6817 1811 6851
rect 3433 6817 3467 6851
rect 8769 6817 8803 6851
rect 13369 6817 13403 6851
rect 14657 6817 14691 6851
rect 15485 6817 15519 6851
rect 2605 6749 2639 6783
rect 4169 6749 4203 6783
rect 5825 6749 5859 6783
rect 5917 6749 5951 6783
rect 10425 6749 10459 6783
rect 11897 6749 11931 6783
rect 13737 6749 13771 6783
rect 14473 6749 14507 6783
rect 15393 6749 15427 6783
rect 2329 6681 2363 6715
rect 4414 6681 4448 6715
rect 6184 6681 6218 6715
rect 8524 6681 8558 6715
rect 11630 6681 11664 6715
rect 13102 6681 13136 6715
rect 15301 6681 15335 6715
rect 2145 6613 2179 6647
rect 2513 6613 2547 6647
rect 2789 6613 2823 6647
rect 3157 6613 3191 6647
rect 3249 6613 3283 6647
rect 3801 6613 3835 6647
rect 5549 6613 5583 6647
rect 7389 6613 7423 6647
rect 10517 6613 10551 6647
rect 11989 6613 12023 6647
rect 13553 6613 13587 6647
rect 14105 6613 14139 6647
rect 14565 6613 14599 6647
rect 14933 6613 14967 6647
rect 2053 6409 2087 6443
rect 2881 6409 2915 6443
rect 6193 6409 6227 6443
rect 11161 6409 11195 6443
rect 11621 6409 11655 6443
rect 11897 6409 11931 6443
rect 12357 6409 12391 6443
rect 13185 6409 13219 6443
rect 13737 6409 13771 6443
rect 14197 6409 14231 6443
rect 14565 6409 14599 6443
rect 14933 6409 14967 6443
rect 2973 6341 3007 6375
rect 4454 6341 4488 6375
rect 10793 6341 10827 6375
rect 11989 6341 12023 6375
rect 13277 6341 13311 6375
rect 1685 6273 1719 6307
rect 1961 6273 1995 6307
rect 2237 6273 2271 6307
rect 4721 6273 4755 6307
rect 4813 6273 4847 6307
rect 5069 6273 5103 6307
rect 7472 6273 7506 6307
rect 8944 6273 8978 6307
rect 12541 6273 12575 6307
rect 14105 6273 14139 6307
rect 15393 6273 15427 6307
rect 2421 6205 2455 6239
rect 3157 6205 3191 6239
rect 6469 6205 6503 6239
rect 6653 6205 6687 6239
rect 7113 6205 7147 6239
rect 7205 6205 7239 6239
rect 8677 6205 8711 6239
rect 13093 6205 13127 6239
rect 14381 6205 14415 6239
rect 15025 6205 15059 6239
rect 15117 6205 15151 6239
rect 1501 6137 1535 6171
rect 13645 6137 13679 6171
rect 1777 6069 1811 6103
rect 2513 6069 2547 6103
rect 3341 6069 3375 6103
rect 6745 6069 6779 6103
rect 8585 6069 8619 6103
rect 10057 6069 10091 6103
rect 11345 6069 11379 6103
rect 12173 6069 12207 6103
rect 12817 6069 12851 6103
rect 15577 6069 15611 6103
rect 2605 5865 2639 5899
rect 3433 5865 3467 5899
rect 5825 5865 5859 5899
rect 7389 5865 7423 5899
rect 8585 5865 8619 5899
rect 9597 5865 9631 5899
rect 11253 5865 11287 5899
rect 13829 5865 13863 5899
rect 14381 5865 14415 5899
rect 15393 5865 15427 5899
rect 3801 5797 3835 5831
rect 7573 5797 7607 5831
rect 7757 5797 7791 5831
rect 7849 5797 7883 5831
rect 8125 5797 8159 5831
rect 11161 5797 11195 5831
rect 2053 5729 2087 5763
rect 2145 5729 2179 5763
rect 2881 5729 2915 5763
rect 7205 5729 7239 5763
rect 9781 5729 9815 5763
rect 13369 5729 13403 5763
rect 15117 5729 15151 5763
rect 1685 5661 1719 5695
rect 3065 5661 3099 5695
rect 4261 5661 4295 5695
rect 4353 5661 4387 5695
rect 6949 5661 6983 5695
rect 12633 5661 12667 5695
rect 13185 5661 13219 5695
rect 13645 5661 13679 5695
rect 15577 5661 15611 5695
rect 4598 5593 4632 5627
rect 10026 5593 10060 5627
rect 12366 5593 12400 5627
rect 14657 5593 14691 5627
rect 1501 5525 1535 5559
rect 2237 5525 2271 5559
rect 2973 5525 3007 5559
rect 3617 5525 3651 5559
rect 3985 5525 4019 5559
rect 5733 5525 5767 5559
rect 8217 5525 8251 5559
rect 8769 5525 8803 5559
rect 12817 5525 12851 5559
rect 13277 5525 13311 5559
rect 14105 5525 14139 5559
rect 14749 5525 14783 5559
rect 15025 5525 15059 5559
rect 2237 5321 2271 5355
rect 2329 5321 2363 5355
rect 3433 5321 3467 5355
rect 3525 5321 3559 5355
rect 3985 5321 4019 5355
rect 4629 5321 4663 5355
rect 5089 5321 5123 5355
rect 5457 5321 5491 5355
rect 6469 5321 6503 5355
rect 7021 5321 7055 5355
rect 8309 5321 8343 5355
rect 9873 5321 9907 5355
rect 11161 5321 11195 5355
rect 13369 5321 13403 5355
rect 14197 5321 14231 5355
rect 15209 5321 15243 5355
rect 3065 5253 3099 5287
rect 11621 5253 11655 5287
rect 13277 5253 13311 5287
rect 1869 5185 1903 5219
rect 2513 5185 2547 5219
rect 3893 5185 3927 5219
rect 4997 5185 5031 5219
rect 5825 5185 5859 5219
rect 6929 5185 6963 5219
rect 7757 5185 7791 5219
rect 8401 5185 8435 5219
rect 8657 5185 8691 5219
rect 10241 5185 10275 5219
rect 12449 5185 12483 5219
rect 14105 5185 14139 5219
rect 14841 5185 14875 5219
rect 15485 5185 15519 5219
rect 1593 5117 1627 5151
rect 1777 5117 1811 5151
rect 2881 5117 2915 5151
rect 2973 5117 3007 5151
rect 4077 5117 4111 5151
rect 4537 5117 4571 5151
rect 5273 5117 5307 5151
rect 5917 5117 5951 5151
rect 6101 5117 6135 5151
rect 7205 5117 7239 5151
rect 7849 5117 7883 5151
rect 7941 5117 7975 5151
rect 10333 5117 10367 5151
rect 10425 5117 10459 5151
rect 11345 5117 11379 5151
rect 11989 5117 12023 5151
rect 12541 5117 12575 5151
rect 12633 5117 12667 5151
rect 13461 5117 13495 5151
rect 14289 5117 14323 5151
rect 14565 5117 14599 5151
rect 7389 5049 7423 5083
rect 6561 4981 6595 5015
rect 9781 4981 9815 5015
rect 10701 4981 10735 5015
rect 10885 4981 10919 5015
rect 12081 4981 12115 5015
rect 12909 4981 12943 5015
rect 13737 4981 13771 5015
rect 15117 4981 15151 5015
rect 15669 4981 15703 5015
rect 1869 4777 1903 4811
rect 3985 4777 4019 4811
rect 5641 4777 5675 4811
rect 6193 4777 6227 4811
rect 8953 4777 8987 4811
rect 9505 4777 9539 4811
rect 10333 4777 10367 4811
rect 10793 4777 10827 4811
rect 10977 4777 11011 4811
rect 11529 4777 11563 4811
rect 14933 4777 14967 4811
rect 2881 4709 2915 4743
rect 4353 4709 4387 4743
rect 8585 4709 8619 4743
rect 11253 4709 11287 4743
rect 2513 4641 2547 4675
rect 3433 4641 3467 4675
rect 4997 4641 5031 4675
rect 6653 4641 6687 4675
rect 6837 4641 6871 4675
rect 7113 4641 7147 4675
rect 7297 4641 7331 4675
rect 8033 4641 8067 4675
rect 9689 4641 9723 4675
rect 12081 4641 12115 4675
rect 12909 4641 12943 4675
rect 13645 4641 13679 4675
rect 13737 4641 13771 4675
rect 14657 4641 14691 4675
rect 1685 4573 1719 4607
rect 3801 4573 3835 4607
rect 4169 4573 4203 4607
rect 6101 4573 6135 4607
rect 9137 4573 9171 4607
rect 10425 4573 10459 4607
rect 10701 4573 10735 4607
rect 11437 4573 11471 4607
rect 12725 4573 12759 4607
rect 14473 4573 14507 4607
rect 15117 4573 15151 4607
rect 15485 4573 15519 4607
rect 2237 4505 2271 4539
rect 7389 4505 7423 4539
rect 8677 4505 8711 4539
rect 9229 4505 9263 4539
rect 11897 4505 11931 4539
rect 13553 4505 13587 4539
rect 1501 4437 1535 4471
rect 2329 4437 2363 4471
rect 2789 4437 2823 4471
rect 3249 4437 3283 4471
rect 3341 4437 3375 4471
rect 4445 4437 4479 4471
rect 4813 4437 4847 4471
rect 4905 4437 4939 4471
rect 5457 4437 5491 4471
rect 5917 4437 5951 4471
rect 6561 4437 6595 4471
rect 7757 4437 7791 4471
rect 8125 4437 8159 4471
rect 8217 4437 8251 4471
rect 9873 4437 9907 4471
rect 9965 4437 9999 4471
rect 11989 4437 12023 4471
rect 12357 4437 12391 4471
rect 12817 4437 12851 4471
rect 13185 4437 13219 4471
rect 14105 4437 14139 4471
rect 14565 4437 14599 4471
rect 15393 4437 15427 4471
rect 1685 4233 1719 4267
rect 2053 4233 2087 4267
rect 2973 4233 3007 4267
rect 3341 4233 3375 4267
rect 3801 4233 3835 4267
rect 5181 4233 5215 4267
rect 5549 4233 5583 4267
rect 6009 4233 6043 4267
rect 7941 4233 7975 4267
rect 8033 4233 8067 4267
rect 8401 4233 8435 4267
rect 9413 4233 9447 4267
rect 10333 4233 10367 4267
rect 10701 4233 10735 4267
rect 11161 4233 11195 4267
rect 11529 4233 11563 4267
rect 11897 4233 11931 4267
rect 13093 4233 13127 4267
rect 13921 4233 13955 4267
rect 12541 4165 12575 4199
rect 1593 4097 1627 4131
rect 2145 4097 2179 4131
rect 2881 4097 2915 4131
rect 4537 4097 4571 4131
rect 5641 4097 5675 4131
rect 6193 4097 6227 4131
rect 6469 4097 6503 4131
rect 7021 4097 7055 4131
rect 7573 4097 7607 4131
rect 8769 4097 8803 4131
rect 8861 4097 8895 4131
rect 9505 4097 9539 4131
rect 9965 4097 9999 4131
rect 11345 4097 11379 4131
rect 11989 4097 12023 4131
rect 14473 4097 14507 4131
rect 15669 4097 15703 4131
rect 2329 4029 2363 4063
rect 2697 4029 2731 4063
rect 3893 4029 3927 4063
rect 4077 4029 4111 4063
rect 4261 4029 4295 4063
rect 5733 4029 5767 4063
rect 7297 4029 7331 4063
rect 7849 4029 7883 4063
rect 9321 4029 9355 4063
rect 10793 4029 10827 4063
rect 10977 4029 11011 4063
rect 12081 4029 12115 4063
rect 12357 4029 12391 4063
rect 13185 4029 13219 4063
rect 13369 4029 13403 4063
rect 14013 4029 14047 4063
rect 14197 4029 14231 4063
rect 15393 4029 15427 4063
rect 6653 3961 6687 3995
rect 9873 3961 9907 3995
rect 10149 3961 10183 3995
rect 1409 3893 1443 3927
rect 3433 3893 3467 3927
rect 6837 3893 6871 3927
rect 7389 3893 7423 3927
rect 8585 3893 8619 3927
rect 9045 3893 9079 3927
rect 12725 3893 12759 3927
rect 13553 3893 13587 3927
rect 14657 3893 14691 3927
rect 2697 3689 2731 3723
rect 3617 3689 3651 3723
rect 6009 3689 6043 3723
rect 7849 3689 7883 3723
rect 9781 3689 9815 3723
rect 10517 3689 10551 3723
rect 11345 3689 11379 3723
rect 12173 3689 12207 3723
rect 1869 3621 1903 3655
rect 5089 3621 5123 3655
rect 14105 3621 14139 3655
rect 14749 3621 14783 3655
rect 3249 3553 3283 3587
rect 4997 3553 5031 3587
rect 5641 3553 5675 3587
rect 6653 3553 6687 3587
rect 7481 3553 7515 3587
rect 8401 3553 8435 3587
rect 9137 3553 9171 3587
rect 11161 3553 11195 3587
rect 11805 3553 11839 3587
rect 11989 3553 12023 3587
rect 12725 3553 12759 3587
rect 13093 3553 13127 3587
rect 13369 3553 13403 3587
rect 14841 3553 14875 3587
rect 1409 3485 1443 3519
rect 2145 3485 2179 3519
rect 2421 3485 2455 3519
rect 3065 3485 3099 3519
rect 4077 3485 4111 3519
rect 4721 3485 4755 3519
rect 5549 3485 5583 3519
rect 7205 3485 7239 3519
rect 7757 3485 7791 3519
rect 8217 3485 8251 3519
rect 10885 3485 10919 3519
rect 12541 3485 12575 3519
rect 14289 3485 14323 3519
rect 15117 3485 15151 3519
rect 2605 3417 2639 3451
rect 6469 3417 6503 3451
rect 8769 3417 8803 3451
rect 10333 3417 10367 3451
rect 11713 3417 11747 3451
rect 14565 3417 14599 3451
rect 1593 3349 1627 3383
rect 1961 3349 1995 3383
rect 2237 3349 2271 3383
rect 3157 3349 3191 3383
rect 3893 3349 3927 3383
rect 5457 3349 5491 3383
rect 6377 3349 6411 3383
rect 6837 3349 6871 3383
rect 7297 3349 7331 3383
rect 8309 3349 8343 3383
rect 9321 3349 9355 3383
rect 9413 3349 9447 3383
rect 10057 3349 10091 3383
rect 10241 3349 10275 3383
rect 10977 3349 11011 3383
rect 12633 3349 12667 3383
rect 3709 3145 3743 3179
rect 4169 3145 4203 3179
rect 5089 3145 5123 3179
rect 5641 3145 5675 3179
rect 6377 3145 6411 3179
rect 6745 3145 6779 3179
rect 8033 3145 8067 3179
rect 8953 3145 8987 3179
rect 9413 3145 9447 3179
rect 9781 3145 9815 3179
rect 10609 3145 10643 3179
rect 10701 3145 10735 3179
rect 11161 3145 11195 3179
rect 12265 3145 12299 3179
rect 12357 3145 12391 3179
rect 12817 3145 12851 3179
rect 4077 3077 4111 3111
rect 11253 3077 11287 3111
rect 11805 3077 11839 3111
rect 12725 3077 12759 3111
rect 1685 3009 1719 3043
rect 1961 3009 1995 3043
rect 2237 3009 2271 3043
rect 2329 3009 2363 3043
rect 2789 3009 2823 3043
rect 2881 3009 2915 3043
rect 3433 3009 3467 3043
rect 4813 3009 4847 3043
rect 4905 3009 4939 3043
rect 5365 3009 5399 3043
rect 5457 3009 5491 3043
rect 5733 3009 5767 3043
rect 7205 3009 7239 3043
rect 7665 3009 7699 3043
rect 8125 3009 8159 3043
rect 9045 3009 9079 3043
rect 9873 3009 9907 3043
rect 11897 3009 11931 3043
rect 14105 3009 14139 3043
rect 14289 3009 14323 3043
rect 14565 3009 14599 3043
rect 15669 3009 15703 3043
rect 4353 2941 4387 2975
rect 6837 2941 6871 2975
rect 7021 2941 7055 2975
rect 7849 2941 7883 2975
rect 9137 2941 9171 2975
rect 9965 2941 9999 2975
rect 10793 2941 10827 2975
rect 11713 2941 11747 2975
rect 13001 2941 13035 2975
rect 13185 2941 13219 2975
rect 13461 2941 13495 2975
rect 14841 2941 14875 2975
rect 1777 2873 1811 2907
rect 2513 2873 2547 2907
rect 3065 2873 3099 2907
rect 3617 2873 3651 2907
rect 8585 2873 8619 2907
rect 10241 2873 10275 2907
rect 1501 2805 1535 2839
rect 2053 2805 2087 2839
rect 2605 2805 2639 2839
rect 3249 2805 3283 2839
rect 4629 2805 4663 2839
rect 5181 2805 5215 2839
rect 5917 2805 5951 2839
rect 6193 2805 6227 2839
rect 7389 2805 7423 2839
rect 8493 2805 8527 2839
rect 15485 2805 15519 2839
rect 7757 2601 7791 2635
rect 9045 2601 9079 2635
rect 9413 2601 9447 2635
rect 10425 2601 10459 2635
rect 12219 2601 12253 2635
rect 3985 2533 4019 2567
rect 7481 2533 7515 2567
rect 8033 2533 8067 2567
rect 11529 2533 11563 2567
rect 8493 2465 8527 2499
rect 8677 2465 8711 2499
rect 9873 2465 9907 2499
rect 9965 2465 9999 2499
rect 15393 2465 15427 2499
rect 1777 2397 1811 2431
rect 1869 2397 1903 2431
rect 2237 2397 2271 2431
rect 2605 2397 2639 2431
rect 2973 2397 3007 2431
rect 3341 2397 3375 2431
rect 3801 2397 3835 2431
rect 4077 2397 4111 2431
rect 4721 2397 4755 2431
rect 5089 2397 5123 2431
rect 5181 2397 5215 2431
rect 5825 2397 5859 2431
rect 6193 2397 6227 2431
rect 6561 2397 6595 2431
rect 7205 2397 7239 2431
rect 7297 2397 7331 2431
rect 7941 2397 7975 2431
rect 8401 2397 8435 2431
rect 10517 2397 10551 2431
rect 10793 2397 10827 2431
rect 11713 2397 11747 2431
rect 11989 2397 12023 2431
rect 12909 2397 12943 2431
rect 13185 2397 13219 2431
rect 14105 2397 14139 2431
rect 14381 2397 14415 2431
rect 15117 2397 15151 2431
rect 9137 2329 9171 2363
rect 9505 2329 9539 2363
rect 1593 2261 1627 2295
rect 2053 2261 2087 2295
rect 2421 2261 2455 2295
rect 2789 2261 2823 2295
rect 3157 2261 3191 2295
rect 3525 2261 3559 2295
rect 4261 2261 4295 2295
rect 4537 2261 4571 2295
rect 4905 2261 4939 2295
rect 5365 2261 5399 2295
rect 5641 2261 5675 2295
rect 6009 2261 6043 2295
rect 6469 2261 6503 2295
rect 6745 2261 6779 2295
rect 7021 2261 7055 2295
rect 10057 2261 10091 2295
rect 13829 2261 13863 2295
<< metal1 >>
rect 4062 17756 4068 17808
rect 4120 17796 4126 17808
rect 15286 17796 15292 17808
rect 4120 17768 15292 17796
rect 4120 17756 4126 17768
rect 15286 17756 15292 17768
rect 15344 17756 15350 17808
rect 5350 17688 5356 17740
rect 5408 17728 5414 17740
rect 13538 17728 13544 17740
rect 5408 17700 13544 17728
rect 5408 17688 5414 17700
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 7466 17620 7472 17672
rect 7524 17660 7530 17672
rect 10134 17660 10140 17672
rect 7524 17632 10140 17660
rect 7524 17620 7530 17632
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 7006 17552 7012 17604
rect 7064 17592 7070 17604
rect 8202 17592 8208 17604
rect 7064 17564 8208 17592
rect 7064 17552 7070 17564
rect 8202 17552 8208 17564
rect 8260 17592 8266 17604
rect 13446 17592 13452 17604
rect 8260 17564 13452 17592
rect 8260 17552 8266 17564
rect 13446 17552 13452 17564
rect 13504 17552 13510 17604
rect 7374 17484 7380 17536
rect 7432 17524 7438 17536
rect 8018 17524 8024 17536
rect 7432 17496 8024 17524
rect 7432 17484 7438 17496
rect 8018 17484 8024 17496
rect 8076 17484 8082 17536
rect 1104 17434 16008 17456
rect 1104 17382 4698 17434
rect 4750 17382 4762 17434
rect 4814 17382 4826 17434
rect 4878 17382 4890 17434
rect 4942 17382 4954 17434
rect 5006 17382 8446 17434
rect 8498 17382 8510 17434
rect 8562 17382 8574 17434
rect 8626 17382 8638 17434
rect 8690 17382 8702 17434
rect 8754 17382 12194 17434
rect 12246 17382 12258 17434
rect 12310 17382 12322 17434
rect 12374 17382 12386 17434
rect 12438 17382 12450 17434
rect 12502 17382 16008 17434
rect 1104 17360 16008 17382
rect 1581 17323 1639 17329
rect 1581 17289 1593 17323
rect 1627 17320 1639 17323
rect 1762 17320 1768 17332
rect 1627 17292 1768 17320
rect 1627 17289 1639 17292
rect 1581 17283 1639 17289
rect 1762 17280 1768 17292
rect 1820 17280 1826 17332
rect 1949 17323 2007 17329
rect 1949 17289 1961 17323
rect 1995 17320 2007 17323
rect 2130 17320 2136 17332
rect 1995 17292 2136 17320
rect 1995 17289 2007 17292
rect 1949 17283 2007 17289
rect 2130 17280 2136 17292
rect 2188 17280 2194 17332
rect 2317 17323 2375 17329
rect 2317 17289 2329 17323
rect 2363 17320 2375 17323
rect 2498 17320 2504 17332
rect 2363 17292 2504 17320
rect 2363 17289 2375 17292
rect 2317 17283 2375 17289
rect 2498 17280 2504 17292
rect 2556 17280 2562 17332
rect 2685 17323 2743 17329
rect 2685 17289 2697 17323
rect 2731 17320 2743 17323
rect 2866 17320 2872 17332
rect 2731 17292 2872 17320
rect 2731 17289 2743 17292
rect 2685 17283 2743 17289
rect 2866 17280 2872 17292
rect 2924 17280 2930 17332
rect 3053 17323 3111 17329
rect 3053 17289 3065 17323
rect 3099 17320 3111 17323
rect 3234 17320 3240 17332
rect 3099 17292 3240 17320
rect 3099 17289 3111 17292
rect 3053 17283 3111 17289
rect 3234 17280 3240 17292
rect 3292 17280 3298 17332
rect 3513 17323 3571 17329
rect 3513 17289 3525 17323
rect 3559 17320 3571 17323
rect 3602 17320 3608 17332
rect 3559 17292 3608 17320
rect 3559 17289 3571 17292
rect 3513 17283 3571 17289
rect 3602 17280 3608 17292
rect 3660 17280 3666 17332
rect 3973 17323 4031 17329
rect 3973 17289 3985 17323
rect 4019 17320 4031 17323
rect 4062 17320 4068 17332
rect 4019 17292 4068 17320
rect 4019 17289 4031 17292
rect 3973 17283 4031 17289
rect 4062 17280 4068 17292
rect 4120 17280 4126 17332
rect 4249 17323 4307 17329
rect 4249 17289 4261 17323
rect 4295 17320 4307 17323
rect 4338 17320 4344 17332
rect 4295 17292 4344 17320
rect 4295 17289 4307 17292
rect 4249 17283 4307 17289
rect 4338 17280 4344 17292
rect 4396 17280 4402 17332
rect 4525 17323 4583 17329
rect 4525 17289 4537 17323
rect 4571 17320 4583 17323
rect 4614 17320 4620 17332
rect 4571 17292 4620 17320
rect 4571 17289 4583 17292
rect 4525 17283 4583 17289
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 4893 17323 4951 17329
rect 4893 17289 4905 17323
rect 4939 17320 4951 17323
rect 5442 17320 5448 17332
rect 4939 17292 5448 17320
rect 4939 17289 4951 17292
rect 4893 17283 4951 17289
rect 5442 17280 5448 17292
rect 5500 17280 5506 17332
rect 5629 17323 5687 17329
rect 5629 17289 5641 17323
rect 5675 17289 5687 17323
rect 5629 17283 5687 17289
rect 6089 17323 6147 17329
rect 6089 17289 6101 17323
rect 6135 17320 6147 17323
rect 6914 17320 6920 17332
rect 6135 17292 6920 17320
rect 6135 17289 6147 17292
rect 6089 17283 6147 17289
rect 4430 17252 4436 17264
rect 2884 17224 4436 17252
rect 1762 17184 1768 17196
rect 1723 17156 1768 17184
rect 1762 17144 1768 17156
rect 1820 17144 1826 17196
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17184 2191 17187
rect 2406 17184 2412 17196
rect 2179 17156 2412 17184
rect 2179 17153 2191 17156
rect 2133 17147 2191 17153
rect 2406 17144 2412 17156
rect 2464 17144 2470 17196
rect 2884 17193 2912 17224
rect 4430 17212 4436 17224
rect 4488 17212 4494 17264
rect 5644 17252 5672 17283
rect 6914 17280 6920 17292
rect 6972 17280 6978 17332
rect 7285 17323 7343 17329
rect 7285 17289 7297 17323
rect 7331 17320 7343 17323
rect 7374 17320 7380 17332
rect 7331 17292 7380 17320
rect 7331 17289 7343 17292
rect 7285 17283 7343 17289
rect 7374 17280 7380 17292
rect 7432 17280 7438 17332
rect 7558 17320 7564 17332
rect 7519 17292 7564 17320
rect 7558 17280 7564 17292
rect 7616 17280 7622 17332
rect 8018 17320 8024 17332
rect 7979 17292 8024 17320
rect 8018 17280 8024 17292
rect 8076 17280 8082 17332
rect 8294 17280 8300 17332
rect 8352 17320 8358 17332
rect 8573 17323 8631 17329
rect 8573 17320 8585 17323
rect 8352 17292 8585 17320
rect 8352 17280 8358 17292
rect 8573 17289 8585 17292
rect 8619 17289 8631 17323
rect 13446 17320 13452 17332
rect 13407 17292 13452 17320
rect 8573 17283 8631 17289
rect 13446 17280 13452 17292
rect 13504 17280 13510 17332
rect 13725 17323 13783 17329
rect 13725 17289 13737 17323
rect 13771 17289 13783 17323
rect 13725 17283 13783 17289
rect 6546 17252 6552 17264
rect 5644 17224 6552 17252
rect 6546 17212 6552 17224
rect 6604 17212 6610 17264
rect 13740 17252 13768 17283
rect 7116 17224 13768 17252
rect 13832 17224 14136 17252
rect 2501 17187 2559 17193
rect 2501 17153 2513 17187
rect 2547 17153 2559 17187
rect 2501 17147 2559 17153
rect 2869 17187 2927 17193
rect 2869 17153 2881 17187
rect 2915 17153 2927 17187
rect 3234 17184 3240 17196
rect 3195 17156 3240 17184
rect 2869 17147 2927 17153
rect 2516 17116 2544 17147
rect 3234 17144 3240 17156
rect 3292 17144 3298 17196
rect 3326 17144 3332 17196
rect 3384 17184 3390 17196
rect 3789 17187 3847 17193
rect 3384 17156 3429 17184
rect 3384 17144 3390 17156
rect 3789 17153 3801 17187
rect 3835 17153 3847 17187
rect 3789 17147 3847 17153
rect 4065 17187 4123 17193
rect 4065 17153 4077 17187
rect 4111 17184 4123 17187
rect 4246 17184 4252 17196
rect 4111 17156 4252 17184
rect 4111 17153 4123 17156
rect 4065 17147 4123 17153
rect 3142 17116 3148 17128
rect 2516 17088 3148 17116
rect 3142 17076 3148 17088
rect 3200 17076 3206 17128
rect 1026 17008 1032 17060
rect 1084 17048 1090 17060
rect 3804 17048 3832 17147
rect 4246 17144 4252 17156
rect 4304 17144 4310 17196
rect 4706 17184 4712 17196
rect 4667 17156 4712 17184
rect 4706 17144 4712 17156
rect 4764 17144 4770 17196
rect 5077 17187 5135 17193
rect 5077 17153 5089 17187
rect 5123 17184 5135 17187
rect 5350 17184 5356 17196
rect 5123 17156 5356 17184
rect 5123 17153 5135 17156
rect 5077 17147 5135 17153
rect 5350 17144 5356 17156
rect 5408 17144 5414 17196
rect 5442 17144 5448 17196
rect 5500 17184 5506 17196
rect 5810 17184 5816 17196
rect 5500 17156 5545 17184
rect 5771 17156 5816 17184
rect 5500 17144 5506 17156
rect 5810 17144 5816 17156
rect 5868 17144 5874 17196
rect 5905 17187 5963 17193
rect 5905 17153 5917 17187
rect 5951 17153 5963 17187
rect 5905 17147 5963 17153
rect 5166 17076 5172 17128
rect 5224 17116 5230 17128
rect 5920 17116 5948 17147
rect 6454 17144 6460 17196
rect 6512 17184 6518 17196
rect 7116 17193 7144 17224
rect 6733 17187 6791 17193
rect 6733 17184 6745 17187
rect 6512 17156 6745 17184
rect 6512 17144 6518 17156
rect 6733 17153 6745 17156
rect 6779 17153 6791 17187
rect 6733 17147 6791 17153
rect 7101 17187 7159 17193
rect 7101 17153 7113 17187
rect 7147 17153 7159 17187
rect 7101 17147 7159 17153
rect 7462 17187 7520 17193
rect 7462 17153 7474 17187
rect 7508 17153 7520 17187
rect 7926 17184 7932 17196
rect 7887 17156 7932 17184
rect 7462 17147 7520 17153
rect 7282 17116 7288 17128
rect 5224 17088 5948 17116
rect 6564 17088 7288 17116
rect 5224 17076 5230 17088
rect 1084 17020 3832 17048
rect 5261 17051 5319 17057
rect 1084 17008 1090 17020
rect 5261 17017 5273 17051
rect 5307 17048 5319 17051
rect 6178 17048 6184 17060
rect 5307 17020 6184 17048
rect 5307 17017 5319 17020
rect 5261 17011 5319 17017
rect 6178 17008 6184 17020
rect 6236 17008 6242 17060
rect 6564 17057 6592 17088
rect 7282 17076 7288 17088
rect 7340 17076 7346 17128
rect 7484 17116 7512 17147
rect 7926 17144 7932 17156
rect 7984 17144 7990 17196
rect 8757 17187 8815 17193
rect 8757 17153 8769 17187
rect 8803 17153 8815 17187
rect 8757 17147 8815 17153
rect 9309 17187 9367 17193
rect 9309 17153 9321 17187
rect 9355 17184 9367 17187
rect 9674 17184 9680 17196
rect 9355 17156 9680 17184
rect 9355 17153 9367 17156
rect 9309 17147 9367 17153
rect 8202 17116 8208 17128
rect 7484 17088 8064 17116
rect 8163 17088 8208 17116
rect 6549 17051 6607 17057
rect 6549 17017 6561 17051
rect 6595 17017 6607 17051
rect 6549 17011 6607 17017
rect 6917 17051 6975 17057
rect 6917 17017 6929 17051
rect 6963 17048 6975 17051
rect 7650 17048 7656 17060
rect 6963 17020 7656 17048
rect 6963 17017 6975 17020
rect 6917 17011 6975 17017
rect 7650 17008 7656 17020
rect 7708 17008 7714 17060
rect 8036 17048 8064 17088
rect 8202 17076 8208 17088
rect 8260 17076 8266 17128
rect 8294 17048 8300 17060
rect 8036 17020 8300 17048
rect 8294 17008 8300 17020
rect 8352 17008 8358 17060
rect 8772 17048 8800 17147
rect 9674 17144 9680 17156
rect 9732 17144 9738 17196
rect 9861 17187 9919 17193
rect 9861 17153 9873 17187
rect 9907 17184 9919 17187
rect 9950 17184 9956 17196
rect 9907 17156 9956 17184
rect 9907 17153 9919 17156
rect 9861 17147 9919 17153
rect 9950 17144 9956 17156
rect 10008 17144 10014 17196
rect 10134 17144 10140 17196
rect 10192 17184 10198 17196
rect 10597 17187 10655 17193
rect 10597 17184 10609 17187
rect 10192 17156 10609 17184
rect 10192 17144 10198 17156
rect 10597 17153 10609 17156
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 10686 17144 10692 17196
rect 10744 17184 10750 17196
rect 10870 17184 10876 17196
rect 10744 17156 10876 17184
rect 10744 17144 10750 17156
rect 10870 17144 10876 17156
rect 10928 17184 10934 17196
rect 11517 17187 11575 17193
rect 11517 17184 11529 17187
rect 10928 17156 11529 17184
rect 10928 17144 10934 17156
rect 11517 17153 11529 17156
rect 11563 17153 11575 17187
rect 11517 17147 11575 17153
rect 11698 17144 11704 17196
rect 11756 17184 11762 17196
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 11756 17156 12449 17184
rect 11756 17144 11762 17156
rect 12437 17153 12449 17156
rect 12483 17153 12495 17187
rect 12437 17147 12495 17153
rect 12526 17144 12532 17196
rect 12584 17184 12590 17196
rect 13078 17184 13084 17196
rect 12584 17156 13084 17184
rect 12584 17144 12590 17156
rect 13078 17144 13084 17156
rect 13136 17184 13142 17196
rect 13541 17187 13599 17193
rect 13541 17184 13553 17187
rect 13136 17156 13553 17184
rect 13136 17144 13142 17156
rect 13541 17153 13553 17156
rect 13587 17153 13599 17187
rect 13541 17147 13599 17153
rect 9398 17076 9404 17128
rect 9456 17116 9462 17128
rect 9585 17119 9643 17125
rect 9585 17116 9597 17119
rect 9456 17088 9597 17116
rect 9456 17076 9462 17088
rect 9585 17085 9597 17088
rect 9631 17085 9643 17119
rect 9585 17079 9643 17085
rect 9769 17119 9827 17125
rect 9769 17085 9781 17119
rect 9815 17116 9827 17119
rect 10042 17116 10048 17128
rect 9815 17088 10048 17116
rect 9815 17085 9827 17088
rect 9769 17079 9827 17085
rect 10042 17076 10048 17088
rect 10100 17076 10106 17128
rect 10226 17076 10232 17128
rect 10284 17116 10290 17128
rect 10321 17119 10379 17125
rect 10321 17116 10333 17119
rect 10284 17088 10333 17116
rect 10284 17076 10290 17088
rect 10321 17085 10333 17088
rect 10367 17085 10379 17119
rect 11790 17116 11796 17128
rect 11751 17088 11796 17116
rect 10321 17079 10379 17085
rect 11790 17076 11796 17088
rect 11848 17076 11854 17128
rect 12710 17116 12716 17128
rect 12671 17088 12716 17116
rect 12710 17076 12716 17088
rect 12768 17076 12774 17128
rect 13170 17076 13176 17128
rect 13228 17116 13234 17128
rect 13832 17116 13860 17224
rect 14108 17193 14136 17224
rect 13909 17187 13967 17193
rect 13909 17153 13921 17187
rect 13955 17153 13967 17187
rect 13909 17147 13967 17153
rect 14093 17187 14151 17193
rect 14093 17153 14105 17187
rect 14139 17184 14151 17187
rect 14458 17184 14464 17196
rect 14139 17156 14464 17184
rect 14139 17153 14151 17156
rect 14093 17147 14151 17153
rect 13228 17088 13860 17116
rect 13228 17076 13234 17088
rect 11054 17048 11060 17060
rect 8772 17020 11060 17048
rect 11054 17008 11060 17020
rect 11112 17008 11118 17060
rect 13924 17048 13952 17147
rect 14458 17144 14464 17156
rect 14516 17144 14522 17196
rect 15105 17187 15163 17193
rect 15105 17153 15117 17187
rect 15151 17184 15163 17187
rect 15378 17184 15384 17196
rect 15151 17156 15384 17184
rect 15151 17153 15163 17156
rect 15105 17147 15163 17153
rect 15378 17144 15384 17156
rect 15436 17144 15442 17196
rect 14366 17116 14372 17128
rect 14327 17088 14372 17116
rect 14366 17076 14372 17088
rect 14424 17076 14430 17128
rect 15194 17076 15200 17128
rect 15252 17116 15258 17128
rect 15289 17119 15347 17125
rect 15289 17116 15301 17119
rect 15252 17088 15301 17116
rect 15252 17076 15258 17088
rect 15289 17085 15301 17088
rect 15335 17085 15347 17119
rect 15289 17079 15347 17085
rect 15102 17048 15108 17060
rect 13924 17020 15108 17048
rect 15102 17008 15108 17020
rect 15160 17008 15166 17060
rect 5442 16940 5448 16992
rect 5500 16980 5506 16992
rect 8018 16980 8024 16992
rect 5500 16952 8024 16980
rect 5500 16940 5506 16952
rect 8018 16940 8024 16952
rect 8076 16940 8082 16992
rect 9030 16980 9036 16992
rect 8991 16952 9036 16980
rect 9030 16940 9036 16952
rect 9088 16940 9094 16992
rect 9217 16983 9275 16989
rect 9217 16949 9229 16983
rect 9263 16980 9275 16983
rect 9582 16980 9588 16992
rect 9263 16952 9588 16980
rect 9263 16949 9275 16952
rect 9217 16943 9275 16949
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 10229 16983 10287 16989
rect 10229 16980 10241 16983
rect 10192 16952 10241 16980
rect 10192 16940 10198 16952
rect 10229 16949 10241 16952
rect 10275 16949 10287 16983
rect 10229 16943 10287 16949
rect 10686 16940 10692 16992
rect 10744 16980 10750 16992
rect 11241 16983 11299 16989
rect 11241 16980 11253 16983
rect 10744 16952 11253 16980
rect 10744 16940 10750 16952
rect 11241 16949 11253 16952
rect 11287 16949 11299 16983
rect 11241 16943 11299 16949
rect 13814 16940 13820 16992
rect 13872 16980 13878 16992
rect 15838 16980 15844 16992
rect 13872 16952 15844 16980
rect 13872 16940 13878 16952
rect 15838 16940 15844 16952
rect 15896 16980 15902 16992
rect 16022 16980 16028 16992
rect 15896 16952 16028 16980
rect 15896 16940 15902 16952
rect 16022 16940 16028 16952
rect 16080 16940 16086 16992
rect 1104 16890 16008 16912
rect 1104 16838 2824 16890
rect 2876 16838 2888 16890
rect 2940 16838 2952 16890
rect 3004 16838 3016 16890
rect 3068 16838 3080 16890
rect 3132 16838 6572 16890
rect 6624 16838 6636 16890
rect 6688 16838 6700 16890
rect 6752 16838 6764 16890
rect 6816 16838 6828 16890
rect 6880 16838 10320 16890
rect 10372 16838 10384 16890
rect 10436 16838 10448 16890
rect 10500 16838 10512 16890
rect 10564 16838 10576 16890
rect 10628 16838 14068 16890
rect 14120 16838 14132 16890
rect 14184 16838 14196 16890
rect 14248 16838 14260 16890
rect 14312 16838 14324 16890
rect 14376 16838 16008 16890
rect 1104 16816 16008 16838
rect 1762 16736 1768 16788
rect 1820 16776 1826 16788
rect 2593 16779 2651 16785
rect 2593 16776 2605 16779
rect 1820 16748 2605 16776
rect 1820 16736 1826 16748
rect 2593 16745 2605 16748
rect 2639 16745 2651 16779
rect 2593 16739 2651 16745
rect 2869 16779 2927 16785
rect 2869 16745 2881 16779
rect 2915 16776 2927 16779
rect 3142 16776 3148 16788
rect 2915 16748 3148 16776
rect 2915 16745 2927 16748
rect 2869 16739 2927 16745
rect 3142 16736 3148 16748
rect 3200 16736 3206 16788
rect 3326 16776 3332 16788
rect 3287 16748 3332 16776
rect 3326 16736 3332 16748
rect 3384 16736 3390 16788
rect 5077 16779 5135 16785
rect 5077 16745 5089 16779
rect 5123 16776 5135 16779
rect 5166 16776 5172 16788
rect 5123 16748 5172 16776
rect 5123 16745 5135 16748
rect 5077 16739 5135 16745
rect 5166 16736 5172 16748
rect 5224 16736 5230 16788
rect 6270 16736 6276 16788
rect 6328 16776 6334 16788
rect 7926 16776 7932 16788
rect 6328 16748 7932 16776
rect 6328 16736 6334 16748
rect 7926 16736 7932 16748
rect 7984 16736 7990 16788
rect 8018 16736 8024 16788
rect 8076 16776 8082 16788
rect 11606 16776 11612 16788
rect 8076 16748 11612 16776
rect 8076 16736 8082 16748
rect 11606 16736 11612 16748
rect 11664 16736 11670 16788
rect 13630 16736 13636 16788
rect 13688 16776 13694 16788
rect 15289 16779 15347 16785
rect 13688 16748 14780 16776
rect 13688 16736 13694 16748
rect 1946 16708 1952 16720
rect 1907 16680 1952 16708
rect 1946 16668 1952 16680
rect 2004 16668 2010 16720
rect 2314 16668 2320 16720
rect 2372 16708 2378 16720
rect 2409 16711 2467 16717
rect 2409 16708 2421 16711
rect 2372 16680 2421 16708
rect 2372 16668 2378 16680
rect 2409 16677 2421 16680
rect 2455 16677 2467 16711
rect 2409 16671 2467 16677
rect 3234 16668 3240 16720
rect 3292 16708 3298 16720
rect 3421 16711 3479 16717
rect 3421 16708 3433 16711
rect 3292 16680 3433 16708
rect 3292 16668 3298 16680
rect 3421 16677 3433 16680
rect 3467 16677 3479 16711
rect 3421 16671 3479 16677
rect 3973 16711 4031 16717
rect 3973 16677 3985 16711
rect 4019 16677 4031 16711
rect 3973 16671 4031 16677
rect 4433 16711 4491 16717
rect 4433 16677 4445 16711
rect 4479 16708 4491 16711
rect 7742 16708 7748 16720
rect 4479 16680 5304 16708
rect 7703 16680 7748 16708
rect 4479 16677 4491 16680
rect 4433 16671 4491 16677
rect 2498 16600 2504 16652
rect 2556 16640 2562 16652
rect 3988 16640 4016 16671
rect 5276 16640 5304 16680
rect 7742 16668 7748 16680
rect 7800 16668 7806 16720
rect 8938 16708 8944 16720
rect 8899 16680 8944 16708
rect 8938 16668 8944 16680
rect 8996 16668 9002 16720
rect 9217 16711 9275 16717
rect 9217 16677 9229 16711
rect 9263 16708 9275 16711
rect 9306 16708 9312 16720
rect 9263 16680 9312 16708
rect 9263 16677 9275 16680
rect 9217 16671 9275 16677
rect 9306 16668 9312 16680
rect 9364 16668 9370 16720
rect 9582 16668 9588 16720
rect 9640 16708 9646 16720
rect 9640 16680 10272 16708
rect 9640 16668 9646 16680
rect 6549 16643 6607 16649
rect 2556 16612 3096 16640
rect 3988 16612 5028 16640
rect 5276 16612 6500 16640
rect 2556 16600 2562 16612
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16541 1823 16575
rect 2130 16572 2136 16584
rect 2091 16544 2136 16572
rect 1765 16535 1823 16541
rect 1780 16504 1808 16535
rect 2130 16532 2136 16544
rect 2188 16532 2194 16584
rect 2222 16532 2228 16584
rect 2280 16572 2286 16584
rect 3068 16581 3096 16612
rect 2777 16575 2835 16581
rect 2280 16544 2325 16572
rect 2280 16532 2286 16544
rect 2777 16541 2789 16575
rect 2823 16541 2835 16575
rect 2777 16535 2835 16541
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16541 3111 16575
rect 3053 16535 3111 16541
rect 3145 16575 3203 16581
rect 3145 16541 3157 16575
rect 3191 16572 3203 16575
rect 3234 16572 3240 16584
rect 3191 16544 3240 16572
rect 3191 16541 3203 16544
rect 3145 16535 3203 16541
rect 2682 16504 2688 16516
rect 1780 16476 2688 16504
rect 2682 16464 2688 16476
rect 2740 16464 2746 16516
rect 1394 16396 1400 16448
rect 1452 16436 1458 16448
rect 1581 16439 1639 16445
rect 1581 16436 1593 16439
rect 1452 16408 1593 16436
rect 1452 16396 1458 16408
rect 1581 16405 1593 16408
rect 1627 16405 1639 16439
rect 2792 16436 2820 16535
rect 3234 16532 3240 16544
rect 3292 16532 3298 16584
rect 3602 16572 3608 16584
rect 3563 16544 3608 16572
rect 3602 16532 3608 16544
rect 3660 16532 3666 16584
rect 3789 16575 3847 16581
rect 3789 16541 3801 16575
rect 3835 16572 3847 16575
rect 3878 16572 3884 16584
rect 3835 16544 3884 16572
rect 3835 16541 3847 16544
rect 3789 16535 3847 16541
rect 3878 16532 3884 16544
rect 3936 16532 3942 16584
rect 4062 16572 4068 16584
rect 4023 16544 4068 16572
rect 4062 16532 4068 16544
rect 4120 16532 4126 16584
rect 4522 16532 4528 16584
rect 4580 16572 4586 16584
rect 4617 16575 4675 16581
rect 4617 16572 4629 16575
rect 4580 16544 4629 16572
rect 4580 16532 4586 16544
rect 4617 16541 4629 16544
rect 4663 16541 4675 16575
rect 4893 16575 4951 16581
rect 4893 16572 4905 16575
rect 4617 16535 4675 16541
rect 4724 16544 4905 16572
rect 4154 16464 4160 16516
rect 4212 16504 4218 16516
rect 4724 16504 4752 16544
rect 4893 16541 4905 16544
rect 4939 16541 4951 16575
rect 5000 16572 5028 16612
rect 5169 16575 5227 16581
rect 5169 16572 5181 16575
rect 5000 16544 5181 16572
rect 4893 16535 4951 16541
rect 5169 16541 5181 16544
rect 5215 16541 5227 16575
rect 5169 16535 5227 16541
rect 5537 16575 5595 16581
rect 5537 16541 5549 16575
rect 5583 16541 5595 16575
rect 6472 16572 6500 16612
rect 6549 16609 6561 16643
rect 6595 16640 6607 16643
rect 7190 16640 7196 16652
rect 6595 16612 7196 16640
rect 6595 16609 6607 16612
rect 6549 16603 6607 16609
rect 7190 16600 7196 16612
rect 7248 16600 7254 16652
rect 7282 16600 7288 16652
rect 7340 16640 7346 16652
rect 7340 16612 7385 16640
rect 7340 16600 7346 16612
rect 8202 16600 8208 16652
rect 8260 16640 8266 16652
rect 8297 16643 8355 16649
rect 8297 16640 8309 16643
rect 8260 16612 8309 16640
rect 8260 16600 8266 16612
rect 8297 16609 8309 16612
rect 8343 16609 8355 16643
rect 10134 16640 10140 16652
rect 8297 16603 8355 16609
rect 8772 16612 8984 16640
rect 10095 16612 10140 16640
rect 7098 16572 7104 16584
rect 6472 16544 6868 16572
rect 7059 16544 7104 16572
rect 5537 16535 5595 16541
rect 5552 16504 5580 16535
rect 4212 16476 4752 16504
rect 4816 16476 5580 16504
rect 4212 16464 4218 16476
rect 3694 16436 3700 16448
rect 2792 16408 3700 16436
rect 1581 16399 1639 16405
rect 3694 16396 3700 16408
rect 3752 16396 3758 16448
rect 3970 16396 3976 16448
rect 4028 16436 4034 16448
rect 4816 16445 4844 16476
rect 5626 16464 5632 16516
rect 5684 16504 5690 16516
rect 6273 16507 6331 16513
rect 5684 16476 5948 16504
rect 5684 16464 5690 16476
rect 4249 16439 4307 16445
rect 4249 16436 4261 16439
rect 4028 16408 4261 16436
rect 4028 16396 4034 16408
rect 4249 16405 4261 16408
rect 4295 16405 4307 16439
rect 4249 16399 4307 16405
rect 4801 16439 4859 16445
rect 4801 16405 4813 16439
rect 4847 16405 4859 16439
rect 4801 16399 4859 16405
rect 5166 16396 5172 16448
rect 5224 16436 5230 16448
rect 5353 16439 5411 16445
rect 5353 16436 5365 16439
rect 5224 16408 5365 16436
rect 5224 16396 5230 16408
rect 5353 16405 5365 16408
rect 5399 16405 5411 16439
rect 5718 16436 5724 16448
rect 5679 16408 5724 16436
rect 5353 16399 5411 16405
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 5920 16445 5948 16476
rect 6273 16473 6285 16507
rect 6319 16504 6331 16507
rect 6319 16476 6776 16504
rect 6319 16473 6331 16476
rect 6273 16467 6331 16473
rect 5905 16439 5963 16445
rect 5905 16405 5917 16439
rect 5951 16405 5963 16439
rect 5905 16399 5963 16405
rect 6362 16396 6368 16448
rect 6420 16436 6426 16448
rect 6748 16445 6776 16476
rect 6733 16439 6791 16445
rect 6420 16408 6465 16436
rect 6420 16396 6426 16408
rect 6733 16405 6745 16439
rect 6779 16405 6791 16439
rect 6840 16436 6868 16544
rect 7098 16532 7104 16544
rect 7156 16532 7162 16584
rect 7374 16532 7380 16584
rect 7432 16572 7438 16584
rect 7561 16575 7619 16581
rect 7561 16572 7573 16575
rect 7432 16544 7573 16572
rect 7432 16532 7438 16544
rect 7561 16541 7573 16544
rect 7607 16541 7619 16575
rect 8573 16575 8631 16581
rect 8573 16572 8585 16575
rect 7561 16535 7619 16541
rect 7852 16544 8585 16572
rect 7193 16507 7251 16513
rect 7193 16473 7205 16507
rect 7239 16504 7251 16507
rect 7650 16504 7656 16516
rect 7239 16476 7656 16504
rect 7239 16473 7251 16476
rect 7193 16467 7251 16473
rect 7650 16464 7656 16476
rect 7708 16464 7714 16516
rect 7852 16436 7880 16544
rect 8573 16541 8585 16544
rect 8619 16572 8631 16575
rect 8772 16572 8800 16612
rect 8619 16544 8800 16572
rect 8619 16541 8631 16544
rect 8573 16535 8631 16541
rect 8846 16532 8852 16584
rect 8904 16532 8910 16584
rect 7926 16464 7932 16516
rect 7984 16504 7990 16516
rect 8864 16504 8892 16532
rect 7984 16476 8892 16504
rect 7984 16464 7990 16476
rect 8110 16436 8116 16448
rect 6840 16408 7880 16436
rect 8071 16408 8116 16436
rect 6733 16399 6791 16405
rect 8110 16396 8116 16408
rect 8168 16396 8174 16448
rect 8205 16439 8263 16445
rect 8205 16405 8217 16439
rect 8251 16436 8263 16439
rect 8386 16436 8392 16448
rect 8251 16408 8392 16436
rect 8251 16405 8263 16408
rect 8205 16399 8263 16405
rect 8386 16396 8392 16408
rect 8444 16396 8450 16448
rect 8757 16439 8815 16445
rect 8757 16405 8769 16439
rect 8803 16436 8815 16439
rect 8846 16436 8852 16448
rect 8803 16408 8852 16436
rect 8803 16405 8815 16408
rect 8757 16399 8815 16405
rect 8846 16396 8852 16408
rect 8904 16396 8910 16448
rect 8956 16436 8984 16612
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 10244 16649 10272 16680
rect 10778 16668 10784 16720
rect 10836 16708 10842 16720
rect 11287 16711 11345 16717
rect 11287 16708 11299 16711
rect 10836 16680 11299 16708
rect 10836 16668 10842 16680
rect 11287 16677 11299 16680
rect 11333 16708 11345 16711
rect 11977 16711 12035 16717
rect 11977 16708 11989 16711
rect 11333 16680 11989 16708
rect 11333 16677 11345 16680
rect 11287 16671 11345 16677
rect 11977 16677 11989 16680
rect 12023 16677 12035 16711
rect 11977 16671 12035 16677
rect 10229 16643 10287 16649
rect 10229 16609 10241 16643
rect 10275 16609 10287 16643
rect 10229 16603 10287 16609
rect 10318 16600 10324 16652
rect 10376 16640 10382 16652
rect 10689 16643 10747 16649
rect 10689 16640 10701 16643
rect 10376 16612 10701 16640
rect 10376 16600 10382 16612
rect 10689 16609 10701 16612
rect 10735 16609 10747 16643
rect 10689 16603 10747 16609
rect 11057 16643 11115 16649
rect 11057 16609 11069 16643
rect 11103 16609 11115 16643
rect 12710 16640 12716 16652
rect 12671 16612 12716 16640
rect 11057 16603 11115 16609
rect 9122 16572 9128 16584
rect 9083 16544 9128 16572
rect 9122 16532 9128 16544
rect 9180 16532 9186 16584
rect 9214 16532 9220 16584
rect 9272 16572 9278 16584
rect 9401 16575 9459 16581
rect 9401 16572 9413 16575
rect 9272 16544 9413 16572
rect 9272 16532 9278 16544
rect 9401 16541 9413 16544
rect 9447 16541 9459 16575
rect 9674 16572 9680 16584
rect 9401 16535 9459 16541
rect 9508 16544 9680 16572
rect 9306 16464 9312 16516
rect 9364 16504 9370 16516
rect 9508 16504 9536 16544
rect 9674 16532 9680 16544
rect 9732 16572 9738 16584
rect 10594 16572 10600 16584
rect 9732 16544 10600 16572
rect 9732 16532 9738 16544
rect 10594 16532 10600 16544
rect 10652 16532 10658 16584
rect 10962 16532 10968 16584
rect 11020 16572 11026 16584
rect 11072 16572 11100 16603
rect 12710 16600 12716 16612
rect 12768 16600 12774 16652
rect 12989 16643 13047 16649
rect 12989 16609 13001 16643
rect 13035 16640 13047 16643
rect 13262 16640 13268 16652
rect 13035 16612 13268 16640
rect 13035 16609 13047 16612
rect 12989 16603 13047 16609
rect 11514 16572 11520 16584
rect 11020 16544 11520 16572
rect 11020 16532 11026 16544
rect 11514 16532 11520 16544
rect 11572 16532 11578 16584
rect 12066 16532 12072 16584
rect 12124 16572 12130 16584
rect 13004 16572 13032 16603
rect 13262 16600 13268 16612
rect 13320 16600 13326 16652
rect 13446 16600 13452 16652
rect 13504 16640 13510 16652
rect 13504 16612 13584 16640
rect 13504 16600 13510 16612
rect 12124 16544 13032 16572
rect 13556 16572 13584 16612
rect 13814 16600 13820 16652
rect 13872 16640 13878 16652
rect 14642 16640 14648 16652
rect 13872 16612 13952 16640
rect 14603 16612 14648 16640
rect 13872 16600 13878 16612
rect 13924 16581 13952 16612
rect 14642 16600 14648 16612
rect 14700 16600 14706 16652
rect 14752 16640 14780 16748
rect 15289 16745 15301 16779
rect 15335 16776 15347 16779
rect 16298 16776 16304 16788
rect 15335 16748 16304 16776
rect 15335 16745 15347 16748
rect 15289 16739 15347 16745
rect 16298 16736 16304 16748
rect 16356 16736 16362 16788
rect 15286 16640 15292 16652
rect 14752 16612 14872 16640
rect 13633 16575 13691 16581
rect 13633 16572 13645 16575
rect 13556 16544 13645 16572
rect 12124 16532 12130 16544
rect 13633 16541 13645 16544
rect 13679 16541 13691 16575
rect 13633 16535 13691 16541
rect 13909 16575 13967 16581
rect 13909 16541 13921 16575
rect 13955 16541 13967 16575
rect 14844 16572 14872 16612
rect 15028 16612 15292 16640
rect 15028 16581 15056 16612
rect 15286 16600 15292 16612
rect 15344 16600 15350 16652
rect 14921 16575 14979 16581
rect 14921 16572 14933 16575
rect 14844 16544 14933 16572
rect 13909 16535 13967 16541
rect 14921 16541 14933 16544
rect 14967 16541 14979 16575
rect 14921 16535 14979 16541
rect 15013 16575 15071 16581
rect 15013 16541 15025 16575
rect 15059 16541 15071 16575
rect 15013 16535 15071 16541
rect 9364 16476 9536 16504
rect 10873 16507 10931 16513
rect 9364 16464 9370 16476
rect 10873 16473 10885 16507
rect 10919 16504 10931 16507
rect 11238 16504 11244 16516
rect 10919 16476 11244 16504
rect 10919 16473 10931 16476
rect 10873 16467 10931 16473
rect 11238 16464 11244 16476
rect 11296 16504 11302 16516
rect 15562 16504 15568 16516
rect 11296 16476 15568 16504
rect 11296 16464 11302 16476
rect 15562 16464 15568 16476
rect 15620 16464 15626 16516
rect 9490 16436 9496 16448
rect 8956 16408 9496 16436
rect 9490 16396 9496 16408
rect 9548 16396 9554 16448
rect 9674 16436 9680 16448
rect 9635 16408 9680 16436
rect 9674 16396 9680 16408
rect 9732 16396 9738 16448
rect 10042 16436 10048 16448
rect 10003 16408 10048 16436
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 10597 16439 10655 16445
rect 10597 16405 10609 16439
rect 10643 16436 10655 16439
rect 10962 16436 10968 16448
rect 10643 16408 10968 16436
rect 10643 16405 10655 16408
rect 10597 16399 10655 16405
rect 10962 16396 10968 16408
rect 11020 16396 11026 16448
rect 15470 16436 15476 16448
rect 15431 16408 15476 16436
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 1104 16346 16008 16368
rect 1104 16294 4698 16346
rect 4750 16294 4762 16346
rect 4814 16294 4826 16346
rect 4878 16294 4890 16346
rect 4942 16294 4954 16346
rect 5006 16294 8446 16346
rect 8498 16294 8510 16346
rect 8562 16294 8574 16346
rect 8626 16294 8638 16346
rect 8690 16294 8702 16346
rect 8754 16294 12194 16346
rect 12246 16294 12258 16346
rect 12310 16294 12322 16346
rect 12374 16294 12386 16346
rect 12438 16294 12450 16346
rect 12502 16294 16008 16346
rect 1104 16272 16008 16294
rect 2130 16232 2136 16244
rect 2091 16204 2136 16232
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 2409 16235 2467 16241
rect 2409 16201 2421 16235
rect 2455 16201 2467 16235
rect 2409 16195 2467 16201
rect 2961 16235 3019 16241
rect 2961 16201 2973 16235
rect 3007 16201 3019 16235
rect 2961 16195 3019 16201
rect 3697 16235 3755 16241
rect 3697 16201 3709 16235
rect 3743 16232 3755 16235
rect 4062 16232 4068 16244
rect 3743 16204 4068 16232
rect 3743 16201 3755 16204
rect 3697 16195 3755 16201
rect 2424 16164 2452 16195
rect 2056 16136 2452 16164
rect 2976 16164 3004 16195
rect 4062 16192 4068 16204
rect 4120 16192 4126 16244
rect 4246 16232 4252 16244
rect 4207 16204 4252 16232
rect 4246 16192 4252 16204
rect 4304 16192 4310 16244
rect 4893 16235 4951 16241
rect 4893 16201 4905 16235
rect 4939 16232 4951 16235
rect 5353 16235 5411 16241
rect 5353 16232 5365 16235
rect 4939 16204 5365 16232
rect 4939 16201 4951 16204
rect 4893 16195 4951 16201
rect 5353 16201 5365 16204
rect 5399 16201 5411 16235
rect 5353 16195 5411 16201
rect 5994 16192 6000 16244
rect 6052 16232 6058 16244
rect 6822 16232 6828 16244
rect 6052 16204 6828 16232
rect 6052 16192 6058 16204
rect 6822 16192 6828 16204
rect 6880 16192 6886 16244
rect 7742 16232 7748 16244
rect 7703 16204 7748 16232
rect 7742 16192 7748 16204
rect 7800 16192 7806 16244
rect 8110 16192 8116 16244
rect 8168 16192 8174 16244
rect 9033 16235 9091 16241
rect 9033 16201 9045 16235
rect 9079 16232 9091 16235
rect 9401 16235 9459 16241
rect 9401 16232 9413 16235
rect 9079 16204 9413 16232
rect 9079 16201 9091 16204
rect 9033 16195 9091 16201
rect 9401 16201 9413 16204
rect 9447 16201 9459 16235
rect 9401 16195 9459 16201
rect 9493 16235 9551 16241
rect 9493 16201 9505 16235
rect 9539 16232 9551 16235
rect 9953 16235 10011 16241
rect 9953 16232 9965 16235
rect 9539 16204 9965 16232
rect 9539 16201 9551 16204
rect 9493 16195 9551 16201
rect 9953 16201 9965 16204
rect 9999 16201 10011 16235
rect 9953 16195 10011 16201
rect 10042 16192 10048 16244
rect 10100 16232 10106 16244
rect 11517 16235 11575 16241
rect 11517 16232 11529 16235
rect 10100 16204 11529 16232
rect 10100 16192 10106 16204
rect 11517 16201 11529 16204
rect 11563 16201 11575 16235
rect 11517 16195 11575 16201
rect 11606 16192 11612 16244
rect 11664 16232 11670 16244
rect 11977 16235 12035 16241
rect 11977 16232 11989 16235
rect 11664 16204 11989 16232
rect 11664 16192 11670 16204
rect 11977 16201 11989 16204
rect 12023 16232 12035 16235
rect 12066 16232 12072 16244
rect 12023 16204 12072 16232
rect 12023 16201 12035 16204
rect 11977 16195 12035 16201
rect 12066 16192 12072 16204
rect 12124 16192 12130 16244
rect 13538 16232 13544 16244
rect 13499 16204 13544 16232
rect 13538 16192 13544 16204
rect 13596 16192 13602 16244
rect 14458 16192 14464 16244
rect 14516 16232 14522 16244
rect 16390 16232 16396 16244
rect 14516 16204 16396 16232
rect 14516 16192 14522 16204
rect 16390 16192 16396 16204
rect 16448 16192 16454 16244
rect 3970 16164 3976 16176
rect 2976 16136 3976 16164
rect 2056 16105 2084 16136
rect 3970 16124 3976 16136
rect 4028 16124 4034 16176
rect 4157 16167 4215 16173
rect 4157 16133 4169 16167
rect 4203 16164 4215 16167
rect 6733 16167 6791 16173
rect 6733 16164 6745 16167
rect 4203 16136 6745 16164
rect 4203 16133 4215 16136
rect 4157 16127 4215 16133
rect 6733 16133 6745 16136
rect 6779 16164 6791 16167
rect 6914 16164 6920 16176
rect 6779 16136 6920 16164
rect 6779 16133 6791 16136
rect 6733 16127 6791 16133
rect 6914 16124 6920 16136
rect 6972 16124 6978 16176
rect 7926 16164 7932 16176
rect 7208 16136 7932 16164
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16065 2099 16099
rect 2314 16096 2320 16108
rect 2275 16068 2320 16096
rect 2041 16059 2099 16065
rect 1688 16028 1716 16059
rect 2314 16056 2320 16068
rect 2372 16056 2378 16108
rect 2590 16096 2596 16108
rect 2551 16068 2596 16096
rect 2590 16056 2596 16068
rect 2648 16056 2654 16108
rect 2682 16056 2688 16108
rect 2740 16096 2746 16108
rect 2777 16099 2835 16105
rect 2777 16096 2789 16099
rect 2740 16068 2789 16096
rect 2740 16056 2746 16068
rect 2777 16065 2789 16068
rect 2823 16065 2835 16099
rect 3510 16096 3516 16108
rect 3471 16068 3516 16096
rect 2777 16059 2835 16065
rect 3510 16056 3516 16068
rect 3568 16056 3574 16108
rect 4338 16056 4344 16108
rect 4396 16096 4402 16108
rect 4433 16099 4491 16105
rect 4433 16096 4445 16099
rect 4396 16068 4445 16096
rect 4396 16056 4402 16068
rect 4433 16065 4445 16068
rect 4479 16096 4491 16099
rect 5258 16096 5264 16108
rect 4479 16068 5264 16096
rect 4479 16065 4491 16068
rect 4433 16059 4491 16065
rect 5258 16056 5264 16068
rect 5316 16056 5322 16108
rect 5718 16096 5724 16108
rect 5679 16068 5724 16096
rect 5718 16056 5724 16068
rect 5776 16056 5782 16108
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 6086 16096 6092 16108
rect 5859 16068 6092 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 6086 16056 6092 16068
rect 6144 16056 6150 16108
rect 7006 16056 7012 16108
rect 7064 16096 7070 16108
rect 7208 16105 7236 16136
rect 7926 16124 7932 16136
rect 7984 16124 7990 16176
rect 8128 16164 8156 16192
rect 9122 16164 9128 16176
rect 8128 16136 9128 16164
rect 9122 16124 9128 16136
rect 9180 16164 9186 16176
rect 9858 16164 9864 16176
rect 9180 16136 9864 16164
rect 9180 16124 9186 16136
rect 9858 16124 9864 16136
rect 9916 16124 9922 16176
rect 10502 16164 10508 16176
rect 10244 16136 10508 16164
rect 7193 16099 7251 16105
rect 7193 16096 7205 16099
rect 7064 16068 7205 16096
rect 7064 16056 7070 16068
rect 7193 16065 7205 16068
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 7837 16099 7895 16105
rect 7837 16065 7849 16099
rect 7883 16096 7895 16099
rect 8110 16096 8116 16108
rect 7883 16068 8116 16096
rect 7883 16065 7895 16068
rect 7837 16059 7895 16065
rect 8110 16056 8116 16068
rect 8168 16056 8174 16108
rect 8665 16099 8723 16105
rect 8665 16065 8677 16099
rect 8711 16096 8723 16099
rect 8938 16096 8944 16108
rect 8711 16068 8944 16096
rect 8711 16065 8723 16068
rect 8665 16059 8723 16065
rect 8938 16056 8944 16068
rect 8996 16056 9002 16108
rect 9490 16056 9496 16108
rect 9548 16096 9554 16108
rect 10244 16096 10272 16136
rect 10502 16124 10508 16136
rect 10560 16124 10566 16176
rect 10594 16124 10600 16176
rect 10652 16124 10658 16176
rect 10965 16167 11023 16173
rect 10965 16133 10977 16167
rect 11011 16164 11023 16167
rect 11885 16167 11943 16173
rect 11885 16164 11897 16167
rect 11011 16136 11897 16164
rect 11011 16133 11023 16136
rect 10965 16127 11023 16133
rect 11885 16133 11897 16136
rect 11931 16133 11943 16167
rect 11885 16127 11943 16133
rect 12802 16124 12808 16176
rect 12860 16164 12866 16176
rect 13357 16167 13415 16173
rect 13357 16164 13369 16167
rect 12860 16136 13369 16164
rect 12860 16124 12866 16136
rect 13357 16133 13369 16136
rect 13403 16164 13415 16167
rect 13446 16164 13452 16176
rect 13403 16136 13452 16164
rect 13403 16133 13415 16136
rect 13357 16127 13415 16133
rect 13446 16124 13452 16136
rect 13504 16124 13510 16176
rect 15654 16164 15660 16176
rect 15615 16136 15660 16164
rect 15654 16124 15660 16136
rect 15712 16124 15718 16176
rect 9548 16068 10272 16096
rect 10321 16099 10379 16105
rect 9548 16056 9554 16068
rect 10321 16065 10333 16099
rect 10367 16065 10379 16099
rect 10612 16096 10640 16124
rect 11057 16099 11115 16105
rect 11057 16096 11069 16099
rect 10612 16068 11069 16096
rect 10321 16059 10379 16065
rect 11057 16065 11069 16068
rect 11103 16065 11115 16099
rect 11057 16059 11115 16065
rect 3418 16028 3424 16040
rect 1688 16000 3424 16028
rect 3418 15988 3424 16000
rect 3476 15988 3482 16040
rect 3973 16031 4031 16037
rect 3973 15997 3985 16031
rect 4019 16028 4031 16031
rect 4062 16028 4068 16040
rect 4019 16000 4068 16028
rect 4019 15997 4031 16000
rect 3973 15991 4031 15997
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 4985 16031 5043 16037
rect 4985 15997 4997 16031
rect 5031 15997 5043 16031
rect 5166 16028 5172 16040
rect 5127 16000 5172 16028
rect 4985 15991 5043 15997
rect 1857 15963 1915 15969
rect 1857 15929 1869 15963
rect 1903 15960 1915 15963
rect 2774 15960 2780 15972
rect 1903 15932 2780 15960
rect 1903 15929 1915 15932
rect 1857 15923 1915 15929
rect 2774 15920 2780 15932
rect 2832 15920 2838 15972
rect 3329 15963 3387 15969
rect 3329 15929 3341 15963
rect 3375 15960 3387 15963
rect 4154 15960 4160 15972
rect 3375 15932 4160 15960
rect 3375 15929 3387 15932
rect 3329 15923 3387 15929
rect 4154 15920 4160 15932
rect 4212 15920 4218 15972
rect 5000 15960 5028 15991
rect 5166 15988 5172 16000
rect 5224 15988 5230 16040
rect 5902 15988 5908 16040
rect 5960 16028 5966 16040
rect 5997 16031 6055 16037
rect 5997 16028 6009 16031
rect 5960 16000 6009 16028
rect 5960 15988 5966 16000
rect 5997 15997 6009 16000
rect 6043 16028 6055 16031
rect 6917 16031 6975 16037
rect 6043 16000 6500 16028
rect 6043 15997 6055 16000
rect 5997 15991 6055 15997
rect 6365 15963 6423 15969
rect 6365 15960 6377 15963
rect 5000 15932 6377 15960
rect 6365 15929 6377 15932
rect 6411 15929 6423 15963
rect 6472 15960 6500 16000
rect 6917 15997 6929 16031
rect 6963 15997 6975 16031
rect 7650 16028 7656 16040
rect 7611 16000 7656 16028
rect 6917 15991 6975 15997
rect 6932 15960 6960 15991
rect 7650 15988 7656 16000
rect 7708 15988 7714 16040
rect 8478 16028 8484 16040
rect 8439 16000 8484 16028
rect 8478 15988 8484 16000
rect 8536 15988 8542 16040
rect 8573 16031 8631 16037
rect 8573 15997 8585 16031
rect 8619 16028 8631 16031
rect 8846 16028 8852 16040
rect 8619 16000 8852 16028
rect 8619 15997 8631 16000
rect 8573 15991 8631 15997
rect 8846 15988 8852 16000
rect 8904 15988 8910 16040
rect 9309 16031 9367 16037
rect 9309 15997 9321 16031
rect 9355 16028 9367 16031
rect 9582 16028 9588 16040
rect 9355 16000 9588 16028
rect 9355 15997 9367 16000
rect 9309 15991 9367 15997
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 9950 15988 9956 16040
rect 10008 16028 10014 16040
rect 10336 16028 10364 16059
rect 11330 16056 11336 16108
rect 11388 16096 11394 16108
rect 12713 16099 12771 16105
rect 12713 16096 12725 16099
rect 11388 16068 12725 16096
rect 11388 16056 11394 16068
rect 12713 16065 12725 16068
rect 12759 16065 12771 16099
rect 12713 16059 12771 16065
rect 12986 16056 12992 16108
rect 13044 16096 13050 16108
rect 13725 16099 13783 16105
rect 13725 16096 13737 16099
rect 13044 16068 13737 16096
rect 13044 16056 13050 16068
rect 13725 16065 13737 16068
rect 13771 16065 13783 16099
rect 13725 16059 13783 16065
rect 10008 16000 10364 16028
rect 10008 15988 10014 16000
rect 10410 15988 10416 16040
rect 10468 16028 10474 16040
rect 10597 16031 10655 16037
rect 10468 16000 10513 16028
rect 10468 15988 10474 16000
rect 10597 15997 10609 16031
rect 10643 16028 10655 16031
rect 12069 16031 12127 16037
rect 12069 16028 12081 16031
rect 10643 16000 12081 16028
rect 10643 15997 10655 16000
rect 10597 15991 10655 15997
rect 12069 15997 12081 16000
rect 12115 15997 12127 16031
rect 12069 15991 12127 15997
rect 8205 15963 8263 15969
rect 6472 15932 6960 15960
rect 7024 15932 7880 15960
rect 6365 15923 6423 15929
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 3237 15895 3295 15901
rect 3237 15861 3249 15895
rect 3283 15892 3295 15895
rect 4338 15892 4344 15904
rect 3283 15864 4344 15892
rect 3283 15861 3295 15864
rect 3237 15855 3295 15861
rect 4338 15852 4344 15864
rect 4396 15852 4402 15904
rect 4522 15892 4528 15904
rect 4483 15864 4528 15892
rect 4522 15852 4528 15864
rect 4580 15852 4586 15904
rect 5534 15852 5540 15904
rect 5592 15892 5598 15904
rect 7024 15892 7052 15932
rect 5592 15864 7052 15892
rect 7377 15895 7435 15901
rect 5592 15852 5598 15864
rect 7377 15861 7389 15895
rect 7423 15892 7435 15895
rect 7558 15892 7564 15904
rect 7423 15864 7564 15892
rect 7423 15861 7435 15864
rect 7377 15855 7435 15861
rect 7558 15852 7564 15864
rect 7616 15852 7622 15904
rect 7852 15892 7880 15932
rect 8205 15929 8217 15963
rect 8251 15960 8263 15963
rect 8251 15932 10364 15960
rect 8251 15929 8263 15932
rect 8205 15923 8263 15929
rect 8386 15892 8392 15904
rect 7852 15864 8392 15892
rect 8386 15852 8392 15864
rect 8444 15852 8450 15904
rect 8478 15852 8484 15904
rect 8536 15892 8542 15904
rect 9490 15892 9496 15904
rect 8536 15864 9496 15892
rect 8536 15852 8542 15864
rect 9490 15852 9496 15864
rect 9548 15852 9554 15904
rect 9861 15895 9919 15901
rect 9861 15861 9873 15895
rect 9907 15892 9919 15895
rect 9950 15892 9956 15904
rect 9907 15864 9956 15892
rect 9907 15861 9919 15864
rect 9861 15855 9919 15861
rect 9950 15852 9956 15864
rect 10008 15852 10014 15904
rect 10336 15892 10364 15932
rect 10502 15920 10508 15972
rect 10560 15960 10566 15972
rect 10612 15960 10640 15991
rect 12618 15988 12624 16040
rect 12676 16028 12682 16040
rect 12805 16031 12863 16037
rect 12805 16028 12817 16031
rect 12676 16000 12817 16028
rect 12676 15988 12682 16000
rect 12805 15997 12817 16000
rect 12851 15997 12863 16031
rect 12805 15991 12863 15997
rect 12897 16031 12955 16037
rect 12897 15997 12909 16031
rect 12943 15997 12955 16031
rect 13814 16028 13820 16040
rect 13775 16000 13820 16028
rect 12897 15991 12955 15997
rect 10560 15932 10640 15960
rect 10560 15920 10566 15932
rect 12526 15920 12532 15972
rect 12584 15960 12590 15972
rect 12912 15960 12940 15991
rect 13814 15988 13820 16000
rect 13872 15988 13878 16040
rect 14001 16031 14059 16037
rect 14001 15997 14013 16031
rect 14047 16028 14059 16031
rect 15470 16028 15476 16040
rect 14047 16000 15476 16028
rect 14047 15997 14059 16000
rect 14001 15991 14059 15997
rect 15470 15988 15476 16000
rect 15528 15988 15534 16040
rect 13170 15960 13176 15972
rect 12584 15932 12940 15960
rect 13131 15932 13176 15960
rect 12584 15920 12590 15932
rect 13170 15920 13176 15932
rect 13228 15920 13234 15972
rect 10686 15892 10692 15904
rect 10336 15864 10692 15892
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 11238 15892 11244 15904
rect 11199 15864 11244 15892
rect 11238 15852 11244 15864
rect 11296 15852 11302 15904
rect 12342 15892 12348 15904
rect 12303 15864 12348 15892
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 1104 15802 16008 15824
rect 1104 15750 2824 15802
rect 2876 15750 2888 15802
rect 2940 15750 2952 15802
rect 3004 15750 3016 15802
rect 3068 15750 3080 15802
rect 3132 15750 6572 15802
rect 6624 15750 6636 15802
rect 6688 15750 6700 15802
rect 6752 15750 6764 15802
rect 6816 15750 6828 15802
rect 6880 15750 10320 15802
rect 10372 15750 10384 15802
rect 10436 15750 10448 15802
rect 10500 15750 10512 15802
rect 10564 15750 10576 15802
rect 10628 15750 14068 15802
rect 14120 15750 14132 15802
rect 14184 15750 14196 15802
rect 14248 15750 14260 15802
rect 14312 15750 14324 15802
rect 14376 15750 16008 15802
rect 1104 15728 16008 15750
rect 1394 15688 1400 15700
rect 1355 15660 1400 15688
rect 1394 15648 1400 15660
rect 1452 15648 1458 15700
rect 1765 15691 1823 15697
rect 1765 15657 1777 15691
rect 1811 15688 1823 15691
rect 2222 15688 2228 15700
rect 1811 15660 2228 15688
rect 1811 15657 1823 15660
rect 1765 15651 1823 15657
rect 2222 15648 2228 15660
rect 2280 15648 2286 15700
rect 2406 15648 2412 15700
rect 2464 15688 2470 15700
rect 2501 15691 2559 15697
rect 2501 15688 2513 15691
rect 2464 15660 2513 15688
rect 2464 15648 2470 15660
rect 2501 15657 2513 15660
rect 2547 15657 2559 15691
rect 3418 15688 3424 15700
rect 3379 15660 3424 15688
rect 2501 15651 2559 15657
rect 3418 15648 3424 15660
rect 3476 15648 3482 15700
rect 4080 15660 4384 15688
rect 1412 15552 1440 15648
rect 2130 15580 2136 15632
rect 2188 15620 2194 15632
rect 2590 15620 2596 15632
rect 2188 15592 2596 15620
rect 2188 15580 2194 15592
rect 2590 15580 2596 15592
rect 2648 15580 2654 15632
rect 2774 15552 2780 15564
rect 1412 15524 1900 15552
rect 1872 15493 1900 15524
rect 2700 15524 2780 15552
rect 2700 15493 2728 15524
rect 2774 15512 2780 15524
rect 2832 15552 2838 15564
rect 3326 15552 3332 15564
rect 2832 15524 3332 15552
rect 2832 15512 2838 15524
rect 3326 15512 3332 15524
rect 3384 15512 3390 15564
rect 3878 15552 3884 15564
rect 3528 15524 3884 15552
rect 1581 15487 1639 15493
rect 1581 15453 1593 15487
rect 1627 15453 1639 15487
rect 1581 15447 1639 15453
rect 1857 15487 1915 15493
rect 1857 15453 1869 15487
rect 1903 15453 1915 15487
rect 1857 15447 1915 15453
rect 2685 15487 2743 15493
rect 2685 15453 2697 15487
rect 2731 15453 2743 15487
rect 2685 15447 2743 15453
rect 2961 15487 3019 15493
rect 2961 15453 2973 15487
rect 3007 15484 3019 15487
rect 3528 15484 3556 15524
rect 3878 15512 3884 15524
rect 3936 15552 3942 15564
rect 4080 15552 4108 15660
rect 4157 15623 4215 15629
rect 4157 15589 4169 15623
rect 4203 15589 4215 15623
rect 4356 15620 4384 15660
rect 4430 15648 4436 15700
rect 4488 15688 4494 15700
rect 4985 15691 5043 15697
rect 4985 15688 4997 15691
rect 4488 15660 4997 15688
rect 4488 15648 4494 15660
rect 4985 15657 4997 15660
rect 5031 15657 5043 15691
rect 5442 15688 5448 15700
rect 5403 15660 5448 15688
rect 4985 15651 5043 15657
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 5810 15688 5816 15700
rect 5771 15660 5816 15688
rect 5810 15648 5816 15660
rect 5868 15648 5874 15700
rect 6362 15688 6368 15700
rect 6323 15660 6368 15688
rect 6362 15648 6368 15660
rect 6420 15648 6426 15700
rect 7466 15688 7472 15700
rect 6472 15660 7472 15688
rect 5350 15620 5356 15632
rect 4356 15592 5356 15620
rect 4157 15583 4215 15589
rect 3936 15524 4108 15552
rect 3936 15512 3942 15524
rect 3007 15456 3556 15484
rect 3605 15487 3663 15493
rect 3007 15453 3019 15456
rect 2961 15447 3019 15453
rect 3605 15453 3617 15487
rect 3651 15484 3663 15487
rect 4172 15484 4200 15583
rect 5350 15580 5356 15592
rect 5408 15580 5414 15632
rect 6472 15620 6500 15660
rect 7466 15648 7472 15660
rect 7524 15648 7530 15700
rect 8938 15688 8944 15700
rect 7852 15660 8064 15688
rect 8899 15660 8944 15688
rect 7852 15620 7880 15660
rect 8036 15629 8064 15660
rect 8938 15648 8944 15660
rect 8996 15648 9002 15700
rect 10226 15688 10232 15700
rect 10187 15660 10232 15688
rect 10226 15648 10232 15660
rect 10284 15648 10290 15700
rect 11054 15648 11060 15700
rect 11112 15688 11118 15700
rect 12618 15688 12624 15700
rect 11112 15660 12480 15688
rect 12579 15660 12624 15688
rect 11112 15648 11118 15660
rect 5552 15592 6500 15620
rect 6748 15592 7880 15620
rect 7929 15623 7987 15629
rect 4246 15512 4252 15564
rect 4304 15552 4310 15564
rect 4801 15555 4859 15561
rect 4304 15524 4660 15552
rect 4304 15512 4310 15524
rect 4522 15484 4528 15496
rect 3651 15456 4200 15484
rect 4483 15456 4528 15484
rect 3651 15453 3663 15456
rect 3605 15447 3663 15453
rect 1596 15416 1624 15447
rect 4522 15444 4528 15456
rect 4580 15444 4586 15496
rect 4632 15484 4660 15524
rect 4801 15521 4813 15555
rect 4847 15552 4859 15555
rect 5442 15552 5448 15564
rect 4847 15524 5448 15552
rect 4847 15521 4859 15524
rect 4801 15515 4859 15521
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 5169 15487 5227 15493
rect 5169 15484 5181 15487
rect 4632 15456 5181 15484
rect 5169 15453 5181 15456
rect 5215 15484 5227 15487
rect 5552 15484 5580 15592
rect 5718 15552 5724 15564
rect 5679 15524 5724 15552
rect 5718 15512 5724 15524
rect 5776 15512 5782 15564
rect 6270 15552 6276 15564
rect 6231 15524 6276 15552
rect 6270 15512 6276 15524
rect 6328 15512 6334 15564
rect 5215 15456 5580 15484
rect 5215 15453 5227 15456
rect 5169 15447 5227 15453
rect 5810 15444 5816 15496
rect 5868 15484 5874 15496
rect 6748 15493 6776 15592
rect 7929 15589 7941 15623
rect 7975 15589 7987 15623
rect 7929 15583 7987 15589
rect 8021 15623 8079 15629
rect 8021 15589 8033 15623
rect 8067 15589 8079 15623
rect 8021 15583 8079 15589
rect 6917 15555 6975 15561
rect 6917 15552 6929 15555
rect 6840 15524 6929 15552
rect 5997 15487 6055 15493
rect 5997 15484 6009 15487
rect 5868 15456 6009 15484
rect 5868 15444 5874 15456
rect 5997 15453 6009 15456
rect 6043 15453 6055 15487
rect 5997 15447 6055 15453
rect 6733 15487 6791 15493
rect 6733 15453 6745 15487
rect 6779 15453 6791 15487
rect 6733 15447 6791 15453
rect 5626 15416 5632 15428
rect 1596 15388 5632 15416
rect 5626 15376 5632 15388
rect 5684 15376 5690 15428
rect 6086 15376 6092 15428
rect 6144 15416 6150 15428
rect 6840 15416 6868 15524
rect 6917 15521 6929 15524
rect 6963 15552 6975 15555
rect 7282 15552 7288 15564
rect 6963 15524 7288 15552
rect 6963 15521 6975 15524
rect 6917 15515 6975 15521
rect 7282 15512 7288 15524
rect 7340 15512 7346 15564
rect 7377 15555 7435 15561
rect 7377 15521 7389 15555
rect 7423 15552 7435 15555
rect 7834 15552 7840 15564
rect 7423 15524 7840 15552
rect 7423 15521 7435 15524
rect 7377 15515 7435 15521
rect 7834 15512 7840 15524
rect 7892 15512 7898 15564
rect 7944 15552 7972 15583
rect 8386 15580 8392 15632
rect 8444 15620 8450 15632
rect 12342 15620 12348 15632
rect 8444 15592 10916 15620
rect 8444 15580 8450 15592
rect 8481 15555 8539 15561
rect 8481 15552 8493 15555
rect 7944 15524 8493 15552
rect 8481 15521 8493 15524
rect 8527 15521 8539 15555
rect 8481 15515 8539 15521
rect 8573 15555 8631 15561
rect 8573 15521 8585 15555
rect 8619 15521 8631 15555
rect 8573 15515 8631 15521
rect 7098 15444 7104 15496
rect 7156 15484 7162 15496
rect 8202 15484 8208 15496
rect 7156 15456 8208 15484
rect 7156 15444 7162 15456
rect 8202 15444 8208 15456
rect 8260 15484 8266 15496
rect 8588 15484 8616 15515
rect 9398 15512 9404 15564
rect 9456 15552 9462 15564
rect 9493 15555 9551 15561
rect 9493 15552 9505 15555
rect 9456 15524 9505 15552
rect 9456 15512 9462 15524
rect 9493 15521 9505 15524
rect 9539 15552 9551 15555
rect 10781 15555 10839 15561
rect 10781 15552 10793 15555
rect 9539 15524 10793 15552
rect 9539 15521 9551 15524
rect 9493 15515 9551 15521
rect 10781 15521 10793 15524
rect 10827 15521 10839 15555
rect 10781 15515 10839 15521
rect 8260 15456 8616 15484
rect 8260 15444 8266 15456
rect 9030 15444 9036 15496
rect 9088 15484 9094 15496
rect 9309 15487 9367 15493
rect 9309 15484 9321 15487
rect 9088 15456 9321 15484
rect 9088 15444 9094 15456
rect 9309 15453 9321 15456
rect 9355 15453 9367 15487
rect 9309 15447 9367 15453
rect 9769 15487 9827 15493
rect 9769 15453 9781 15487
rect 9815 15484 9827 15487
rect 9858 15484 9864 15496
rect 9815 15456 9864 15484
rect 9815 15453 9827 15456
rect 9769 15447 9827 15453
rect 9858 15444 9864 15456
rect 9916 15484 9922 15496
rect 10045 15487 10103 15493
rect 10045 15484 10057 15487
rect 9916 15456 10057 15484
rect 9916 15444 9922 15456
rect 10045 15453 10057 15456
rect 10091 15453 10103 15487
rect 10045 15447 10103 15453
rect 10689 15487 10747 15493
rect 10689 15453 10701 15487
rect 10735 15484 10747 15487
rect 10888 15484 10916 15592
rect 11532 15592 12348 15620
rect 11532 15561 11560 15592
rect 12342 15580 12348 15592
rect 12400 15580 12406 15632
rect 12452 15620 12480 15660
rect 12618 15648 12624 15660
rect 12676 15648 12682 15700
rect 13725 15623 13783 15629
rect 13725 15620 13737 15623
rect 12452 15592 13737 15620
rect 13725 15589 13737 15592
rect 13771 15589 13783 15623
rect 13725 15583 13783 15589
rect 11517 15555 11575 15561
rect 11517 15521 11529 15555
rect 11563 15521 11575 15555
rect 11517 15515 11575 15521
rect 11609 15555 11667 15561
rect 11609 15521 11621 15555
rect 11655 15521 11667 15555
rect 11609 15515 11667 15521
rect 10962 15484 10968 15496
rect 10735 15456 10968 15484
rect 10735 15453 10747 15456
rect 10689 15447 10747 15453
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 11054 15444 11060 15496
rect 11112 15484 11118 15496
rect 11624 15484 11652 15515
rect 11790 15512 11796 15564
rect 11848 15552 11854 15564
rect 11977 15555 12035 15561
rect 11977 15552 11989 15555
rect 11848 15524 11989 15552
rect 11848 15512 11854 15524
rect 11977 15521 11989 15524
rect 12023 15521 12035 15555
rect 11977 15515 12035 15521
rect 12066 15512 12072 15564
rect 12124 15552 12130 15564
rect 12124 15524 12434 15552
rect 12124 15512 12130 15524
rect 11112 15456 11652 15484
rect 11112 15444 11118 15456
rect 11882 15444 11888 15496
rect 11940 15484 11946 15496
rect 12253 15487 12311 15493
rect 12253 15484 12265 15487
rect 11940 15456 12265 15484
rect 11940 15444 11946 15456
rect 12253 15453 12265 15456
rect 12299 15453 12311 15487
rect 12406 15484 12434 15524
rect 12894 15512 12900 15564
rect 12952 15552 12958 15564
rect 12989 15555 13047 15561
rect 12989 15552 13001 15555
rect 12952 15524 13001 15552
rect 12952 15512 12958 15524
rect 12989 15521 13001 15524
rect 13035 15521 13047 15555
rect 14274 15552 14280 15564
rect 12989 15515 13047 15521
rect 13188 15524 14280 15552
rect 12710 15484 12716 15496
rect 12406 15456 12716 15484
rect 12253 15447 12311 15453
rect 12710 15444 12716 15456
rect 12768 15484 12774 15496
rect 13188 15484 13216 15524
rect 14274 15512 14280 15524
rect 14332 15512 14338 15564
rect 14829 15555 14887 15561
rect 14829 15521 14841 15555
rect 14875 15552 14887 15555
rect 15010 15552 15016 15564
rect 14875 15524 15016 15552
rect 14875 15521 14887 15524
rect 14829 15515 14887 15521
rect 15010 15512 15016 15524
rect 15068 15552 15074 15564
rect 15286 15552 15292 15564
rect 15068 15524 15292 15552
rect 15068 15512 15074 15524
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 13909 15487 13967 15493
rect 13909 15484 13921 15487
rect 12768 15456 13216 15484
rect 13832 15456 13921 15484
rect 12768 15444 12774 15456
rect 6144 15388 6868 15416
rect 6144 15376 6150 15388
rect 7374 15376 7380 15428
rect 7432 15416 7438 15428
rect 7561 15419 7619 15425
rect 7561 15416 7573 15419
rect 7432 15388 7573 15416
rect 7432 15376 7438 15388
rect 7561 15385 7573 15388
rect 7607 15385 7619 15419
rect 10502 15416 10508 15428
rect 7561 15379 7619 15385
rect 9968 15388 10508 15416
rect 2038 15348 2044 15360
rect 1999 15320 2044 15348
rect 2038 15308 2044 15320
rect 2096 15308 2102 15360
rect 2130 15308 2136 15360
rect 2188 15348 2194 15360
rect 2406 15348 2412 15360
rect 2188 15320 2233 15348
rect 2367 15320 2412 15348
rect 2188 15308 2194 15320
rect 2406 15308 2412 15320
rect 2464 15308 2470 15360
rect 2774 15308 2780 15360
rect 2832 15348 2838 15360
rect 3050 15348 3056 15360
rect 2832 15320 3056 15348
rect 2832 15308 2838 15320
rect 3050 15308 3056 15320
rect 3108 15308 3114 15360
rect 3329 15351 3387 15357
rect 3329 15317 3341 15351
rect 3375 15348 3387 15351
rect 3418 15348 3424 15360
rect 3375 15320 3424 15348
rect 3375 15317 3387 15320
rect 3329 15311 3387 15317
rect 3418 15308 3424 15320
rect 3476 15308 3482 15360
rect 3786 15348 3792 15360
rect 3747 15320 3792 15348
rect 3786 15308 3792 15320
rect 3844 15308 3850 15360
rect 4614 15348 4620 15360
rect 4575 15320 4620 15348
rect 4614 15308 4620 15320
rect 4672 15308 4678 15360
rect 6822 15308 6828 15360
rect 6880 15348 6886 15360
rect 7466 15348 7472 15360
rect 6880 15320 6925 15348
rect 7427 15320 7472 15348
rect 6880 15308 6886 15320
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 8202 15308 8208 15360
rect 8260 15348 8266 15360
rect 8386 15348 8392 15360
rect 8260 15320 8392 15348
rect 8260 15308 8266 15320
rect 8386 15308 8392 15320
rect 8444 15308 8450 15360
rect 8938 15308 8944 15360
rect 8996 15348 9002 15360
rect 9968 15357 9996 15388
rect 10502 15376 10508 15388
rect 10560 15376 10566 15428
rect 10778 15416 10784 15428
rect 10612 15388 10784 15416
rect 9401 15351 9459 15357
rect 9401 15348 9413 15351
rect 8996 15320 9413 15348
rect 8996 15308 9002 15320
rect 9401 15317 9413 15320
rect 9447 15317 9459 15351
rect 9401 15311 9459 15317
rect 9953 15351 10011 15357
rect 9953 15317 9965 15351
rect 9999 15317 10011 15351
rect 9953 15311 10011 15317
rect 10226 15308 10232 15360
rect 10284 15348 10290 15360
rect 10612 15357 10640 15388
rect 10778 15376 10784 15388
rect 10836 15376 10842 15428
rect 11974 15376 11980 15428
rect 12032 15416 12038 15428
rect 13173 15419 13231 15425
rect 13173 15416 13185 15419
rect 12032 15388 13185 15416
rect 12032 15376 12038 15388
rect 13173 15385 13185 15388
rect 13219 15385 13231 15419
rect 13173 15379 13231 15385
rect 13265 15419 13323 15425
rect 13265 15385 13277 15419
rect 13311 15416 13323 15419
rect 13538 15416 13544 15428
rect 13311 15388 13544 15416
rect 13311 15385 13323 15388
rect 13265 15379 13323 15385
rect 13538 15376 13544 15388
rect 13596 15376 13602 15428
rect 13832 15360 13860 15456
rect 13909 15453 13921 15456
rect 13955 15453 13967 15487
rect 13909 15447 13967 15453
rect 14550 15444 14556 15496
rect 14608 15484 14614 15496
rect 14645 15487 14703 15493
rect 14645 15484 14657 15487
rect 14608 15456 14657 15484
rect 14608 15444 14614 15456
rect 14645 15453 14657 15456
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 13998 15376 14004 15428
rect 14056 15416 14062 15428
rect 14277 15419 14335 15425
rect 14277 15416 14289 15419
rect 14056 15388 14289 15416
rect 14056 15376 14062 15388
rect 14277 15385 14289 15388
rect 14323 15416 14335 15419
rect 14458 15416 14464 15428
rect 14323 15388 14464 15416
rect 14323 15385 14335 15388
rect 14277 15379 14335 15385
rect 14458 15376 14464 15388
rect 14516 15376 14522 15428
rect 14660 15416 14688 15447
rect 14734 15444 14740 15496
rect 14792 15484 14798 15496
rect 15105 15487 15163 15493
rect 15105 15484 15117 15487
rect 14792 15456 15117 15484
rect 14792 15444 14798 15456
rect 15105 15453 15117 15456
rect 15151 15453 15163 15487
rect 15105 15447 15163 15453
rect 14918 15416 14924 15428
rect 14660 15388 14924 15416
rect 14918 15376 14924 15388
rect 14976 15376 14982 15428
rect 10597 15351 10655 15357
rect 10597 15348 10609 15351
rect 10284 15320 10609 15348
rect 10284 15308 10290 15320
rect 10597 15317 10609 15320
rect 10643 15317 10655 15351
rect 10597 15311 10655 15317
rect 11057 15351 11115 15357
rect 11057 15317 11069 15351
rect 11103 15348 11115 15351
rect 11146 15348 11152 15360
rect 11103 15320 11152 15348
rect 11103 15317 11115 15320
rect 11057 15311 11115 15317
rect 11146 15308 11152 15320
rect 11204 15308 11210 15360
rect 11422 15348 11428 15360
rect 11383 15320 11428 15348
rect 11422 15308 11428 15320
rect 11480 15308 11486 15360
rect 12066 15308 12072 15360
rect 12124 15348 12130 15360
rect 12161 15351 12219 15357
rect 12161 15348 12173 15351
rect 12124 15320 12173 15348
rect 12124 15308 12130 15320
rect 12161 15317 12173 15320
rect 12207 15317 12219 15351
rect 12802 15348 12808 15360
rect 12763 15320 12808 15348
rect 12161 15311 12219 15317
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 13630 15348 13636 15360
rect 13591 15320 13636 15348
rect 13630 15308 13636 15320
rect 13688 15308 13694 15360
rect 13814 15308 13820 15360
rect 13872 15308 13878 15360
rect 13906 15308 13912 15360
rect 13964 15348 13970 15360
rect 14185 15351 14243 15357
rect 14185 15348 14197 15351
rect 13964 15320 14197 15348
rect 13964 15308 13970 15320
rect 14185 15317 14197 15320
rect 14231 15317 14243 15351
rect 14550 15348 14556 15360
rect 14511 15320 14556 15348
rect 14185 15311 14243 15317
rect 14550 15308 14556 15320
rect 14608 15308 14614 15360
rect 1104 15258 16008 15280
rect 1104 15206 4698 15258
rect 4750 15206 4762 15258
rect 4814 15206 4826 15258
rect 4878 15206 4890 15258
rect 4942 15206 4954 15258
rect 5006 15206 8446 15258
rect 8498 15206 8510 15258
rect 8562 15206 8574 15258
rect 8626 15206 8638 15258
rect 8690 15206 8702 15258
rect 8754 15206 12194 15258
rect 12246 15206 12258 15258
rect 12310 15206 12322 15258
rect 12374 15206 12386 15258
rect 12438 15206 12450 15258
rect 12502 15206 16008 15258
rect 1104 15184 16008 15206
rect 3053 15147 3111 15153
rect 3053 15113 3065 15147
rect 3099 15144 3111 15147
rect 3418 15144 3424 15156
rect 3099 15116 3424 15144
rect 3099 15113 3111 15116
rect 3053 15107 3111 15113
rect 3418 15104 3424 15116
rect 3476 15104 3482 15156
rect 3513 15147 3571 15153
rect 3513 15113 3525 15147
rect 3559 15144 3571 15147
rect 3786 15144 3792 15156
rect 3559 15116 3792 15144
rect 3559 15113 3571 15116
rect 3513 15107 3571 15113
rect 3786 15104 3792 15116
rect 3844 15104 3850 15156
rect 4157 15147 4215 15153
rect 4157 15113 4169 15147
rect 4203 15113 4215 15147
rect 4157 15107 4215 15113
rect 4433 15147 4491 15153
rect 4433 15113 4445 15147
rect 4479 15144 4491 15147
rect 4614 15144 4620 15156
rect 4479 15116 4620 15144
rect 4479 15113 4491 15116
rect 4433 15107 4491 15113
rect 2501 15079 2559 15085
rect 2501 15045 2513 15079
rect 2547 15076 2559 15079
rect 2547 15048 2774 15076
rect 2547 15045 2559 15048
rect 2501 15039 2559 15045
rect 1578 14968 1584 15020
rect 1636 15008 1642 15020
rect 1673 15011 1731 15017
rect 1673 15008 1685 15011
rect 1636 14980 1685 15008
rect 1636 14968 1642 14980
rect 1673 14977 1685 14980
rect 1719 14977 1731 15011
rect 1946 15008 1952 15020
rect 1907 14980 1952 15008
rect 1673 14971 1731 14977
rect 1946 14968 1952 14980
rect 2004 14968 2010 15020
rect 2746 15008 2774 15048
rect 3142 15036 3148 15088
rect 3200 15076 3206 15088
rect 4172 15076 4200 15107
rect 4614 15104 4620 15116
rect 4672 15104 4678 15156
rect 4893 15147 4951 15153
rect 4893 15113 4905 15147
rect 4939 15144 4951 15147
rect 5261 15147 5319 15153
rect 5261 15144 5273 15147
rect 4939 15116 5273 15144
rect 4939 15113 4951 15116
rect 4893 15107 4951 15113
rect 5261 15113 5273 15116
rect 5307 15113 5319 15147
rect 5261 15107 5319 15113
rect 5350 15104 5356 15156
rect 5408 15144 5414 15156
rect 5408 15116 5764 15144
rect 5408 15104 5414 15116
rect 5629 15079 5687 15085
rect 5629 15076 5641 15079
rect 3200 15048 4200 15076
rect 4724 15048 5641 15076
rect 3200 15036 3206 15048
rect 3694 15008 3700 15020
rect 2746 14980 3700 15008
rect 3694 14968 3700 14980
rect 3752 14968 3758 15020
rect 4065 15011 4123 15017
rect 4065 14977 4077 15011
rect 4111 15008 4123 15011
rect 4246 15008 4252 15020
rect 4111 14980 4252 15008
rect 4111 14977 4123 14980
rect 4065 14971 4123 14977
rect 4246 14968 4252 14980
rect 4304 14968 4310 15020
rect 4341 15011 4399 15017
rect 4341 14977 4353 15011
rect 4387 15008 4399 15011
rect 4430 15008 4436 15020
rect 4387 14980 4436 15008
rect 4387 14977 4399 14980
rect 4341 14971 4399 14977
rect 4430 14968 4436 14980
rect 4488 14968 4494 15020
rect 3418 14900 3424 14952
rect 3476 14940 3482 14952
rect 3602 14940 3608 14952
rect 3476 14912 3608 14940
rect 3476 14900 3482 14912
rect 3602 14900 3608 14912
rect 3660 14900 3666 14952
rect 3786 14940 3792 14952
rect 3747 14912 3792 14940
rect 3786 14900 3792 14912
rect 3844 14900 3850 14952
rect 3970 14900 3976 14952
rect 4028 14940 4034 14952
rect 4724 14940 4752 15048
rect 5629 15045 5641 15048
rect 5675 15045 5687 15079
rect 5736 15076 5764 15116
rect 5994 15104 6000 15156
rect 6052 15144 6058 15156
rect 6365 15147 6423 15153
rect 6365 15144 6377 15147
rect 6052 15116 6377 15144
rect 6052 15104 6058 15116
rect 6365 15113 6377 15116
rect 6411 15113 6423 15147
rect 6365 15107 6423 15113
rect 6549 15147 6607 15153
rect 6549 15113 6561 15147
rect 6595 15144 6607 15147
rect 6822 15144 6828 15156
rect 6595 15116 6828 15144
rect 6595 15113 6607 15116
rect 6549 15107 6607 15113
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 7009 15147 7067 15153
rect 7009 15113 7021 15147
rect 7055 15144 7067 15147
rect 7377 15147 7435 15153
rect 7377 15144 7389 15147
rect 7055 15116 7389 15144
rect 7055 15113 7067 15116
rect 7009 15107 7067 15113
rect 7377 15113 7389 15116
rect 7423 15113 7435 15147
rect 7377 15107 7435 15113
rect 7558 15104 7564 15156
rect 7616 15144 7622 15156
rect 7742 15144 7748 15156
rect 7616 15116 7748 15144
rect 7616 15104 7622 15116
rect 7742 15104 7748 15116
rect 7800 15104 7806 15156
rect 8665 15147 8723 15153
rect 8665 15113 8677 15147
rect 8711 15144 8723 15147
rect 8846 15144 8852 15156
rect 8711 15116 8852 15144
rect 8711 15113 8723 15116
rect 8665 15107 8723 15113
rect 8846 15104 8852 15116
rect 8904 15104 8910 15156
rect 9398 15144 9404 15156
rect 9324 15116 9404 15144
rect 6178 15076 6184 15088
rect 5736 15048 6184 15076
rect 5629 15039 5687 15045
rect 4801 15011 4859 15017
rect 4801 14977 4813 15011
rect 4847 15008 4859 15011
rect 5074 15008 5080 15020
rect 4847 14980 5080 15008
rect 4847 14977 4859 14980
rect 4801 14971 4859 14977
rect 5074 14968 5080 14980
rect 5132 14968 5138 15020
rect 5644 15008 5672 15039
rect 6178 15036 6184 15048
rect 6236 15036 6242 15088
rect 6454 15036 6460 15088
rect 6512 15076 6518 15088
rect 7650 15076 7656 15088
rect 6512 15048 7656 15076
rect 6512 15036 6518 15048
rect 7650 15036 7656 15048
rect 7708 15036 7714 15088
rect 8110 15036 8116 15088
rect 8168 15076 8174 15088
rect 8754 15076 8760 15088
rect 8168 15048 8760 15076
rect 8168 15036 8174 15048
rect 8754 15036 8760 15048
rect 8812 15036 8818 15088
rect 6822 15008 6828 15020
rect 5644 14980 6828 15008
rect 6822 14968 6828 14980
rect 6880 14968 6886 15020
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 15008 6975 15011
rect 7282 15008 7288 15020
rect 6963 14980 7288 15008
rect 6963 14977 6975 14980
rect 6917 14971 6975 14977
rect 7282 14968 7288 14980
rect 7340 14968 7346 15020
rect 7742 14968 7748 15020
rect 7800 15012 7806 15020
rect 7800 15008 7972 15012
rect 8202 15008 8208 15020
rect 7800 14984 8208 15008
rect 7800 14968 7806 14984
rect 7944 14980 8208 14984
rect 8202 14968 8208 14980
rect 8260 15008 8266 15020
rect 8389 15011 8447 15017
rect 8389 15008 8401 15011
rect 8260 14980 8401 15008
rect 8260 14968 8266 14980
rect 8389 14977 8401 14980
rect 8435 15008 8447 15011
rect 9033 15011 9091 15017
rect 9033 15008 9045 15011
rect 8435 14980 9045 15008
rect 8435 14977 8447 14980
rect 8389 14971 8447 14977
rect 9033 14977 9045 14980
rect 9079 14977 9091 15011
rect 9033 14971 9091 14977
rect 9324 14952 9352 15116
rect 9398 15104 9404 15116
rect 9456 15104 9462 15156
rect 9674 15104 9680 15156
rect 9732 15144 9738 15156
rect 9861 15147 9919 15153
rect 9861 15144 9873 15147
rect 9732 15116 9873 15144
rect 9732 15104 9738 15116
rect 9861 15113 9873 15116
rect 9907 15113 9919 15147
rect 9861 15107 9919 15113
rect 9950 15104 9956 15156
rect 10008 15144 10014 15156
rect 10008 15116 10053 15144
rect 10008 15104 10014 15116
rect 10134 15104 10140 15156
rect 10192 15144 10198 15156
rect 10410 15144 10416 15156
rect 10192 15116 10416 15144
rect 10192 15104 10198 15116
rect 10410 15104 10416 15116
rect 10468 15144 10474 15156
rect 11330 15144 11336 15156
rect 10468 15116 11100 15144
rect 11291 15116 11336 15144
rect 10468 15104 10474 15116
rect 10962 15076 10968 15088
rect 10923 15048 10968 15076
rect 10962 15036 10968 15048
rect 11020 15036 11026 15088
rect 11072 15076 11100 15116
rect 11330 15104 11336 15116
rect 11388 15104 11394 15156
rect 11885 15147 11943 15153
rect 11885 15144 11897 15147
rect 11440 15116 11897 15144
rect 11440 15076 11468 15116
rect 11885 15113 11897 15116
rect 11931 15113 11943 15147
rect 11885 15107 11943 15113
rect 12066 15104 12072 15156
rect 12124 15144 12130 15156
rect 12345 15147 12403 15153
rect 12345 15144 12357 15147
rect 12124 15116 12357 15144
rect 12124 15104 12130 15116
rect 12345 15113 12357 15116
rect 12391 15113 12403 15147
rect 12345 15107 12403 15113
rect 12452 15116 12848 15144
rect 11072 15048 11468 15076
rect 11790 15036 11796 15088
rect 11848 15076 11854 15088
rect 12452 15076 12480 15116
rect 11848 15048 12480 15076
rect 12820 15076 12848 15116
rect 13630 15104 13636 15156
rect 13688 15144 13694 15156
rect 13725 15147 13783 15153
rect 13725 15144 13737 15147
rect 13688 15116 13737 15144
rect 13688 15104 13694 15116
rect 13725 15113 13737 15116
rect 13771 15113 13783 15147
rect 13725 15107 13783 15113
rect 14093 15147 14151 15153
rect 14093 15113 14105 15147
rect 14139 15144 14151 15147
rect 14550 15144 14556 15156
rect 14139 15116 14556 15144
rect 14139 15113 14151 15116
rect 14093 15107 14151 15113
rect 14550 15104 14556 15116
rect 14608 15104 14614 15156
rect 15562 15144 15568 15156
rect 15523 15116 15568 15144
rect 15562 15104 15568 15116
rect 15620 15104 15626 15156
rect 13173 15079 13231 15085
rect 13173 15076 13185 15079
rect 12820 15048 13185 15076
rect 11848 15036 11854 15048
rect 13173 15045 13185 15048
rect 13219 15045 13231 15079
rect 13173 15039 13231 15045
rect 14461 15079 14519 15085
rect 14461 15045 14473 15079
rect 14507 15076 14519 15079
rect 14826 15076 14832 15088
rect 14507 15048 14832 15076
rect 14507 15045 14519 15048
rect 14461 15039 14519 15045
rect 14826 15036 14832 15048
rect 14884 15076 14890 15088
rect 15838 15076 15844 15088
rect 14884 15048 15844 15076
rect 14884 15036 14890 15048
rect 15838 15036 15844 15048
rect 15896 15036 15902 15088
rect 10873 15011 10931 15017
rect 10873 14977 10885 15011
rect 10919 15008 10931 15011
rect 11238 15008 11244 15020
rect 10919 14980 11244 15008
rect 10919 14977 10931 14980
rect 10873 14971 10931 14977
rect 11238 14968 11244 14980
rect 11296 15008 11302 15020
rect 11900 15008 12112 15012
rect 11296 14984 12112 15008
rect 11296 14980 11928 14984
rect 11296 14968 11302 14980
rect 12084 14952 12112 14984
rect 12434 14968 12440 15020
rect 12492 15008 12498 15020
rect 12713 15011 12771 15017
rect 12713 15008 12725 15011
rect 12492 14980 12725 15008
rect 12492 14968 12498 14980
rect 12713 14977 12725 14980
rect 12759 14977 12771 15011
rect 12713 14971 12771 14977
rect 12805 15011 12863 15017
rect 12805 14977 12817 15011
rect 12851 15008 12863 15011
rect 14274 15008 14280 15020
rect 12851 14980 14136 15008
rect 14235 14980 14280 15008
rect 12851 14977 12863 14980
rect 12805 14971 12863 14977
rect 4028 14912 4752 14940
rect 4985 14943 5043 14949
rect 4028 14900 4034 14912
rect 4985 14909 4997 14943
rect 5031 14940 5043 14943
rect 5166 14940 5172 14952
rect 5031 14912 5172 14940
rect 5031 14909 5043 14912
rect 4985 14903 5043 14909
rect 5166 14900 5172 14912
rect 5224 14900 5230 14952
rect 5718 14940 5724 14952
rect 5679 14912 5724 14940
rect 5718 14900 5724 14912
rect 5776 14900 5782 14952
rect 5902 14940 5908 14952
rect 5863 14912 5908 14940
rect 5902 14900 5908 14912
rect 5960 14900 5966 14952
rect 7098 14940 7104 14952
rect 7059 14912 7104 14940
rect 7098 14900 7104 14912
rect 7156 14900 7162 14952
rect 7558 14900 7564 14952
rect 7616 14940 7622 14952
rect 7837 14943 7895 14949
rect 7837 14940 7849 14943
rect 7616 14912 7849 14940
rect 7616 14900 7622 14912
rect 7837 14909 7849 14912
rect 7883 14909 7895 14943
rect 7837 14903 7895 14909
rect 8021 14943 8079 14949
rect 8021 14909 8033 14943
rect 8067 14909 8079 14943
rect 8021 14903 8079 14909
rect 2406 14832 2412 14884
rect 2464 14872 2470 14884
rect 2869 14875 2927 14881
rect 2869 14872 2881 14875
rect 2464 14844 2881 14872
rect 2464 14832 2470 14844
rect 2869 14841 2881 14844
rect 2915 14872 2927 14875
rect 3234 14872 3240 14884
rect 2915 14844 3240 14872
rect 2915 14841 2927 14844
rect 2869 14835 2927 14841
rect 3234 14832 3240 14844
rect 3292 14872 3298 14884
rect 5534 14872 5540 14884
rect 3292 14844 5540 14872
rect 3292 14832 3298 14844
rect 5534 14832 5540 14844
rect 5592 14832 5598 14884
rect 5626 14832 5632 14884
rect 5684 14872 5690 14884
rect 7742 14872 7748 14884
rect 5684 14844 7748 14872
rect 5684 14832 5690 14844
rect 7742 14832 7748 14844
rect 7800 14832 7806 14884
rect 7926 14832 7932 14884
rect 7984 14872 7990 14884
rect 8036 14872 8064 14903
rect 8110 14900 8116 14952
rect 8168 14940 8174 14952
rect 9125 14943 9183 14949
rect 9125 14940 9137 14943
rect 8168 14912 9137 14940
rect 8168 14900 8174 14912
rect 9125 14909 9137 14912
rect 9171 14909 9183 14943
rect 9306 14940 9312 14952
rect 9267 14912 9312 14940
rect 9125 14903 9183 14909
rect 9306 14900 9312 14912
rect 9364 14900 9370 14952
rect 10134 14940 10140 14952
rect 10095 14912 10140 14940
rect 10134 14900 10140 14912
rect 10192 14900 10198 14952
rect 10689 14943 10747 14949
rect 10689 14909 10701 14943
rect 10735 14940 10747 14943
rect 10778 14940 10784 14952
rect 10735 14912 10784 14940
rect 10735 14909 10747 14912
rect 10689 14903 10747 14909
rect 7984 14844 8064 14872
rect 7984 14832 7990 14844
rect 8662 14832 8668 14884
rect 8720 14872 8726 14884
rect 9493 14875 9551 14881
rect 9493 14872 9505 14875
rect 8720 14844 9505 14872
rect 8720 14832 8726 14844
rect 9493 14841 9505 14844
rect 9539 14841 9551 14875
rect 9950 14872 9956 14884
rect 9493 14835 9551 14841
rect 9600 14844 9956 14872
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 1670 14764 1676 14816
rect 1728 14804 1734 14816
rect 1765 14807 1823 14813
rect 1765 14804 1777 14807
rect 1728 14776 1777 14804
rect 1728 14764 1734 14776
rect 1765 14773 1777 14776
rect 1811 14773 1823 14807
rect 1765 14767 1823 14773
rect 2498 14764 2504 14816
rect 2556 14804 2562 14816
rect 2593 14807 2651 14813
rect 2593 14804 2605 14807
rect 2556 14776 2605 14804
rect 2556 14764 2562 14776
rect 2593 14773 2605 14776
rect 2639 14773 2651 14807
rect 3142 14804 3148 14816
rect 3103 14776 3148 14804
rect 2593 14767 2651 14773
rect 3142 14764 3148 14776
rect 3200 14764 3206 14816
rect 3602 14764 3608 14816
rect 3660 14804 3666 14816
rect 4338 14804 4344 14816
rect 3660 14776 4344 14804
rect 3660 14764 3666 14776
rect 4338 14764 4344 14776
rect 4396 14764 4402 14816
rect 6454 14764 6460 14816
rect 6512 14804 6518 14816
rect 8205 14807 8263 14813
rect 8205 14804 8217 14807
rect 6512 14776 8217 14804
rect 6512 14764 6518 14776
rect 8205 14773 8217 14776
rect 8251 14773 8263 14807
rect 8205 14767 8263 14773
rect 8386 14764 8392 14816
rect 8444 14804 8450 14816
rect 8481 14807 8539 14813
rect 8481 14804 8493 14807
rect 8444 14776 8493 14804
rect 8444 14764 8450 14776
rect 8481 14773 8493 14776
rect 8527 14773 8539 14807
rect 8481 14767 8539 14773
rect 8570 14764 8576 14816
rect 8628 14804 8634 14816
rect 9600 14804 9628 14844
rect 9950 14832 9956 14844
rect 10008 14872 10014 14884
rect 10704 14872 10732 14903
rect 10778 14900 10784 14912
rect 10836 14900 10842 14952
rect 11606 14940 11612 14952
rect 11567 14912 11612 14940
rect 11606 14900 11612 14912
rect 11664 14900 11670 14952
rect 11790 14940 11796 14952
rect 11751 14912 11796 14940
rect 11790 14900 11796 14912
rect 11848 14900 11854 14952
rect 12066 14900 12072 14952
rect 12124 14940 12130 14952
rect 12124 14912 12434 14940
rect 12124 14900 12130 14912
rect 10008 14844 10732 14872
rect 10008 14832 10014 14844
rect 11974 14832 11980 14884
rect 12032 14872 12038 14884
rect 12253 14875 12311 14881
rect 12253 14872 12265 14875
rect 12032 14844 12265 14872
rect 12032 14832 12038 14844
rect 12253 14841 12265 14844
rect 12299 14841 12311 14875
rect 12406 14872 12434 14912
rect 12618 14900 12624 14952
rect 12676 14940 12682 14952
rect 12897 14943 12955 14949
rect 12897 14940 12909 14943
rect 12676 14912 12909 14940
rect 12676 14900 12682 14912
rect 12897 14909 12909 14912
rect 12943 14909 12955 14943
rect 12897 14903 12955 14909
rect 12986 14900 12992 14952
rect 13044 14940 13050 14952
rect 13449 14943 13507 14949
rect 13449 14940 13461 14943
rect 13044 14912 13461 14940
rect 13044 14900 13050 14912
rect 13449 14909 13461 14912
rect 13495 14909 13507 14943
rect 13449 14903 13507 14909
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14940 13691 14943
rect 13722 14940 13728 14952
rect 13679 14912 13728 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 14108 14940 14136 14980
rect 14274 14968 14280 14980
rect 14332 14968 14338 15020
rect 15654 15008 15660 15020
rect 14568 14980 15660 15008
rect 14568 14940 14596 14980
rect 15654 14968 15660 14980
rect 15712 14968 15718 15020
rect 14108 14912 14596 14940
rect 14645 14943 14703 14949
rect 14645 14909 14657 14943
rect 14691 14909 14703 14943
rect 14645 14903 14703 14909
rect 12406 14844 12664 14872
rect 12253 14835 12311 14841
rect 8628 14776 9628 14804
rect 8628 14764 8634 14776
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 10410 14804 10416 14816
rect 9732 14776 10416 14804
rect 9732 14764 9738 14776
rect 10410 14764 10416 14776
rect 10468 14764 10474 14816
rect 10502 14764 10508 14816
rect 10560 14804 10566 14816
rect 12434 14804 12440 14816
rect 10560 14776 12440 14804
rect 10560 14764 10566 14776
rect 12434 14764 12440 14776
rect 12492 14764 12498 14816
rect 12636 14804 12664 14844
rect 14660 14804 14688 14903
rect 14826 14900 14832 14952
rect 14884 14940 14890 14952
rect 14921 14943 14979 14949
rect 14921 14940 14933 14943
rect 14884 14912 14933 14940
rect 14884 14900 14890 14912
rect 14921 14909 14933 14912
rect 14967 14909 14979 14943
rect 14921 14903 14979 14909
rect 12636 14776 14688 14804
rect 1104 14714 16008 14736
rect 1104 14662 2824 14714
rect 2876 14662 2888 14714
rect 2940 14662 2952 14714
rect 3004 14662 3016 14714
rect 3068 14662 3080 14714
rect 3132 14662 6572 14714
rect 6624 14662 6636 14714
rect 6688 14662 6700 14714
rect 6752 14662 6764 14714
rect 6816 14662 6828 14714
rect 6880 14662 10320 14714
rect 10372 14662 10384 14714
rect 10436 14662 10448 14714
rect 10500 14662 10512 14714
rect 10564 14662 10576 14714
rect 10628 14662 14068 14714
rect 14120 14662 14132 14714
rect 14184 14662 14196 14714
rect 14248 14662 14260 14714
rect 14312 14662 14324 14714
rect 14376 14662 16008 14714
rect 1104 14640 16008 14662
rect 1489 14603 1547 14609
rect 1489 14569 1501 14603
rect 1535 14600 1547 14603
rect 1578 14600 1584 14612
rect 1535 14572 1584 14600
rect 1535 14569 1547 14572
rect 1489 14563 1547 14569
rect 1578 14560 1584 14572
rect 1636 14560 1642 14612
rect 5074 14600 5080 14612
rect 5035 14572 5080 14600
rect 5074 14560 5080 14572
rect 5132 14560 5138 14612
rect 5718 14560 5724 14612
rect 5776 14600 5782 14612
rect 5905 14603 5963 14609
rect 5905 14600 5917 14603
rect 5776 14572 5917 14600
rect 5776 14560 5782 14572
rect 5905 14569 5917 14572
rect 5951 14569 5963 14603
rect 7006 14600 7012 14612
rect 6967 14572 7012 14600
rect 5905 14563 5963 14569
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 7282 14600 7288 14612
rect 7243 14572 7288 14600
rect 7282 14560 7288 14572
rect 7340 14560 7346 14612
rect 7650 14560 7656 14612
rect 7708 14600 7714 14612
rect 7708 14572 8248 14600
rect 7708 14560 7714 14572
rect 2590 14492 2596 14544
rect 2648 14532 2654 14544
rect 8113 14535 8171 14541
rect 8113 14532 8125 14535
rect 2648 14504 8125 14532
rect 2648 14492 2654 14504
rect 2961 14467 3019 14473
rect 2961 14433 2973 14467
rect 3007 14464 3019 14467
rect 3050 14464 3056 14476
rect 3007 14436 3056 14464
rect 3007 14433 3019 14436
rect 2961 14427 3019 14433
rect 3050 14424 3056 14436
rect 3108 14424 3114 14476
rect 3786 14424 3792 14476
rect 3844 14464 3850 14476
rect 5552 14473 5580 14504
rect 8113 14501 8125 14504
rect 8159 14501 8171 14535
rect 8220 14532 8248 14572
rect 8294 14560 8300 14612
rect 8352 14600 8358 14612
rect 8389 14603 8447 14609
rect 8389 14600 8401 14603
rect 8352 14572 8401 14600
rect 8352 14560 8358 14572
rect 8389 14569 8401 14572
rect 8435 14569 8447 14603
rect 8389 14563 8447 14569
rect 8754 14560 8760 14612
rect 8812 14600 8818 14612
rect 8812 14572 9168 14600
rect 8812 14560 8818 14572
rect 8941 14535 8999 14541
rect 8941 14532 8953 14535
rect 8220 14504 8953 14532
rect 8113 14495 8171 14501
rect 8941 14501 8953 14504
rect 8987 14501 8999 14535
rect 9140 14532 9168 14572
rect 9214 14560 9220 14612
rect 9272 14600 9278 14612
rect 9401 14603 9459 14609
rect 9401 14600 9413 14603
rect 9272 14572 9413 14600
rect 9272 14560 9278 14572
rect 9401 14569 9413 14572
rect 9447 14569 9459 14603
rect 9401 14563 9459 14569
rect 11422 14560 11428 14612
rect 11480 14600 11486 14612
rect 11701 14603 11759 14609
rect 11701 14600 11713 14603
rect 11480 14572 11713 14600
rect 11480 14560 11486 14572
rect 11701 14569 11713 14572
rect 11747 14569 11759 14603
rect 11701 14563 11759 14569
rect 12434 14560 12440 14612
rect 12492 14600 12498 14612
rect 12492 14572 13308 14600
rect 12492 14560 12498 14572
rect 9140 14504 9352 14532
rect 8941 14495 8999 14501
rect 4341 14467 4399 14473
rect 4341 14464 4353 14467
rect 3844 14436 4353 14464
rect 3844 14424 3850 14436
rect 4341 14433 4353 14436
rect 4387 14433 4399 14467
rect 4341 14427 4399 14433
rect 5537 14467 5595 14473
rect 5537 14433 5549 14467
rect 5583 14433 5595 14467
rect 5537 14427 5595 14433
rect 5721 14467 5779 14473
rect 5721 14433 5733 14467
rect 5767 14464 5779 14467
rect 5902 14464 5908 14476
rect 5767 14436 5908 14464
rect 5767 14433 5779 14436
rect 5721 14427 5779 14433
rect 5902 14424 5908 14436
rect 5960 14424 5966 14476
rect 6362 14424 6368 14476
rect 6420 14464 6426 14476
rect 6457 14467 6515 14473
rect 6457 14464 6469 14467
rect 6420 14436 6469 14464
rect 6420 14424 6426 14436
rect 6457 14433 6469 14436
rect 6503 14433 6515 14467
rect 7834 14464 7840 14476
rect 7795 14436 7840 14464
rect 6457 14427 6515 14433
rect 7834 14424 7840 14436
rect 7892 14424 7898 14476
rect 9030 14464 9036 14476
rect 8312 14436 9036 14464
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 2682 14396 2688 14408
rect 1719 14368 2688 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 3142 14396 3148 14408
rect 3103 14368 3148 14396
rect 3142 14356 3148 14368
rect 3200 14356 3206 14408
rect 4430 14356 4436 14408
rect 4488 14396 4494 14408
rect 4617 14399 4675 14405
rect 4617 14396 4629 14399
rect 4488 14368 4629 14396
rect 4488 14356 4494 14368
rect 4617 14365 4629 14368
rect 4663 14365 4675 14399
rect 4617 14359 4675 14365
rect 5350 14356 5356 14408
rect 5408 14396 5414 14408
rect 5445 14399 5503 14405
rect 5445 14396 5457 14399
rect 5408 14368 5457 14396
rect 5408 14356 5414 14368
rect 5445 14365 5457 14368
rect 5491 14365 5503 14399
rect 5445 14359 5503 14365
rect 5626 14356 5632 14408
rect 5684 14396 5690 14408
rect 6270 14396 6276 14408
rect 5684 14368 6276 14396
rect 5684 14356 5690 14368
rect 6270 14356 6276 14368
rect 6328 14356 6334 14408
rect 8312 14405 8340 14436
rect 9030 14424 9036 14436
rect 9088 14424 9094 14476
rect 9122 14424 9128 14476
rect 9180 14464 9186 14476
rect 9217 14467 9275 14473
rect 9217 14464 9229 14467
rect 9180 14436 9229 14464
rect 9180 14424 9186 14436
rect 9217 14433 9229 14436
rect 9263 14433 9275 14467
rect 9217 14427 9275 14433
rect 7653 14399 7711 14405
rect 7653 14365 7665 14399
rect 7699 14396 7711 14399
rect 8297 14399 8355 14405
rect 8297 14396 8309 14399
rect 7699 14368 8309 14396
rect 7699 14365 7711 14368
rect 7653 14359 7711 14365
rect 8297 14365 8309 14368
rect 8343 14365 8355 14399
rect 8297 14359 8355 14365
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14396 8631 14399
rect 8757 14399 8815 14405
rect 8757 14396 8769 14399
rect 8619 14368 8769 14396
rect 8619 14365 8631 14368
rect 8573 14359 8631 14365
rect 8757 14365 8769 14368
rect 8803 14396 8815 14399
rect 8846 14396 8852 14408
rect 8803 14368 8852 14396
rect 8803 14365 8815 14368
rect 8757 14359 8815 14365
rect 8846 14356 8852 14368
rect 8904 14356 8910 14408
rect 9125 14375 9183 14381
rect 9125 14341 9137 14375
rect 9171 14372 9183 14375
rect 9223 14372 9251 14427
rect 9171 14344 9251 14372
rect 9171 14341 9183 14344
rect 3053 14331 3111 14337
rect 3053 14297 3065 14331
rect 3099 14328 3111 14331
rect 4985 14331 5043 14337
rect 3099 14300 3832 14328
rect 3099 14297 3111 14300
rect 3053 14291 3111 14297
rect 3510 14260 3516 14272
rect 3471 14232 3516 14260
rect 3510 14220 3516 14232
rect 3568 14220 3574 14272
rect 3804 14269 3832 14300
rect 4985 14297 4997 14331
rect 5031 14328 5043 14331
rect 5718 14328 5724 14340
rect 5031 14300 5724 14328
rect 5031 14297 5043 14300
rect 4985 14291 5043 14297
rect 5718 14288 5724 14300
rect 5776 14288 5782 14340
rect 5994 14288 6000 14340
rect 6052 14328 6058 14340
rect 6178 14328 6184 14340
rect 6052 14300 6184 14328
rect 6052 14288 6058 14300
rect 6178 14288 6184 14300
rect 6236 14288 6242 14340
rect 6822 14328 6828 14340
rect 6380 14300 6828 14328
rect 3789 14263 3847 14269
rect 3789 14229 3801 14263
rect 3835 14229 3847 14263
rect 4154 14260 4160 14272
rect 4115 14232 4160 14260
rect 3789 14223 3847 14229
rect 4154 14220 4160 14232
rect 4212 14220 4218 14272
rect 4246 14220 4252 14272
rect 4304 14260 4310 14272
rect 6380 14269 6408 14300
rect 6822 14288 6828 14300
rect 6880 14288 6886 14340
rect 6914 14288 6920 14340
rect 6972 14328 6978 14340
rect 9125 14335 9183 14341
rect 9324 14328 9352 14504
rect 11514 14492 11520 14544
rect 11572 14532 11578 14544
rect 11974 14532 11980 14544
rect 11572 14504 11980 14532
rect 11572 14492 11578 14504
rect 11974 14492 11980 14504
rect 12032 14492 12038 14544
rect 13280 14532 13308 14572
rect 13354 14560 13360 14612
rect 13412 14600 13418 14612
rect 13541 14603 13599 14609
rect 13541 14600 13553 14603
rect 13412 14572 13553 14600
rect 13412 14560 13418 14572
rect 13541 14569 13553 14572
rect 13587 14569 13599 14603
rect 13541 14563 13599 14569
rect 14366 14532 14372 14544
rect 13280 14504 14372 14532
rect 14366 14492 14372 14504
rect 14424 14532 14430 14544
rect 14424 14504 14596 14532
rect 14424 14492 14430 14504
rect 9398 14424 9404 14476
rect 9456 14464 9462 14476
rect 9677 14467 9735 14473
rect 9677 14464 9689 14467
rect 9456 14436 9689 14464
rect 9456 14424 9462 14436
rect 9677 14433 9689 14436
rect 9723 14433 9735 14467
rect 9677 14427 9735 14433
rect 9950 14424 9956 14476
rect 10008 14464 10014 14476
rect 10229 14467 10287 14473
rect 10229 14464 10241 14467
rect 10008 14436 10241 14464
rect 10008 14424 10014 14436
rect 10229 14433 10241 14436
rect 10275 14433 10287 14467
rect 10229 14427 10287 14433
rect 11149 14467 11207 14473
rect 11149 14433 11161 14467
rect 11195 14464 11207 14467
rect 11238 14464 11244 14476
rect 11195 14436 11244 14464
rect 11195 14433 11207 14436
rect 11149 14427 11207 14433
rect 11238 14424 11244 14436
rect 11296 14464 11302 14476
rect 14568 14473 14596 14504
rect 13265 14467 13323 14473
rect 13265 14464 13277 14467
rect 11296 14436 12112 14464
rect 11296 14424 11302 14436
rect 12084 14396 12112 14436
rect 13096 14436 13277 14464
rect 12526 14396 12532 14408
rect 10612 14368 12020 14396
rect 12084 14368 12532 14396
rect 10612 14328 10640 14368
rect 6972 14300 7788 14328
rect 9324 14300 10640 14328
rect 6972 14288 6978 14300
rect 4801 14263 4859 14269
rect 4304 14232 4349 14260
rect 4304 14220 4310 14232
rect 4801 14229 4813 14263
rect 4847 14260 4859 14263
rect 6365 14263 6423 14269
rect 6365 14260 6377 14263
rect 4847 14232 6377 14260
rect 4847 14229 4859 14232
rect 4801 14223 4859 14229
rect 6365 14229 6377 14232
rect 6411 14229 6423 14263
rect 6365 14223 6423 14229
rect 6454 14220 6460 14272
rect 6512 14260 6518 14272
rect 6733 14263 6791 14269
rect 6733 14260 6745 14263
rect 6512 14232 6745 14260
rect 6512 14220 6518 14232
rect 6733 14229 6745 14232
rect 6779 14229 6791 14263
rect 6733 14223 6791 14229
rect 7193 14263 7251 14269
rect 7193 14229 7205 14263
rect 7239 14260 7251 14263
rect 7466 14260 7472 14272
rect 7239 14232 7472 14260
rect 7239 14229 7251 14232
rect 7193 14223 7251 14229
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 7760 14269 7788 14300
rect 10686 14288 10692 14340
rect 10744 14328 10750 14340
rect 11333 14331 11391 14337
rect 11333 14328 11345 14331
rect 10744 14300 11345 14328
rect 10744 14288 10750 14300
rect 11333 14297 11345 14300
rect 11379 14297 11391 14331
rect 11992 14328 12020 14368
rect 12526 14356 12532 14368
rect 12584 14356 12590 14408
rect 13096 14396 13124 14436
rect 13265 14433 13277 14436
rect 13311 14433 13323 14467
rect 13265 14427 13323 14433
rect 14553 14467 14611 14473
rect 14553 14433 14565 14467
rect 14599 14433 14611 14467
rect 14553 14427 14611 14433
rect 12820 14368 13124 14396
rect 13173 14399 13231 14405
rect 12820 14328 12848 14368
rect 13173 14365 13185 14399
rect 13219 14365 13231 14399
rect 13173 14359 13231 14365
rect 11992 14300 12848 14328
rect 11333 14291 11391 14297
rect 12894 14288 12900 14340
rect 12952 14337 12958 14340
rect 12952 14328 12964 14337
rect 12952 14300 12997 14328
rect 12952 14291 12964 14300
rect 12952 14288 12958 14291
rect 13078 14288 13084 14340
rect 13136 14328 13142 14340
rect 13188 14328 13216 14359
rect 13630 14356 13636 14408
rect 13688 14396 13694 14408
rect 13725 14399 13783 14405
rect 13725 14396 13737 14399
rect 13688 14368 13737 14396
rect 13688 14356 13694 14368
rect 13725 14365 13737 14368
rect 13771 14365 13783 14399
rect 13725 14359 13783 14365
rect 14829 14399 14887 14405
rect 14829 14365 14841 14399
rect 14875 14396 14887 14399
rect 15010 14396 15016 14408
rect 14875 14368 15016 14396
rect 14875 14365 14887 14368
rect 14829 14359 14887 14365
rect 15010 14356 15016 14368
rect 15068 14356 15074 14408
rect 15470 14356 15476 14408
rect 15528 14396 15534 14408
rect 15622 14399 15680 14405
rect 15622 14396 15634 14399
rect 15528 14368 15634 14396
rect 15528 14356 15534 14368
rect 15622 14365 15634 14368
rect 15668 14396 15680 14399
rect 16206 14396 16212 14408
rect 15668 14368 16212 14396
rect 15668 14365 15680 14368
rect 15622 14359 15680 14365
rect 16206 14356 16212 14368
rect 16264 14356 16270 14408
rect 13136 14300 13216 14328
rect 14369 14331 14427 14337
rect 13136 14288 13142 14300
rect 14369 14297 14381 14331
rect 14415 14328 14427 14331
rect 15746 14328 15752 14340
rect 14415 14300 15752 14328
rect 14415 14297 14427 14300
rect 14369 14291 14427 14297
rect 15746 14288 15752 14300
rect 15804 14328 15810 14340
rect 15930 14328 15936 14340
rect 15804 14300 15936 14328
rect 15804 14288 15810 14300
rect 15930 14288 15936 14300
rect 15988 14288 15994 14340
rect 7745 14263 7803 14269
rect 7745 14229 7757 14263
rect 7791 14260 7803 14263
rect 8938 14260 8944 14272
rect 7791 14232 8944 14260
rect 7791 14229 7803 14232
rect 7745 14223 7803 14229
rect 8938 14220 8944 14232
rect 8996 14220 9002 14272
rect 9766 14260 9772 14272
rect 9727 14232 9772 14260
rect 9766 14220 9772 14232
rect 9824 14220 9830 14272
rect 9950 14260 9956 14272
rect 9911 14232 9956 14260
rect 9950 14220 9956 14232
rect 10008 14260 10014 14272
rect 10413 14263 10471 14269
rect 10413 14260 10425 14263
rect 10008 14232 10425 14260
rect 10008 14220 10014 14232
rect 10413 14229 10425 14232
rect 10459 14229 10471 14263
rect 10413 14223 10471 14229
rect 10505 14263 10563 14269
rect 10505 14229 10517 14263
rect 10551 14260 10563 14263
rect 10778 14260 10784 14272
rect 10551 14232 10784 14260
rect 10551 14229 10563 14232
rect 10505 14223 10563 14229
rect 10778 14220 10784 14232
rect 10836 14220 10842 14272
rect 10873 14263 10931 14269
rect 10873 14229 10885 14263
rect 10919 14260 10931 14263
rect 11241 14263 11299 14269
rect 11241 14260 11253 14263
rect 10919 14232 11253 14260
rect 10919 14229 10931 14232
rect 10873 14223 10931 14229
rect 11241 14229 11253 14232
rect 11287 14229 11299 14263
rect 11790 14260 11796 14272
rect 11751 14232 11796 14260
rect 11241 14223 11299 14229
rect 11790 14220 11796 14232
rect 11848 14220 11854 14272
rect 11974 14220 11980 14272
rect 12032 14260 12038 14272
rect 13909 14263 13967 14269
rect 13909 14260 13921 14263
rect 12032 14232 13921 14260
rect 12032 14220 12038 14232
rect 13909 14229 13921 14232
rect 13955 14229 13967 14263
rect 14274 14260 14280 14272
rect 14235 14232 14280 14260
rect 13909 14223 13967 14229
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 15470 14220 15476 14272
rect 15528 14269 15534 14272
rect 15528 14263 15577 14269
rect 15528 14229 15531 14263
rect 15565 14229 15577 14263
rect 15528 14223 15577 14229
rect 15528 14220 15534 14223
rect 1104 14170 16008 14192
rect 1104 14118 4698 14170
rect 4750 14118 4762 14170
rect 4814 14118 4826 14170
rect 4878 14118 4890 14170
rect 4942 14118 4954 14170
rect 5006 14118 8446 14170
rect 8498 14118 8510 14170
rect 8562 14118 8574 14170
rect 8626 14118 8638 14170
rect 8690 14118 8702 14170
rect 8754 14118 12194 14170
rect 12246 14118 12258 14170
rect 12310 14118 12322 14170
rect 12374 14118 12386 14170
rect 12438 14118 12450 14170
rect 12502 14118 16008 14170
rect 1104 14096 16008 14118
rect 1026 14016 1032 14068
rect 1084 14056 1090 14068
rect 3605 14059 3663 14065
rect 3605 14056 3617 14059
rect 1084 14028 3617 14056
rect 1084 14016 1090 14028
rect 3605 14025 3617 14028
rect 3651 14025 3663 14059
rect 3605 14019 3663 14025
rect 4709 14059 4767 14065
rect 4709 14025 4721 14059
rect 4755 14025 4767 14059
rect 4709 14019 4767 14025
rect 2774 13948 2780 14000
rect 2832 13948 2838 14000
rect 2866 13948 2872 14000
rect 2924 13988 2930 14000
rect 3418 13988 3424 14000
rect 2924 13960 3424 13988
rect 2924 13948 2930 13960
rect 3418 13948 3424 13960
rect 3476 13948 3482 14000
rect 4246 13988 4252 14000
rect 4207 13960 4252 13988
rect 4246 13948 4252 13960
rect 4304 13948 4310 14000
rect 4724 13988 4752 14019
rect 5442 14016 5448 14068
rect 5500 14056 5506 14068
rect 7650 14056 7656 14068
rect 5500 14028 7656 14056
rect 5500 14016 5506 14028
rect 7650 14016 7656 14028
rect 7708 14056 7714 14068
rect 7745 14059 7803 14065
rect 7745 14056 7757 14059
rect 7708 14028 7757 14056
rect 7708 14016 7714 14028
rect 7745 14025 7757 14028
rect 7791 14025 7803 14059
rect 8018 14056 8024 14068
rect 7979 14028 8024 14056
rect 7745 14019 7803 14025
rect 8018 14016 8024 14028
rect 8076 14016 8082 14068
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 8481 14059 8539 14065
rect 8481 14056 8493 14059
rect 8260 14028 8493 14056
rect 8260 14016 8266 14028
rect 8481 14025 8493 14028
rect 8527 14025 8539 14059
rect 8481 14019 8539 14025
rect 8849 14059 8907 14065
rect 8849 14025 8861 14059
rect 8895 14025 8907 14059
rect 8849 14019 8907 14025
rect 5166 13988 5172 14000
rect 4724 13960 5172 13988
rect 5166 13948 5172 13960
rect 5224 13988 5230 14000
rect 6610 13991 6668 13997
rect 6610 13988 6622 13991
rect 5224 13960 6622 13988
rect 5224 13948 5230 13960
rect 6610 13957 6622 13960
rect 6656 13957 6668 13991
rect 6610 13951 6668 13957
rect 6822 13948 6828 14000
rect 6880 13988 6886 14000
rect 7558 13988 7564 14000
rect 6880 13960 7564 13988
rect 6880 13948 6886 13960
rect 7558 13948 7564 13960
rect 7616 13988 7622 14000
rect 8110 13988 8116 14000
rect 7616 13960 8116 13988
rect 7616 13948 7622 13960
rect 8110 13948 8116 13960
rect 8168 13988 8174 14000
rect 8389 13991 8447 13997
rect 8389 13988 8401 13991
rect 8168 13960 8401 13988
rect 8168 13948 8174 13960
rect 8389 13957 8401 13960
rect 8435 13957 8447 13991
rect 8864 13988 8892 14019
rect 9030 14016 9036 14068
rect 9088 14056 9094 14068
rect 9309 14059 9367 14065
rect 9309 14056 9321 14059
rect 9088 14028 9321 14056
rect 9088 14016 9094 14028
rect 9309 14025 9321 14028
rect 9355 14025 9367 14059
rect 9309 14019 9367 14025
rect 9677 14059 9735 14065
rect 9677 14025 9689 14059
rect 9723 14056 9735 14059
rect 10137 14059 10195 14065
rect 10137 14056 10149 14059
rect 9723 14028 10149 14056
rect 9723 14025 9735 14028
rect 9677 14019 9735 14025
rect 10137 14025 10149 14028
rect 10183 14025 10195 14059
rect 10137 14019 10195 14025
rect 10505 14059 10563 14065
rect 10505 14025 10517 14059
rect 10551 14056 10563 14059
rect 10686 14056 10692 14068
rect 10551 14028 10692 14056
rect 10551 14025 10563 14028
rect 10505 14019 10563 14025
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 13722 14056 13728 14068
rect 13683 14028 13728 14056
rect 13722 14016 13728 14028
rect 13780 14016 13786 14068
rect 10045 13991 10103 13997
rect 10045 13988 10057 13991
rect 8864 13960 10057 13988
rect 8389 13951 8447 13957
rect 10045 13957 10057 13960
rect 10091 13957 10103 13991
rect 10962 13988 10968 14000
rect 10923 13960 10968 13988
rect 10045 13951 10103 13957
rect 10962 13948 10968 13960
rect 11020 13948 11026 14000
rect 13078 13988 13084 14000
rect 11532 13960 13084 13988
rect 1670 13920 1676 13932
rect 1631 13892 1676 13920
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 2685 13923 2743 13929
rect 2685 13920 2697 13923
rect 2148 13892 2697 13920
rect 1394 13812 1400 13864
rect 1452 13852 1458 13864
rect 2148 13852 2176 13892
rect 2685 13889 2697 13892
rect 2731 13920 2743 13923
rect 2792 13920 2820 13948
rect 3145 13923 3203 13929
rect 3145 13920 3157 13923
rect 2731 13892 3157 13920
rect 2731 13889 2743 13892
rect 2685 13883 2743 13889
rect 3145 13889 3157 13892
rect 3191 13889 3203 13923
rect 3145 13883 3203 13889
rect 5810 13880 5816 13932
rect 5868 13929 5874 13932
rect 5868 13920 5880 13929
rect 5868 13892 5913 13920
rect 5868 13883 5880 13892
rect 5868 13880 5874 13883
rect 5994 13880 6000 13932
rect 6052 13920 6058 13932
rect 6089 13923 6147 13929
rect 6089 13920 6101 13923
rect 6052 13892 6101 13920
rect 6052 13880 6058 13892
rect 6089 13889 6101 13892
rect 6135 13920 6147 13923
rect 6365 13923 6423 13929
rect 6365 13920 6377 13923
rect 6135 13892 6377 13920
rect 6135 13889 6147 13892
rect 6089 13883 6147 13889
rect 6365 13889 6377 13892
rect 6411 13920 6423 13923
rect 6454 13920 6460 13932
rect 6411 13892 6460 13920
rect 6411 13889 6423 13892
rect 6365 13883 6423 13889
rect 6454 13880 6460 13892
rect 6512 13880 6518 13932
rect 8938 13880 8944 13932
rect 8996 13920 9002 13932
rect 9217 13923 9275 13929
rect 9217 13920 9229 13923
rect 8996 13892 9229 13920
rect 8996 13880 9002 13892
rect 9217 13889 9229 13892
rect 9263 13889 9275 13923
rect 9217 13883 9275 13889
rect 9950 13880 9956 13932
rect 10008 13920 10014 13932
rect 11532 13929 11560 13960
rect 13078 13948 13084 13960
rect 13136 13948 13142 14000
rect 13814 13988 13820 14000
rect 13775 13960 13820 13988
rect 13814 13948 13820 13960
rect 13872 13948 13878 14000
rect 15470 13988 15476 14000
rect 15431 13960 15476 13988
rect 15470 13948 15476 13960
rect 15528 13948 15534 14000
rect 11517 13923 11575 13929
rect 10008 13892 10824 13920
rect 10008 13880 10014 13892
rect 1452 13824 2176 13852
rect 1452 13812 1458 13824
rect 2222 13812 2228 13864
rect 2280 13852 2286 13864
rect 2777 13855 2835 13861
rect 2777 13852 2789 13855
rect 2280 13824 2789 13852
rect 2280 13812 2286 13824
rect 2777 13821 2789 13824
rect 2823 13852 2835 13855
rect 2866 13852 2872 13864
rect 2823 13824 2872 13852
rect 2823 13821 2835 13824
rect 2777 13815 2835 13821
rect 2866 13812 2872 13824
rect 2924 13812 2930 13864
rect 2961 13855 3019 13861
rect 2961 13821 2973 13855
rect 3007 13852 3019 13855
rect 3786 13852 3792 13864
rect 3007 13824 3792 13852
rect 3007 13821 3019 13824
rect 2961 13815 3019 13821
rect 3786 13812 3792 13824
rect 3844 13812 3850 13864
rect 4154 13812 4160 13864
rect 4212 13852 4218 13864
rect 4341 13855 4399 13861
rect 4341 13852 4353 13855
rect 4212 13824 4353 13852
rect 4212 13812 4218 13824
rect 4341 13821 4353 13824
rect 4387 13821 4399 13855
rect 4341 13815 4399 13821
rect 8297 13855 8355 13861
rect 8297 13821 8309 13855
rect 8343 13821 8355 13855
rect 8297 13815 8355 13821
rect 9125 13855 9183 13861
rect 9125 13821 9137 13855
rect 9171 13821 9183 13855
rect 9125 13815 9183 13821
rect 9861 13855 9919 13861
rect 9861 13821 9873 13855
rect 9907 13821 9919 13855
rect 9861 13815 9919 13821
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13821 10747 13855
rect 10796 13852 10824 13892
rect 11517 13889 11529 13923
rect 11563 13889 11575 13923
rect 11517 13883 11575 13889
rect 11784 13923 11842 13929
rect 11784 13889 11796 13923
rect 11830 13920 11842 13923
rect 12802 13920 12808 13932
rect 11830 13892 12808 13920
rect 11830 13889 11842 13892
rect 11784 13883 11842 13889
rect 12802 13880 12808 13892
rect 12860 13920 12866 13932
rect 13354 13920 13360 13932
rect 12860 13892 13216 13920
rect 13315 13892 13360 13920
rect 12860 13880 12866 13892
rect 13188 13864 13216 13892
rect 13354 13880 13360 13892
rect 13412 13880 13418 13932
rect 10873 13855 10931 13861
rect 10873 13852 10885 13855
rect 10796 13824 10885 13852
rect 10689 13815 10747 13821
rect 10873 13821 10885 13824
rect 10919 13852 10931 13855
rect 13170 13852 13176 13864
rect 10919 13824 11008 13852
rect 13131 13824 13176 13852
rect 10919 13821 10931 13824
rect 10873 13815 10931 13821
rect 1486 13784 1492 13796
rect 1447 13756 1492 13784
rect 1486 13744 1492 13756
rect 1544 13744 1550 13796
rect 8312 13784 8340 13815
rect 9140 13784 9168 13815
rect 8312 13756 9168 13784
rect 9876 13784 9904 13815
rect 9950 13784 9956 13796
rect 9876 13756 9956 13784
rect 2314 13716 2320 13728
rect 2275 13688 2320 13716
rect 2314 13676 2320 13688
rect 2372 13676 2378 13728
rect 4522 13716 4528 13728
rect 4483 13688 4528 13716
rect 4522 13676 4528 13688
rect 4580 13676 4586 13728
rect 9140 13716 9168 13756
rect 9950 13744 9956 13756
rect 10008 13744 10014 13796
rect 9858 13716 9864 13728
rect 9140 13688 9864 13716
rect 9858 13676 9864 13688
rect 9916 13716 9922 13728
rect 10704 13716 10732 13815
rect 10980 13784 11008 13824
rect 13170 13812 13176 13824
rect 13228 13812 13234 13864
rect 13265 13855 13323 13861
rect 13265 13821 13277 13855
rect 13311 13852 13323 13855
rect 13722 13852 13728 13864
rect 13311 13824 13728 13852
rect 13311 13821 13323 13824
rect 13265 13815 13323 13821
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 15654 13852 15660 13864
rect 15615 13824 15660 13852
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 11422 13784 11428 13796
rect 10980 13756 11428 13784
rect 11422 13744 11428 13756
rect 11480 13744 11486 13796
rect 14642 13784 14648 13796
rect 12820 13756 14648 13784
rect 11330 13716 11336 13728
rect 9916 13688 10732 13716
rect 11291 13688 11336 13716
rect 9916 13676 9922 13688
rect 11330 13676 11336 13688
rect 11388 13676 11394 13728
rect 11790 13676 11796 13728
rect 11848 13716 11854 13728
rect 12820 13716 12848 13756
rect 14642 13744 14648 13756
rect 14700 13744 14706 13796
rect 11848 13688 12848 13716
rect 11848 13676 11854 13688
rect 12894 13676 12900 13728
rect 12952 13716 12958 13728
rect 12952 13688 12997 13716
rect 12952 13676 12958 13688
rect 14366 13676 14372 13728
rect 14424 13716 14430 13728
rect 15470 13716 15476 13728
rect 14424 13688 15476 13716
rect 14424 13676 14430 13688
rect 15470 13676 15476 13688
rect 15528 13676 15534 13728
rect 1104 13626 16008 13648
rect 1104 13574 2824 13626
rect 2876 13574 2888 13626
rect 2940 13574 2952 13626
rect 3004 13574 3016 13626
rect 3068 13574 3080 13626
rect 3132 13574 6572 13626
rect 6624 13574 6636 13626
rect 6688 13574 6700 13626
rect 6752 13574 6764 13626
rect 6816 13574 6828 13626
rect 6880 13574 10320 13626
rect 10372 13574 10384 13626
rect 10436 13574 10448 13626
rect 10500 13574 10512 13626
rect 10564 13574 10576 13626
rect 10628 13574 14068 13626
rect 14120 13574 14132 13626
rect 14184 13574 14196 13626
rect 14248 13574 14260 13626
rect 14312 13574 14324 13626
rect 14376 13574 16008 13626
rect 1104 13552 16008 13574
rect 3142 13472 3148 13524
rect 3200 13512 3206 13524
rect 4062 13512 4068 13524
rect 3200 13484 4068 13512
rect 3200 13472 3206 13484
rect 4062 13472 4068 13484
rect 4120 13512 4126 13524
rect 5261 13515 5319 13521
rect 5261 13512 5273 13515
rect 4120 13484 5273 13512
rect 4120 13472 4126 13484
rect 5261 13481 5273 13484
rect 5307 13481 5319 13515
rect 5261 13475 5319 13481
rect 5629 13515 5687 13521
rect 5629 13481 5641 13515
rect 5675 13512 5687 13515
rect 5902 13512 5908 13524
rect 5675 13484 5908 13512
rect 5675 13481 5687 13484
rect 5629 13475 5687 13481
rect 5902 13472 5908 13484
rect 5960 13472 5966 13524
rect 6270 13472 6276 13524
rect 6328 13512 6334 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 6328 13484 8953 13512
rect 6328 13472 6334 13484
rect 8941 13481 8953 13484
rect 8987 13481 8999 13515
rect 9122 13512 9128 13524
rect 9083 13484 9128 13512
rect 8941 13475 8999 13481
rect 1765 13447 1823 13453
rect 1765 13413 1777 13447
rect 1811 13413 1823 13447
rect 2869 13447 2927 13453
rect 2869 13444 2881 13447
rect 1765 13407 1823 13413
rect 1964 13416 2881 13444
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 1780 13308 1808 13407
rect 1964 13317 1992 13416
rect 2869 13413 2881 13416
rect 2915 13413 2927 13447
rect 8956 13444 8984 13475
rect 9122 13472 9128 13484
rect 9180 13472 9186 13524
rect 9766 13512 9772 13524
rect 9727 13484 9772 13512
rect 9766 13472 9772 13484
rect 9824 13472 9830 13524
rect 11241 13515 11299 13521
rect 11241 13481 11253 13515
rect 11287 13512 11299 13515
rect 11606 13512 11612 13524
rect 11287 13484 11612 13512
rect 11287 13481 11299 13484
rect 11241 13475 11299 13481
rect 11606 13472 11612 13484
rect 11664 13472 11670 13524
rect 11974 13472 11980 13524
rect 12032 13512 12038 13524
rect 12802 13512 12808 13524
rect 12032 13484 12808 13512
rect 12032 13472 12038 13484
rect 12802 13472 12808 13484
rect 12860 13472 12866 13524
rect 12897 13515 12955 13521
rect 12897 13481 12909 13515
rect 12943 13512 12955 13515
rect 13078 13512 13084 13524
rect 12943 13484 13084 13512
rect 12943 13481 12955 13484
rect 12897 13475 12955 13481
rect 9030 13444 9036 13456
rect 8956 13416 9036 13444
rect 2869 13407 2927 13413
rect 9030 13404 9036 13416
rect 9088 13404 9094 13456
rect 9585 13447 9643 13453
rect 9585 13413 9597 13447
rect 9631 13444 9643 13447
rect 9674 13444 9680 13456
rect 9631 13416 9680 13444
rect 9631 13413 9643 13416
rect 9585 13407 9643 13413
rect 9674 13404 9680 13416
rect 9732 13404 9738 13456
rect 2225 13379 2283 13385
rect 2225 13345 2237 13379
rect 2271 13376 2283 13379
rect 3142 13376 3148 13388
rect 2271 13348 3148 13376
rect 2271 13345 2283 13348
rect 2225 13339 2283 13345
rect 3142 13336 3148 13348
rect 3200 13336 3206 13388
rect 3418 13376 3424 13388
rect 3379 13348 3424 13376
rect 3418 13336 3424 13348
rect 3476 13336 3482 13388
rect 9784 13376 9812 13472
rect 11146 13404 11152 13456
rect 11204 13444 11210 13456
rect 11333 13447 11391 13453
rect 11333 13444 11345 13447
rect 11204 13416 11345 13444
rect 11204 13404 11210 13416
rect 11333 13413 11345 13416
rect 11379 13413 11391 13447
rect 11333 13407 11391 13413
rect 9861 13379 9919 13385
rect 9861 13376 9873 13379
rect 9784 13348 9873 13376
rect 9861 13345 9873 13348
rect 9907 13345 9919 13379
rect 9861 13339 9919 13345
rect 12713 13379 12771 13385
rect 12713 13345 12725 13379
rect 12759 13376 12771 13379
rect 12912 13376 12940 13475
rect 13078 13472 13084 13484
rect 13136 13472 13142 13524
rect 13173 13515 13231 13521
rect 13173 13481 13185 13515
rect 13219 13512 13231 13515
rect 13354 13512 13360 13524
rect 13219 13484 13360 13512
rect 13219 13481 13231 13484
rect 13173 13475 13231 13481
rect 13354 13472 13360 13484
rect 13412 13472 13418 13524
rect 13722 13472 13728 13524
rect 13780 13512 13786 13524
rect 14921 13515 14979 13521
rect 14921 13512 14933 13515
rect 13780 13484 14933 13512
rect 13780 13472 13786 13484
rect 14921 13481 14933 13484
rect 14967 13481 14979 13515
rect 14921 13475 14979 13481
rect 13740 13416 15516 13444
rect 13740 13385 13768 13416
rect 12759 13348 12940 13376
rect 13725 13379 13783 13385
rect 12759 13345 12771 13348
rect 12713 13339 12771 13345
rect 13725 13345 13737 13379
rect 13771 13345 13783 13379
rect 14642 13376 14648 13388
rect 14603 13348 14648 13376
rect 13725 13339 13783 13345
rect 1719 13280 1808 13308
rect 1949 13311 2007 13317
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 1949 13277 1961 13311
rect 1995 13277 2007 13311
rect 1949 13271 2007 13277
rect 2314 13268 2320 13320
rect 2372 13308 2378 13320
rect 2409 13311 2467 13317
rect 2409 13308 2421 13311
rect 2372 13280 2421 13308
rect 2372 13268 2378 13280
rect 2409 13277 2421 13280
rect 2455 13277 2467 13311
rect 2409 13271 2467 13277
rect 3237 13311 3295 13317
rect 3237 13277 3249 13311
rect 3283 13308 3295 13311
rect 3510 13308 3516 13320
rect 3283 13280 3516 13308
rect 3283 13277 3295 13280
rect 3237 13271 3295 13277
rect 3510 13268 3516 13280
rect 3568 13268 3574 13320
rect 3881 13311 3939 13317
rect 3881 13277 3893 13311
rect 3927 13308 3939 13311
rect 4522 13308 4528 13320
rect 3927 13280 4528 13308
rect 3927 13277 3939 13280
rect 3881 13271 3939 13277
rect 4522 13268 4528 13280
rect 4580 13308 4586 13320
rect 5445 13311 5503 13317
rect 5445 13308 5457 13311
rect 4580 13280 5457 13308
rect 4580 13268 4586 13280
rect 5445 13277 5457 13280
rect 5491 13308 5503 13311
rect 5994 13308 6000 13320
rect 5491 13280 6000 13308
rect 5491 13277 5503 13280
rect 5445 13271 5503 13277
rect 5994 13268 6000 13280
rect 6052 13308 6058 13320
rect 7650 13317 7656 13320
rect 7009 13311 7067 13317
rect 7009 13308 7021 13311
rect 6052 13280 7021 13308
rect 6052 13268 6058 13280
rect 6656 13252 6684 13280
rect 7009 13277 7021 13280
rect 7055 13308 7067 13311
rect 7193 13311 7251 13317
rect 7193 13308 7205 13311
rect 7055 13280 7205 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 7193 13277 7205 13280
rect 7239 13308 7251 13311
rect 7377 13311 7435 13317
rect 7377 13308 7389 13311
rect 7239 13280 7389 13308
rect 7239 13277 7251 13280
rect 7193 13271 7251 13277
rect 7377 13277 7389 13280
rect 7423 13277 7435 13311
rect 7644 13308 7656 13317
rect 7611 13280 7656 13308
rect 7377 13271 7435 13277
rect 7644 13271 7656 13280
rect 7650 13268 7656 13271
rect 7708 13268 7714 13320
rect 10134 13317 10140 13320
rect 10128 13308 10140 13317
rect 10095 13280 10140 13308
rect 10128 13271 10140 13280
rect 10134 13268 10140 13271
rect 10192 13268 10198 13320
rect 11606 13268 11612 13320
rect 11664 13308 11670 13320
rect 13740 13308 13768 13339
rect 14642 13336 14648 13348
rect 14700 13336 14706 13388
rect 15488 13385 15516 13416
rect 15473 13379 15531 13385
rect 15473 13345 15485 13379
rect 15519 13345 15531 13379
rect 15473 13339 15531 13345
rect 14550 13308 14556 13320
rect 11664 13280 13768 13308
rect 14511 13280 14556 13308
rect 11664 13268 11670 13280
rect 14550 13268 14556 13280
rect 14608 13268 14614 13320
rect 15381 13311 15439 13317
rect 15381 13277 15393 13311
rect 15427 13308 15439 13311
rect 15746 13308 15752 13320
rect 15427 13280 15752 13308
rect 15427 13277 15439 13280
rect 15381 13271 15439 13277
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 3329 13243 3387 13249
rect 3329 13240 3341 13243
rect 2792 13212 3341 13240
rect 1486 13172 1492 13184
rect 1447 13144 1492 13172
rect 1486 13132 1492 13144
rect 1544 13132 1550 13184
rect 2314 13172 2320 13184
rect 2275 13144 2320 13172
rect 2314 13132 2320 13144
rect 2372 13132 2378 13184
rect 2792 13181 2820 13212
rect 3329 13209 3341 13212
rect 3375 13209 3387 13243
rect 3329 13203 3387 13209
rect 3786 13200 3792 13252
rect 3844 13240 3850 13252
rect 4126 13243 4184 13249
rect 4126 13240 4138 13243
rect 3844 13212 4138 13240
rect 3844 13200 3850 13212
rect 4126 13209 4138 13212
rect 4172 13209 4184 13243
rect 4126 13203 4184 13209
rect 6638 13200 6644 13252
rect 6696 13200 6702 13252
rect 6742 13243 6800 13249
rect 6742 13209 6754 13243
rect 6788 13209 6800 13243
rect 12468 13243 12526 13249
rect 12468 13240 12480 13243
rect 6742 13203 6800 13209
rect 8772 13212 12480 13240
rect 2777 13175 2835 13181
rect 2777 13141 2789 13175
rect 2823 13141 2835 13175
rect 2777 13135 2835 13141
rect 6362 13132 6368 13184
rect 6420 13172 6426 13184
rect 6748 13172 6776 13203
rect 8772 13181 8800 13212
rect 12468 13209 12480 13212
rect 12514 13240 12526 13243
rect 12618 13240 12624 13252
rect 12514 13212 12624 13240
rect 12514 13209 12526 13212
rect 12468 13203 12526 13209
rect 12618 13200 12624 13212
rect 12676 13200 12682 13252
rect 12802 13200 12808 13252
rect 12860 13240 12866 13252
rect 13354 13240 13360 13252
rect 12860 13212 13360 13240
rect 12860 13200 12866 13212
rect 13354 13200 13360 13212
rect 13412 13240 13418 13252
rect 13633 13243 13691 13249
rect 13633 13240 13645 13243
rect 13412 13212 13645 13240
rect 13412 13200 13418 13212
rect 13633 13209 13645 13212
rect 13679 13209 13691 13243
rect 13633 13203 13691 13209
rect 14366 13200 14372 13252
rect 14424 13240 14430 13252
rect 15102 13240 15108 13252
rect 14424 13212 15108 13240
rect 14424 13200 14430 13212
rect 15102 13200 15108 13212
rect 15160 13200 15166 13252
rect 15289 13243 15347 13249
rect 15289 13209 15301 13243
rect 15335 13240 15347 13243
rect 15470 13240 15476 13252
rect 15335 13212 15476 13240
rect 15335 13209 15347 13212
rect 15289 13203 15347 13209
rect 15470 13200 15476 13212
rect 15528 13200 15534 13252
rect 6420 13144 6776 13172
rect 8757 13175 8815 13181
rect 6420 13132 6426 13144
rect 8757 13141 8769 13175
rect 8803 13141 8815 13175
rect 8757 13135 8815 13141
rect 9401 13175 9459 13181
rect 9401 13141 9413 13175
rect 9447 13172 9459 13175
rect 10042 13172 10048 13184
rect 9447 13144 10048 13172
rect 9447 13141 9459 13144
rect 9401 13135 9459 13141
rect 10042 13132 10048 13144
rect 10100 13132 10106 13184
rect 10778 13132 10784 13184
rect 10836 13172 10842 13184
rect 10962 13172 10968 13184
rect 10836 13144 10968 13172
rect 10836 13132 10842 13144
rect 10962 13132 10968 13144
rect 11020 13132 11026 13184
rect 12066 13132 12072 13184
rect 12124 13172 12130 13184
rect 13541 13175 13599 13181
rect 13541 13172 13553 13175
rect 12124 13144 13553 13172
rect 12124 13132 12130 13144
rect 13541 13141 13553 13144
rect 13587 13141 13599 13175
rect 14090 13172 14096 13184
rect 14051 13144 14096 13172
rect 13541 13135 13599 13141
rect 14090 13132 14096 13144
rect 14148 13132 14154 13184
rect 14182 13132 14188 13184
rect 14240 13172 14246 13184
rect 14461 13175 14519 13181
rect 14461 13172 14473 13175
rect 14240 13144 14473 13172
rect 14240 13132 14246 13144
rect 14461 13141 14473 13144
rect 14507 13141 14519 13175
rect 14461 13135 14519 13141
rect 1104 13082 16008 13104
rect 1104 13030 4698 13082
rect 4750 13030 4762 13082
rect 4814 13030 4826 13082
rect 4878 13030 4890 13082
rect 4942 13030 4954 13082
rect 5006 13030 8446 13082
rect 8498 13030 8510 13082
rect 8562 13030 8574 13082
rect 8626 13030 8638 13082
rect 8690 13030 8702 13082
rect 8754 13030 12194 13082
rect 12246 13030 12258 13082
rect 12310 13030 12322 13082
rect 12374 13030 12386 13082
rect 12438 13030 12450 13082
rect 12502 13030 16008 13082
rect 1104 13008 16008 13030
rect 2314 12928 2320 12980
rect 2372 12968 2378 12980
rect 2409 12971 2467 12977
rect 2409 12968 2421 12971
rect 2372 12940 2421 12968
rect 2372 12928 2378 12940
rect 2409 12937 2421 12940
rect 2455 12937 2467 12971
rect 2409 12931 2467 12937
rect 3329 12971 3387 12977
rect 3329 12937 3341 12971
rect 3375 12937 3387 12971
rect 3329 12931 3387 12937
rect 3344 12900 3372 12931
rect 3418 12928 3424 12980
rect 3476 12968 3482 12980
rect 6181 12971 6239 12977
rect 6181 12968 6193 12971
rect 3476 12940 6193 12968
rect 3476 12928 3482 12940
rect 6181 12937 6193 12940
rect 6227 12937 6239 12971
rect 6181 12931 6239 12937
rect 3786 12900 3792 12912
rect 3344 12872 3792 12900
rect 2317 12835 2375 12841
rect 2317 12801 2329 12835
rect 2363 12832 2375 12835
rect 2498 12832 2504 12844
rect 2363 12804 2504 12832
rect 2363 12801 2375 12804
rect 2317 12795 2375 12801
rect 2498 12792 2504 12804
rect 2556 12832 2562 12844
rect 2777 12835 2835 12841
rect 2777 12832 2789 12835
rect 2556 12804 2789 12832
rect 2556 12792 2562 12804
rect 2777 12801 2789 12804
rect 2823 12801 2835 12835
rect 2777 12795 2835 12801
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12832 2927 12835
rect 3142 12832 3148 12844
rect 2915 12804 3148 12832
rect 2915 12801 2927 12804
rect 2869 12795 2927 12801
rect 2792 12764 2820 12795
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 3053 12767 3111 12773
rect 2792 12736 2912 12764
rect 2884 12696 2912 12736
rect 3053 12733 3065 12767
rect 3099 12764 3111 12767
rect 3344 12764 3372 12872
rect 3786 12860 3792 12872
rect 3844 12860 3850 12912
rect 4062 12860 4068 12912
rect 4120 12900 4126 12912
rect 5046 12903 5104 12909
rect 5046 12900 5058 12903
rect 4120 12872 5058 12900
rect 4120 12860 4126 12872
rect 5046 12869 5058 12872
rect 5092 12869 5104 12903
rect 5046 12863 5104 12869
rect 4154 12792 4160 12844
rect 4212 12832 4218 12844
rect 4442 12835 4500 12841
rect 4442 12832 4454 12835
rect 4212 12804 4454 12832
rect 4212 12792 4218 12804
rect 4442 12801 4454 12804
rect 4488 12801 4500 12835
rect 4442 12795 4500 12801
rect 3099 12736 3372 12764
rect 4709 12767 4767 12773
rect 3099 12733 3111 12736
rect 3053 12727 3111 12733
rect 4709 12733 4721 12767
rect 4755 12764 4767 12767
rect 4798 12764 4804 12776
rect 4755 12736 4804 12764
rect 4755 12733 4767 12736
rect 4709 12727 4767 12733
rect 4798 12724 4804 12736
rect 4856 12724 4862 12776
rect 6196 12764 6224 12931
rect 6638 12928 6644 12980
rect 6696 12968 6702 12980
rect 7193 12971 7251 12977
rect 7193 12968 7205 12971
rect 6696 12940 7205 12968
rect 6696 12928 6702 12940
rect 7193 12937 7205 12940
rect 7239 12937 7251 12971
rect 7193 12931 7251 12937
rect 8757 12971 8815 12977
rect 8757 12937 8769 12971
rect 8803 12937 8815 12971
rect 8757 12931 8815 12937
rect 7208 12832 7236 12931
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 7208 12804 7389 12832
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7633 12835 7691 12841
rect 7633 12832 7645 12835
rect 7377 12795 7435 12801
rect 7484 12804 7645 12832
rect 7484 12764 7512 12804
rect 7633 12801 7645 12804
rect 7679 12801 7691 12835
rect 8772 12832 8800 12931
rect 9122 12928 9128 12980
rect 9180 12968 9186 12980
rect 10042 12968 10048 12980
rect 9180 12940 10048 12968
rect 9180 12928 9186 12940
rect 10042 12928 10048 12940
rect 10100 12968 10106 12980
rect 10505 12971 10563 12977
rect 10505 12968 10517 12971
rect 10100 12940 10517 12968
rect 10100 12928 10106 12940
rect 10505 12937 10517 12940
rect 10551 12937 10563 12971
rect 10505 12931 10563 12937
rect 10594 12928 10600 12980
rect 10652 12968 10658 12980
rect 10689 12971 10747 12977
rect 10689 12968 10701 12971
rect 10652 12940 10701 12968
rect 10652 12928 10658 12940
rect 10689 12937 10701 12940
rect 10735 12937 10747 12971
rect 10689 12931 10747 12937
rect 10778 12928 10784 12980
rect 10836 12968 10842 12980
rect 10873 12971 10931 12977
rect 10873 12968 10885 12971
rect 10836 12940 10885 12968
rect 10836 12928 10842 12940
rect 10873 12937 10885 12940
rect 10919 12937 10931 12971
rect 10873 12931 10931 12937
rect 11146 12928 11152 12980
rect 11204 12968 11210 12980
rect 12342 12968 12348 12980
rect 11204 12940 12348 12968
rect 11204 12928 11210 12940
rect 12342 12928 12348 12940
rect 12400 12928 12406 12980
rect 12710 12928 12716 12980
rect 12768 12968 12774 12980
rect 12989 12971 13047 12977
rect 12989 12968 13001 12971
rect 12768 12940 13001 12968
rect 12768 12928 12774 12940
rect 12989 12937 13001 12940
rect 13035 12937 13047 12971
rect 13262 12968 13268 12980
rect 13223 12940 13268 12968
rect 12989 12931 13047 12937
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 13725 12971 13783 12977
rect 13725 12937 13737 12971
rect 13771 12968 13783 12971
rect 14277 12971 14335 12977
rect 14277 12968 14289 12971
rect 13771 12940 14289 12968
rect 13771 12937 13783 12940
rect 13725 12931 13783 12937
rect 14277 12937 14289 12940
rect 14323 12937 14335 12971
rect 14734 12968 14740 12980
rect 14695 12940 14740 12968
rect 14277 12931 14335 12937
rect 14734 12928 14740 12940
rect 14792 12968 14798 12980
rect 15102 12968 15108 12980
rect 14792 12940 15108 12968
rect 14792 12928 14798 12940
rect 15102 12928 15108 12940
rect 15160 12928 15166 12980
rect 15381 12971 15439 12977
rect 15381 12937 15393 12971
rect 15427 12968 15439 12971
rect 16114 12968 16120 12980
rect 15427 12940 16120 12968
rect 15427 12937 15439 12940
rect 15381 12931 15439 12937
rect 16114 12928 16120 12940
rect 16172 12928 16178 12980
rect 8941 12903 8999 12909
rect 8941 12869 8953 12903
rect 8987 12900 8999 12903
rect 9766 12900 9772 12912
rect 8987 12872 9772 12900
rect 8987 12869 8999 12872
rect 8941 12863 8999 12869
rect 9766 12860 9772 12872
rect 9824 12900 9830 12912
rect 10962 12900 10968 12912
rect 9824 12872 10968 12900
rect 9824 12860 9830 12872
rect 9306 12832 9312 12844
rect 8772 12804 9312 12832
rect 7633 12795 7691 12801
rect 9306 12792 9312 12804
rect 9364 12832 9370 12844
rect 10428 12841 10456 12872
rect 10962 12860 10968 12872
rect 11020 12900 11026 12912
rect 11241 12903 11299 12909
rect 11241 12900 11253 12903
rect 11020 12872 11253 12900
rect 11020 12860 11026 12872
rect 11241 12869 11253 12872
rect 11287 12869 11299 12903
rect 13078 12900 13084 12912
rect 11241 12863 11299 12869
rect 11532 12872 13084 12900
rect 10146 12835 10204 12841
rect 10146 12832 10158 12835
rect 9364 12804 10158 12832
rect 9364 12792 9370 12804
rect 10146 12801 10158 12804
rect 10192 12801 10204 12835
rect 10146 12795 10204 12801
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12801 10471 12835
rect 11256 12832 11284 12863
rect 11532 12841 11560 12872
rect 13078 12860 13084 12872
rect 13136 12860 13142 12912
rect 14366 12860 14372 12912
rect 14424 12900 14430 12912
rect 14645 12903 14703 12909
rect 14645 12900 14657 12903
rect 14424 12872 14657 12900
rect 14424 12860 14430 12872
rect 14645 12869 14657 12872
rect 14691 12869 14703 12903
rect 14645 12863 14703 12869
rect 11517 12835 11575 12841
rect 11517 12832 11529 12835
rect 11256 12804 11529 12832
rect 10413 12795 10471 12801
rect 11517 12801 11529 12804
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 11606 12792 11612 12844
rect 11664 12832 11670 12844
rect 11773 12835 11831 12841
rect 11773 12832 11785 12835
rect 11664 12804 11785 12832
rect 11664 12792 11670 12804
rect 11773 12801 11785 12804
rect 11819 12801 11831 12835
rect 13814 12832 13820 12844
rect 13775 12804 13820 12832
rect 11773 12795 11831 12801
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 14734 12792 14740 12844
rect 14792 12832 14798 12844
rect 14918 12832 14924 12844
rect 14792 12804 14924 12832
rect 14792 12792 14798 12804
rect 14918 12792 14924 12804
rect 14976 12792 14982 12844
rect 15194 12832 15200 12844
rect 15155 12804 15200 12832
rect 15194 12792 15200 12804
rect 15252 12792 15258 12844
rect 15473 12835 15531 12841
rect 15473 12801 15485 12835
rect 15519 12832 15531 12835
rect 15562 12832 15568 12844
rect 15519 12804 15568 12832
rect 15519 12801 15531 12804
rect 15473 12795 15531 12801
rect 15562 12792 15568 12804
rect 15620 12792 15626 12844
rect 6196 12736 7512 12764
rect 11149 12767 11207 12773
rect 11149 12733 11161 12767
rect 11195 12764 11207 12767
rect 11422 12764 11428 12776
rect 11195 12736 11428 12764
rect 11195 12733 11207 12736
rect 11149 12727 11207 12733
rect 11422 12724 11428 12736
rect 11480 12724 11486 12776
rect 12894 12724 12900 12776
rect 12952 12764 12958 12776
rect 13541 12767 13599 12773
rect 13541 12764 13553 12767
rect 12952 12736 13553 12764
rect 12952 12724 12958 12736
rect 13541 12733 13553 12736
rect 13587 12733 13599 12767
rect 13541 12727 13599 12733
rect 14829 12767 14887 12773
rect 14829 12733 14841 12767
rect 14875 12764 14887 12767
rect 14875 12736 14964 12764
rect 14875 12733 14887 12736
rect 14829 12727 14887 12733
rect 14936 12708 14964 12736
rect 3418 12696 3424 12708
rect 2884 12668 3424 12696
rect 3418 12656 3424 12668
rect 3476 12656 3482 12708
rect 8846 12656 8852 12708
rect 8904 12696 8910 12708
rect 9306 12696 9312 12708
rect 8904 12668 9312 12696
rect 8904 12656 8910 12668
rect 9306 12656 9312 12668
rect 9364 12656 9370 12708
rect 10778 12656 10784 12708
rect 10836 12656 10842 12708
rect 14182 12696 14188 12708
rect 14143 12668 14188 12696
rect 14182 12656 14188 12668
rect 14240 12656 14246 12708
rect 14918 12656 14924 12708
rect 14976 12656 14982 12708
rect 15654 12696 15660 12708
rect 15615 12668 15660 12696
rect 15654 12656 15660 12668
rect 15712 12656 15718 12708
rect 9030 12628 9036 12640
rect 8991 12600 9036 12628
rect 9030 12588 9036 12600
rect 9088 12628 9094 12640
rect 9490 12628 9496 12640
rect 9088 12600 9496 12628
rect 9088 12588 9094 12600
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 9766 12588 9772 12640
rect 9824 12628 9830 12640
rect 10796 12628 10824 12656
rect 9824 12600 10824 12628
rect 12897 12631 12955 12637
rect 9824 12588 9830 12600
rect 12897 12597 12909 12631
rect 12943 12628 12955 12631
rect 13170 12628 13176 12640
rect 12943 12600 13176 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 13170 12588 13176 12600
rect 13228 12628 13234 12640
rect 14936 12628 14964 12656
rect 13228 12600 14964 12628
rect 13228 12588 13234 12600
rect 1104 12538 16008 12560
rect 1104 12486 2824 12538
rect 2876 12486 2888 12538
rect 2940 12486 2952 12538
rect 3004 12486 3016 12538
rect 3068 12486 3080 12538
rect 3132 12486 6572 12538
rect 6624 12486 6636 12538
rect 6688 12486 6700 12538
rect 6752 12486 6764 12538
rect 6816 12486 6828 12538
rect 6880 12486 10320 12538
rect 10372 12486 10384 12538
rect 10436 12486 10448 12538
rect 10500 12486 10512 12538
rect 10564 12486 10576 12538
rect 10628 12486 14068 12538
rect 14120 12486 14132 12538
rect 14184 12486 14196 12538
rect 14248 12486 14260 12538
rect 14312 12486 14324 12538
rect 14376 12486 16008 12538
rect 1104 12464 16008 12486
rect 2869 12427 2927 12433
rect 2869 12393 2881 12427
rect 2915 12424 2927 12427
rect 3142 12424 3148 12436
rect 2915 12396 3148 12424
rect 2915 12393 2927 12396
rect 2869 12387 2927 12393
rect 3142 12384 3148 12396
rect 3200 12384 3206 12436
rect 6362 12384 6368 12436
rect 6420 12424 6426 12436
rect 6733 12427 6791 12433
rect 6733 12424 6745 12427
rect 6420 12396 6745 12424
rect 6420 12384 6426 12396
rect 6733 12393 6745 12396
rect 6779 12393 6791 12427
rect 6733 12387 6791 12393
rect 7834 12384 7840 12436
rect 7892 12424 7898 12436
rect 8941 12427 8999 12433
rect 8941 12424 8953 12427
rect 7892 12396 8953 12424
rect 7892 12384 7898 12396
rect 8941 12393 8953 12396
rect 8987 12393 8999 12427
rect 10870 12424 10876 12436
rect 10831 12396 10876 12424
rect 8941 12387 8999 12393
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 14093 12427 14151 12433
rect 14093 12424 14105 12427
rect 13872 12396 14105 12424
rect 13872 12384 13878 12396
rect 14093 12393 14105 12396
rect 14139 12393 14151 12427
rect 15562 12424 15568 12436
rect 15523 12396 15568 12424
rect 14093 12387 14151 12393
rect 15562 12384 15568 12396
rect 15620 12384 15626 12436
rect 3694 12356 3700 12368
rect 3344 12328 3700 12356
rect 3344 12297 3372 12328
rect 3694 12316 3700 12328
rect 3752 12356 3758 12368
rect 5258 12356 5264 12368
rect 3752 12328 5264 12356
rect 3752 12316 3758 12328
rect 5258 12316 5264 12328
rect 5316 12316 5322 12368
rect 11054 12316 11060 12368
rect 11112 12316 11118 12368
rect 12894 12316 12900 12368
rect 12952 12356 12958 12368
rect 15473 12359 15531 12365
rect 12952 12328 14596 12356
rect 12952 12316 12958 12328
rect 1765 12291 1823 12297
rect 1765 12257 1777 12291
rect 1811 12257 1823 12291
rect 1765 12251 1823 12257
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12288 2835 12291
rect 3329 12291 3387 12297
rect 3329 12288 3341 12291
rect 2823 12260 3341 12288
rect 2823 12257 2835 12260
rect 2777 12251 2835 12257
rect 3329 12257 3341 12260
rect 3375 12257 3387 12291
rect 3329 12251 3387 12257
rect 3513 12291 3571 12297
rect 3513 12257 3525 12291
rect 3559 12288 3571 12291
rect 4154 12288 4160 12300
rect 3559 12260 4160 12288
rect 3559 12257 3571 12260
rect 3513 12251 3571 12257
rect 1780 12152 1808 12251
rect 4154 12248 4160 12260
rect 4212 12248 4218 12300
rect 11072 12288 11100 12316
rect 14568 12300 14596 12328
rect 15473 12325 15485 12359
rect 15519 12356 15531 12359
rect 15838 12356 15844 12368
rect 15519 12328 15844 12356
rect 15519 12325 15531 12328
rect 15473 12319 15531 12325
rect 15838 12316 15844 12328
rect 15896 12316 15902 12368
rect 10244 12260 11100 12288
rect 12621 12291 12679 12297
rect 2593 12223 2651 12229
rect 2593 12189 2605 12223
rect 2639 12220 2651 12223
rect 3878 12220 3884 12232
rect 2639 12192 3884 12220
rect 2639 12189 2651 12192
rect 2593 12183 2651 12189
rect 3878 12180 3884 12192
rect 3936 12180 3942 12232
rect 4617 12223 4675 12229
rect 4617 12189 4629 12223
rect 4663 12220 4675 12223
rect 4798 12220 4804 12232
rect 4663 12192 4804 12220
rect 4663 12189 4675 12192
rect 4617 12183 4675 12189
rect 4798 12180 4804 12192
rect 4856 12220 4862 12232
rect 4985 12223 5043 12229
rect 4985 12220 4997 12223
rect 4856 12192 4997 12220
rect 4856 12180 4862 12192
rect 4985 12189 4997 12192
rect 5031 12220 5043 12223
rect 5169 12223 5227 12229
rect 5169 12220 5181 12223
rect 5031 12192 5181 12220
rect 5031 12189 5043 12192
rect 4985 12183 5043 12189
rect 5169 12189 5181 12192
rect 5215 12220 5227 12223
rect 5445 12223 5503 12229
rect 5445 12220 5457 12223
rect 5215 12192 5457 12220
rect 5215 12189 5227 12192
rect 5169 12183 5227 12189
rect 5445 12189 5457 12192
rect 5491 12220 5503 12223
rect 6454 12220 6460 12232
rect 5491 12192 6460 12220
rect 5491 12189 5503 12192
rect 5445 12183 5503 12189
rect 6454 12180 6460 12192
rect 6512 12220 6518 12232
rect 6641 12223 6699 12229
rect 6641 12220 6653 12223
rect 6512 12192 6653 12220
rect 6512 12180 6518 12192
rect 6641 12189 6653 12192
rect 6687 12220 6699 12223
rect 8113 12223 8171 12229
rect 8113 12220 8125 12223
rect 6687 12192 8125 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 8113 12189 8125 12192
rect 8159 12189 8171 12223
rect 8113 12183 8171 12189
rect 4522 12152 4528 12164
rect 1780 12124 4528 12152
rect 4522 12112 4528 12124
rect 4580 12112 4586 12164
rect 7868 12155 7926 12161
rect 7868 12121 7880 12155
rect 7914 12152 7926 12155
rect 8128 12152 8156 12183
rect 9490 12180 9496 12232
rect 9548 12220 9554 12232
rect 10065 12223 10123 12229
rect 10065 12220 10077 12223
rect 9548 12192 10077 12220
rect 9548 12180 9554 12192
rect 10065 12189 10077 12192
rect 10111 12220 10123 12223
rect 10244 12220 10272 12260
rect 12621 12257 12633 12291
rect 12667 12288 12679 12291
rect 13078 12288 13084 12300
rect 12667 12260 13084 12288
rect 12667 12257 12679 12260
rect 12621 12251 12679 12257
rect 13078 12248 13084 12260
rect 13136 12248 13142 12300
rect 13357 12291 13415 12297
rect 13357 12257 13369 12291
rect 13403 12257 13415 12291
rect 13357 12251 13415 12257
rect 10111 12192 10272 12220
rect 10321 12223 10379 12229
rect 10111 12189 10123 12192
rect 10065 12183 10123 12189
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 10870 12220 10876 12232
rect 10367 12192 10876 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 10870 12180 10876 12192
rect 10928 12220 10934 12232
rect 11057 12223 11115 12229
rect 11057 12220 11069 12223
rect 10928 12192 11069 12220
rect 10928 12180 10934 12192
rect 11057 12189 11069 12192
rect 11103 12189 11115 12223
rect 11057 12183 11115 12189
rect 11330 12180 11336 12232
rect 11388 12220 11394 12232
rect 13265 12223 13323 12229
rect 13265 12220 13277 12223
rect 11388 12192 13277 12220
rect 11388 12180 11394 12192
rect 13265 12189 13277 12192
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 13372 12220 13400 12251
rect 13446 12248 13452 12300
rect 13504 12288 13510 12300
rect 13817 12291 13875 12297
rect 13817 12288 13829 12291
rect 13504 12260 13829 12288
rect 13504 12248 13510 12260
rect 13817 12257 13829 12260
rect 13863 12257 13875 12291
rect 14550 12288 14556 12300
rect 14511 12260 14556 12288
rect 13817 12251 13875 12257
rect 14550 12248 14556 12260
rect 14608 12248 14614 12300
rect 14737 12291 14795 12297
rect 14737 12257 14749 12291
rect 14783 12288 14795 12291
rect 14918 12288 14924 12300
rect 14783 12260 14924 12288
rect 14783 12257 14795 12260
rect 14737 12251 14795 12257
rect 14918 12248 14924 12260
rect 14976 12248 14982 12300
rect 15289 12291 15347 12297
rect 15289 12257 15301 12291
rect 15335 12288 15347 12291
rect 15930 12288 15936 12300
rect 15335 12260 15936 12288
rect 15335 12257 15347 12260
rect 15289 12251 15347 12257
rect 15930 12248 15936 12260
rect 15988 12248 15994 12300
rect 14642 12220 14648 12232
rect 13372 12192 14648 12220
rect 8757 12155 8815 12161
rect 8757 12152 8769 12155
rect 7914 12124 8064 12152
rect 8128 12124 8769 12152
rect 7914 12121 7926 12124
rect 7868 12115 7926 12121
rect 1854 12084 1860 12096
rect 1815 12056 1860 12084
rect 1854 12044 1860 12056
rect 1912 12044 1918 12096
rect 1949 12087 2007 12093
rect 1949 12053 1961 12087
rect 1995 12084 2007 12087
rect 2038 12084 2044 12096
rect 1995 12056 2044 12084
rect 1995 12053 2007 12056
rect 1949 12047 2007 12053
rect 2038 12044 2044 12056
rect 2096 12044 2102 12096
rect 2314 12084 2320 12096
rect 2275 12056 2320 12084
rect 2314 12044 2320 12056
rect 2372 12044 2378 12096
rect 3234 12084 3240 12096
rect 3195 12056 3240 12084
rect 3234 12044 3240 12056
rect 3292 12044 3298 12096
rect 3970 12044 3976 12096
rect 4028 12084 4034 12096
rect 5718 12084 5724 12096
rect 4028 12056 5724 12084
rect 4028 12044 4034 12056
rect 5718 12044 5724 12056
rect 5776 12044 5782 12096
rect 8036 12084 8064 12124
rect 8757 12121 8769 12124
rect 8803 12152 8815 12155
rect 9214 12152 9220 12164
rect 8803 12124 9220 12152
rect 8803 12121 8815 12124
rect 8757 12115 8815 12121
rect 9214 12112 9220 12124
rect 9272 12112 9278 12164
rect 11790 12152 11796 12164
rect 11072 12124 11796 12152
rect 11072 12084 11100 12124
rect 11790 12112 11796 12124
rect 11848 12112 11854 12164
rect 12342 12152 12348 12164
rect 12400 12161 12406 12164
rect 12312 12124 12348 12152
rect 12342 12112 12348 12124
rect 12400 12115 12412 12161
rect 13372 12152 13400 12192
rect 14642 12180 14648 12192
rect 14700 12180 14706 12232
rect 12636 12124 13400 12152
rect 14461 12155 14519 12161
rect 12400 12112 12406 12115
rect 11238 12084 11244 12096
rect 8036 12056 11100 12084
rect 11199 12056 11244 12084
rect 11238 12044 11244 12056
rect 11296 12044 11302 12096
rect 11330 12044 11336 12096
rect 11388 12084 11394 12096
rect 12636 12084 12664 12124
rect 14461 12121 14473 12155
rect 14507 12152 14519 12155
rect 14921 12155 14979 12161
rect 14921 12152 14933 12155
rect 14507 12124 14933 12152
rect 14507 12121 14519 12124
rect 14461 12115 14519 12121
rect 14921 12121 14933 12124
rect 14967 12121 14979 12155
rect 14921 12115 14979 12121
rect 12802 12084 12808 12096
rect 11388 12056 12664 12084
rect 12763 12056 12808 12084
rect 11388 12044 11394 12056
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 13173 12087 13231 12093
rect 13173 12053 13185 12087
rect 13219 12084 13231 12087
rect 13722 12084 13728 12096
rect 13219 12056 13728 12084
rect 13219 12053 13231 12056
rect 13173 12047 13231 12053
rect 13722 12044 13728 12056
rect 13780 12044 13786 12096
rect 1104 11994 16008 12016
rect 1104 11942 4698 11994
rect 4750 11942 4762 11994
rect 4814 11942 4826 11994
rect 4878 11942 4890 11994
rect 4942 11942 4954 11994
rect 5006 11942 8446 11994
rect 8498 11942 8510 11994
rect 8562 11942 8574 11994
rect 8626 11942 8638 11994
rect 8690 11942 8702 11994
rect 8754 11942 12194 11994
rect 12246 11942 12258 11994
rect 12310 11942 12322 11994
rect 12374 11942 12386 11994
rect 12438 11942 12450 11994
rect 12502 11942 16008 11994
rect 1104 11920 16008 11942
rect 1486 11880 1492 11892
rect 1447 11852 1492 11880
rect 1486 11840 1492 11852
rect 1544 11840 1550 11892
rect 2590 11880 2596 11892
rect 2551 11852 2596 11880
rect 2590 11840 2596 11852
rect 2648 11840 2654 11892
rect 4065 11883 4123 11889
rect 4065 11849 4077 11883
rect 4111 11880 4123 11883
rect 4154 11880 4160 11892
rect 4111 11852 4160 11880
rect 4111 11849 4123 11852
rect 4065 11843 4123 11849
rect 4154 11840 4160 11852
rect 4212 11840 4218 11892
rect 4338 11840 4344 11892
rect 4396 11880 4402 11892
rect 9490 11880 9496 11892
rect 4396 11852 5304 11880
rect 9451 11852 9496 11880
rect 4396 11840 4402 11852
rect 2406 11772 2412 11824
rect 2464 11812 2470 11824
rect 2501 11815 2559 11821
rect 2501 11812 2513 11815
rect 2464 11784 2513 11812
rect 2464 11772 2470 11784
rect 2501 11781 2513 11784
rect 2547 11781 2559 11815
rect 3970 11812 3976 11824
rect 2501 11775 2559 11781
rect 3344 11784 3976 11812
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 1949 11747 2007 11753
rect 1719 11716 1808 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 1780 11617 1808 11716
rect 1949 11713 1961 11747
rect 1995 11744 2007 11747
rect 2314 11744 2320 11756
rect 1995 11716 2320 11744
rect 1995 11713 2007 11716
rect 1949 11707 2007 11713
rect 2314 11704 2320 11716
rect 2372 11704 2378 11756
rect 3142 11704 3148 11756
rect 3200 11744 3206 11756
rect 3344 11753 3372 11784
rect 3970 11772 3976 11784
rect 4028 11772 4034 11824
rect 4522 11772 4528 11824
rect 4580 11812 4586 11824
rect 5178 11815 5236 11821
rect 5178 11812 5190 11815
rect 4580 11784 5190 11812
rect 4580 11772 4586 11784
rect 5178 11781 5190 11784
rect 5224 11781 5236 11815
rect 5276 11812 5304 11852
rect 9490 11840 9496 11852
rect 9548 11840 9554 11892
rect 9950 11840 9956 11892
rect 10008 11880 10014 11892
rect 11330 11880 11336 11892
rect 10008 11852 11336 11880
rect 10008 11840 10014 11852
rect 11330 11840 11336 11852
rect 11388 11840 11394 11892
rect 11698 11840 11704 11892
rect 11756 11880 11762 11892
rect 12713 11883 12771 11889
rect 12713 11880 12725 11883
rect 11756 11852 12725 11880
rect 11756 11840 11762 11852
rect 12713 11849 12725 11852
rect 12759 11849 12771 11883
rect 12986 11880 12992 11892
rect 12947 11852 12992 11880
rect 12713 11843 12771 11849
rect 12986 11840 12992 11852
rect 13044 11840 13050 11892
rect 13170 11880 13176 11892
rect 13131 11852 13176 11880
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 13814 11880 13820 11892
rect 13775 11852 13820 11880
rect 13814 11840 13820 11852
rect 13872 11880 13878 11892
rect 14369 11883 14427 11889
rect 14369 11880 14381 11883
rect 13872 11852 14381 11880
rect 13872 11840 13878 11852
rect 14369 11849 14381 11852
rect 14415 11849 14427 11883
rect 14369 11843 14427 11849
rect 14458 11840 14464 11892
rect 14516 11880 14522 11892
rect 14553 11883 14611 11889
rect 14553 11880 14565 11883
rect 14516 11852 14565 11880
rect 14516 11840 14522 11852
rect 14553 11849 14565 11852
rect 14599 11849 14611 11883
rect 14734 11880 14740 11892
rect 14695 11852 14740 11880
rect 14553 11843 14611 11849
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 15286 11840 15292 11892
rect 15344 11880 15350 11892
rect 15565 11883 15623 11889
rect 15565 11880 15577 11883
rect 15344 11852 15577 11880
rect 15344 11840 15350 11852
rect 15565 11849 15577 11852
rect 15611 11849 15623 11883
rect 15565 11843 15623 11849
rect 10628 11815 10686 11821
rect 5276 11784 10364 11812
rect 5178 11775 5236 11781
rect 3329 11747 3387 11753
rect 3329 11744 3341 11747
rect 3200 11716 3341 11744
rect 3200 11704 3206 11716
rect 3329 11713 3341 11716
rect 3375 11713 3387 11747
rect 3329 11707 3387 11713
rect 3421 11747 3479 11753
rect 3421 11713 3433 11747
rect 3467 11744 3479 11747
rect 4062 11744 4068 11756
rect 3467 11716 4068 11744
rect 3467 11713 3479 11716
rect 3421 11707 3479 11713
rect 4062 11704 4068 11716
rect 4120 11744 4126 11756
rect 10226 11744 10232 11756
rect 4120 11716 10232 11744
rect 4120 11704 4126 11716
rect 10226 11704 10232 11716
rect 10284 11704 10290 11756
rect 10336 11744 10364 11784
rect 10628 11781 10640 11815
rect 10674 11812 10686 11815
rect 11238 11812 11244 11824
rect 10674 11784 11244 11812
rect 10674 11781 10686 11784
rect 10628 11775 10686 11781
rect 11238 11772 11244 11784
rect 11296 11772 11302 11824
rect 12253 11815 12311 11821
rect 12253 11781 12265 11815
rect 12299 11812 12311 11815
rect 12299 11784 12756 11812
rect 12299 11781 12311 11784
rect 12253 11775 12311 11781
rect 12728 11756 12756 11784
rect 12345 11747 12403 11753
rect 10336 11716 11008 11744
rect 2777 11679 2835 11685
rect 2777 11645 2789 11679
rect 2823 11676 2835 11679
rect 3510 11676 3516 11688
rect 2823 11648 3516 11676
rect 2823 11645 2835 11648
rect 2777 11639 2835 11645
rect 3510 11636 3516 11648
rect 3568 11636 3574 11688
rect 5442 11636 5448 11688
rect 5500 11676 5506 11688
rect 10870 11676 10876 11688
rect 5500 11648 5672 11676
rect 10831 11648 10876 11676
rect 5500 11636 5506 11648
rect 1765 11611 1823 11617
rect 1765 11577 1777 11611
rect 1811 11577 1823 11611
rect 1765 11571 1823 11577
rect 2130 11540 2136 11552
rect 2091 11512 2136 11540
rect 2130 11500 2136 11512
rect 2188 11500 2194 11552
rect 2498 11500 2504 11552
rect 2556 11540 2562 11552
rect 2961 11543 3019 11549
rect 2961 11540 2973 11543
rect 2556 11512 2973 11540
rect 2556 11500 2562 11512
rect 2961 11509 2973 11512
rect 3007 11509 3019 11543
rect 2961 11503 3019 11509
rect 3234 11500 3240 11552
rect 3292 11540 3298 11552
rect 5644 11549 5672 11648
rect 10870 11636 10876 11648
rect 10928 11636 10934 11688
rect 10980 11608 11008 11716
rect 12345 11713 12357 11747
rect 12391 11744 12403 11747
rect 12618 11744 12624 11756
rect 12391 11716 12624 11744
rect 12391 11713 12403 11716
rect 12345 11707 12403 11713
rect 12618 11704 12624 11716
rect 12676 11704 12682 11756
rect 12710 11704 12716 11756
rect 12768 11704 12774 11756
rect 12066 11636 12072 11688
rect 12124 11676 12130 11688
rect 12437 11679 12495 11685
rect 12437 11676 12449 11679
rect 12124 11648 12449 11676
rect 12124 11636 12130 11648
rect 12437 11645 12449 11648
rect 12483 11645 12495 11679
rect 13188 11676 13216 11840
rect 13538 11772 13544 11824
rect 13596 11812 13602 11824
rect 14921 11815 14979 11821
rect 14921 11812 14933 11815
rect 13596 11784 14933 11812
rect 13596 11772 13602 11784
rect 14921 11781 14933 11784
rect 14967 11781 14979 11815
rect 14921 11775 14979 11781
rect 15381 11815 15439 11821
rect 15381 11781 15393 11815
rect 15427 11812 15439 11815
rect 15746 11812 15752 11824
rect 15427 11784 15752 11812
rect 15427 11781 15439 11784
rect 15381 11775 15439 11781
rect 15746 11772 15752 11784
rect 15804 11772 15810 11824
rect 13725 11747 13783 11753
rect 13725 11713 13737 11747
rect 13771 11744 13783 11747
rect 15197 11747 15255 11753
rect 13771 11716 14780 11744
rect 13771 11713 13783 11716
rect 13725 11707 13783 11713
rect 14001 11679 14059 11685
rect 13188 11648 13952 11676
rect 12437 11639 12495 11645
rect 13814 11608 13820 11620
rect 10980 11580 13820 11608
rect 13814 11568 13820 11580
rect 13872 11568 13878 11620
rect 13924 11552 13952 11648
rect 14001 11645 14013 11679
rect 14047 11676 14059 11679
rect 14642 11676 14648 11688
rect 14047 11648 14648 11676
rect 14047 11645 14059 11648
rect 14001 11639 14059 11645
rect 14642 11636 14648 11648
rect 14700 11636 14706 11688
rect 3881 11543 3939 11549
rect 3881 11540 3893 11543
rect 3292 11512 3893 11540
rect 3292 11500 3298 11512
rect 3881 11509 3893 11512
rect 3927 11509 3939 11543
rect 3881 11503 3939 11509
rect 5629 11543 5687 11549
rect 5629 11509 5641 11543
rect 5675 11540 5687 11543
rect 5813 11543 5871 11549
rect 5813 11540 5825 11543
rect 5675 11512 5825 11540
rect 5675 11509 5687 11512
rect 5629 11503 5687 11509
rect 5813 11509 5825 11512
rect 5859 11540 5871 11543
rect 5997 11543 6055 11549
rect 5997 11540 6009 11543
rect 5859 11512 6009 11540
rect 5859 11509 5871 11512
rect 5813 11503 5871 11509
rect 5997 11509 6009 11512
rect 6043 11540 6055 11543
rect 7285 11543 7343 11549
rect 7285 11540 7297 11543
rect 6043 11512 7297 11540
rect 6043 11509 6055 11512
rect 5997 11503 6055 11509
rect 7285 11509 7297 11512
rect 7331 11540 7343 11543
rect 9214 11540 9220 11552
rect 7331 11512 9220 11540
rect 7331 11509 7343 11512
rect 7285 11503 7343 11509
rect 9214 11500 9220 11512
rect 9272 11540 9278 11552
rect 9309 11543 9367 11549
rect 9309 11540 9321 11543
rect 9272 11512 9321 11540
rect 9272 11500 9278 11512
rect 9309 11509 9321 11512
rect 9355 11509 9367 11543
rect 9309 11503 9367 11509
rect 11054 11500 11060 11552
rect 11112 11540 11118 11552
rect 11885 11543 11943 11549
rect 11885 11540 11897 11543
rect 11112 11512 11897 11540
rect 11112 11500 11118 11512
rect 11885 11509 11897 11512
rect 11931 11509 11943 11543
rect 13354 11540 13360 11552
rect 13315 11512 13360 11540
rect 11885 11503 11943 11509
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 13906 11500 13912 11552
rect 13964 11500 13970 11552
rect 14277 11543 14335 11549
rect 14277 11509 14289 11543
rect 14323 11540 14335 11543
rect 14752 11540 14780 11716
rect 15197 11713 15209 11747
rect 15243 11744 15255 11747
rect 16022 11744 16028 11756
rect 15243 11716 16028 11744
rect 15243 11713 15255 11716
rect 15197 11707 15255 11713
rect 16022 11704 16028 11716
rect 16080 11704 16086 11756
rect 15194 11540 15200 11552
rect 14323 11512 15200 11540
rect 14323 11509 14335 11512
rect 14277 11503 14335 11509
rect 15194 11500 15200 11512
rect 15252 11500 15258 11552
rect 1104 11450 16008 11472
rect 1104 11398 2824 11450
rect 2876 11398 2888 11450
rect 2940 11398 2952 11450
rect 3004 11398 3016 11450
rect 3068 11398 3080 11450
rect 3132 11398 6572 11450
rect 6624 11398 6636 11450
rect 6688 11398 6700 11450
rect 6752 11398 6764 11450
rect 6816 11398 6828 11450
rect 6880 11398 10320 11450
rect 10372 11398 10384 11450
rect 10436 11398 10448 11450
rect 10500 11398 10512 11450
rect 10564 11398 10576 11450
rect 10628 11398 14068 11450
rect 14120 11398 14132 11450
rect 14184 11398 14196 11450
rect 14248 11398 14260 11450
rect 14312 11398 14324 11450
rect 14376 11398 16008 11450
rect 1104 11376 16008 11398
rect 2038 11336 2044 11348
rect 1999 11308 2044 11336
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 5810 11336 5816 11348
rect 3252 11308 5816 11336
rect 2869 11271 2927 11277
rect 2869 11268 2881 11271
rect 2424 11240 2881 11268
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11132 1731 11135
rect 1762 11132 1768 11144
rect 1719 11104 1768 11132
rect 1719 11101 1731 11104
rect 1673 11095 1731 11101
rect 1762 11092 1768 11104
rect 1820 11092 1826 11144
rect 2424 11141 2452 11240
rect 2869 11237 2881 11240
rect 2915 11237 2927 11271
rect 2869 11231 2927 11237
rect 2498 11160 2504 11212
rect 2556 11200 2562 11212
rect 2685 11203 2743 11209
rect 2556 11172 2601 11200
rect 2556 11160 2562 11172
rect 2685 11169 2697 11203
rect 2731 11200 2743 11203
rect 3252 11200 3280 11308
rect 5810 11296 5816 11308
rect 5868 11296 5874 11348
rect 7282 11336 7288 11348
rect 7243 11308 7288 11336
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 8757 11339 8815 11345
rect 8757 11305 8769 11339
rect 8803 11336 8815 11339
rect 9490 11336 9496 11348
rect 8803 11308 9496 11336
rect 8803 11305 8815 11308
rect 8757 11299 8815 11305
rect 9490 11296 9496 11308
rect 9548 11296 9554 11348
rect 10134 11296 10140 11348
rect 10192 11336 10198 11348
rect 10505 11339 10563 11345
rect 10505 11336 10517 11339
rect 10192 11308 10517 11336
rect 10192 11296 10198 11308
rect 10505 11305 10517 11308
rect 10551 11305 10563 11339
rect 10870 11336 10876 11348
rect 10505 11299 10563 11305
rect 10612 11308 10876 11336
rect 3344 11240 3740 11268
rect 3344 11209 3372 11240
rect 2731 11172 3280 11200
rect 3329 11203 3387 11209
rect 2731 11169 2743 11172
rect 2685 11163 2743 11169
rect 3329 11169 3341 11203
rect 3375 11169 3387 11203
rect 3329 11163 3387 11169
rect 2409 11135 2467 11141
rect 2409 11101 2421 11135
rect 2455 11101 2467 11135
rect 2409 11095 2467 11101
rect 2590 11092 2596 11144
rect 2648 11132 2654 11144
rect 2700 11132 2728 11163
rect 3510 11160 3516 11212
rect 3568 11200 3574 11212
rect 3712 11200 3740 11240
rect 4062 11228 4068 11280
rect 4120 11268 4126 11280
rect 4249 11271 4307 11277
rect 4249 11268 4261 11271
rect 4120 11240 4261 11268
rect 4120 11228 4126 11240
rect 4249 11237 4261 11240
rect 4295 11237 4307 11271
rect 4249 11231 4307 11237
rect 4338 11200 4344 11212
rect 3568 11172 3613 11200
rect 3712 11172 4344 11200
rect 3568 11160 3574 11172
rect 4338 11160 4344 11172
rect 4396 11160 4402 11212
rect 2648 11104 2728 11132
rect 3528 11132 3556 11160
rect 3528 11104 3924 11132
rect 2648 11092 2654 11104
rect 3237 11067 3295 11073
rect 3237 11033 3249 11067
rect 3283 11064 3295 11067
rect 3789 11067 3847 11073
rect 3789 11064 3801 11067
rect 3283 11036 3801 11064
rect 3283 11033 3295 11036
rect 3237 11027 3295 11033
rect 3789 11033 3801 11036
rect 3835 11033 3847 11067
rect 3896 11064 3924 11104
rect 3970 11092 3976 11144
rect 4028 11132 4034 11144
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 4028 11104 4077 11132
rect 4028 11092 4034 11104
rect 4065 11101 4077 11104
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11132 4491 11135
rect 5442 11132 5448 11144
rect 4479 11104 5448 11132
rect 4479 11101 4491 11104
rect 4433 11095 4491 11101
rect 5442 11092 5448 11104
rect 5500 11132 5506 11144
rect 5905 11135 5963 11141
rect 5905 11132 5917 11135
rect 5500 11104 5917 11132
rect 5500 11092 5506 11104
rect 5905 11101 5917 11104
rect 5951 11101 5963 11135
rect 5905 11095 5963 11101
rect 6172 11135 6230 11141
rect 6172 11101 6184 11135
rect 6218 11101 6230 11135
rect 6172 11095 6230 11101
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11132 7435 11135
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 7423 11104 9137 11132
rect 7423 11101 7435 11104
rect 7377 11095 7435 11101
rect 4678 11067 4736 11073
rect 4678 11064 4690 11067
rect 3896 11036 4690 11064
rect 3789 11027 3847 11033
rect 4678 11033 4690 11036
rect 4724 11033 4736 11067
rect 4678 11027 4736 11033
rect 6086 11024 6092 11076
rect 6144 11064 6150 11076
rect 6196 11064 6224 11095
rect 6144 11036 6224 11064
rect 7644 11067 7702 11073
rect 6144 11024 6150 11036
rect 7644 11033 7656 11067
rect 7690 11064 7702 11067
rect 8846 11064 8852 11076
rect 7690 11036 8852 11064
rect 7690 11033 7702 11036
rect 7644 11027 7702 11033
rect 8846 11024 8852 11036
rect 8904 11024 8910 11076
rect 8956 11008 8984 11104
rect 9125 11101 9137 11104
rect 9171 11132 9183 11135
rect 9214 11132 9220 11144
rect 9171 11104 9220 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 9214 11092 9220 11104
rect 9272 11132 9278 11144
rect 10612 11141 10640 11308
rect 10870 11296 10876 11308
rect 10928 11336 10934 11348
rect 12526 11336 12532 11348
rect 10928 11308 12532 11336
rect 10928 11296 10934 11308
rect 12526 11296 12532 11308
rect 12584 11336 12590 11348
rect 15197 11339 15255 11345
rect 12584 11308 13492 11336
rect 12584 11296 12590 11308
rect 13464 11209 13492 11308
rect 15197 11305 15209 11339
rect 15243 11336 15255 11339
rect 15286 11336 15292 11348
rect 15243 11308 15292 11336
rect 15243 11305 15255 11308
rect 15197 11299 15255 11305
rect 15286 11296 15292 11308
rect 15344 11336 15350 11348
rect 16298 11336 16304 11348
rect 15344 11308 16304 11336
rect 15344 11296 15350 11308
rect 16298 11296 16304 11308
rect 16356 11296 16362 11348
rect 13449 11203 13507 11209
rect 13449 11169 13461 11203
rect 13495 11169 13507 11203
rect 14642 11200 14648 11212
rect 14603 11172 14648 11200
rect 13449 11163 13507 11169
rect 14642 11160 14648 11172
rect 14700 11160 14706 11212
rect 15194 11160 15200 11212
rect 15252 11160 15258 11212
rect 10597 11135 10655 11141
rect 10597 11132 10609 11135
rect 9272 11104 10609 11132
rect 9272 11092 9278 11104
rect 10597 11101 10609 11104
rect 10643 11101 10655 11135
rect 15212 11132 15240 11160
rect 16022 11132 16028 11144
rect 10597 11095 10655 11101
rect 10704 11104 16028 11132
rect 9392 11067 9450 11073
rect 9392 11033 9404 11067
rect 9438 11064 9450 11067
rect 9582 11064 9588 11076
rect 9438 11036 9588 11064
rect 9438 11033 9450 11036
rect 9392 11027 9450 11033
rect 9582 11024 9588 11036
rect 9640 11024 9646 11076
rect 10704 11064 10732 11104
rect 16022 11092 16028 11104
rect 16080 11092 16086 11144
rect 10853 11067 10911 11073
rect 10853 11064 10865 11067
rect 9692 11036 10732 11064
rect 10796 11036 10865 11064
rect 1486 10996 1492 11008
rect 1447 10968 1492 10996
rect 1486 10956 1492 10968
rect 1544 10956 1550 11008
rect 3142 10956 3148 11008
rect 3200 10996 3206 11008
rect 3326 10996 3332 11008
rect 3200 10968 3332 10996
rect 3200 10956 3206 10968
rect 3326 10956 3332 10968
rect 3384 10956 3390 11008
rect 8938 10996 8944 11008
rect 8899 10968 8944 10996
rect 8938 10956 8944 10968
rect 8996 10956 9002 11008
rect 9306 10956 9312 11008
rect 9364 10996 9370 11008
rect 9692 10996 9720 11036
rect 9364 10968 9720 10996
rect 9364 10956 9370 10968
rect 9950 10956 9956 11008
rect 10008 10996 10014 11008
rect 10796 10996 10824 11036
rect 10853 11033 10865 11036
rect 10899 11033 10911 11067
rect 13182 11067 13240 11073
rect 13182 11064 13194 11067
rect 10853 11027 10911 11033
rect 11992 11036 13194 11064
rect 10008 10968 10824 10996
rect 10008 10956 10014 10968
rect 11882 10956 11888 11008
rect 11940 10996 11946 11008
rect 11992 11005 12020 11036
rect 13182 11033 13194 11036
rect 13228 11033 13240 11067
rect 13182 11027 13240 11033
rect 13909 11067 13967 11073
rect 13909 11033 13921 11067
rect 13955 11064 13967 11067
rect 14461 11067 14519 11073
rect 14461 11064 14473 11067
rect 13955 11036 14473 11064
rect 13955 11033 13967 11036
rect 13909 11027 13967 11033
rect 14461 11033 14473 11036
rect 14507 11033 14519 11067
rect 14461 11027 14519 11033
rect 14550 11024 14556 11076
rect 14608 11064 14614 11076
rect 14921 11067 14979 11073
rect 14921 11064 14933 11067
rect 14608 11036 14933 11064
rect 14608 11024 14614 11036
rect 14921 11033 14933 11036
rect 14967 11033 14979 11067
rect 14921 11027 14979 11033
rect 15194 11024 15200 11076
rect 15252 11064 15258 11076
rect 15289 11067 15347 11073
rect 15289 11064 15301 11067
rect 15252 11036 15301 11064
rect 15252 11024 15258 11036
rect 15289 11033 15301 11036
rect 15335 11064 15347 11067
rect 15378 11064 15384 11076
rect 15335 11036 15384 11064
rect 15335 11033 15347 11036
rect 15289 11027 15347 11033
rect 15378 11024 15384 11036
rect 15436 11024 15442 11076
rect 11977 10999 12035 11005
rect 11977 10996 11989 10999
rect 11940 10968 11989 10996
rect 11940 10956 11946 10968
rect 11977 10965 11989 10968
rect 12023 10965 12035 10999
rect 11977 10959 12035 10965
rect 12066 10956 12072 11008
rect 12124 10996 12130 11008
rect 14090 10996 14096 11008
rect 12124 10968 12169 10996
rect 14051 10968 14096 10996
rect 12124 10956 12130 10968
rect 14090 10956 14096 10968
rect 14148 10956 14154 11008
rect 14642 10956 14648 11008
rect 14700 10996 14706 11008
rect 15010 10996 15016 11008
rect 14700 10968 15016 10996
rect 14700 10956 14706 10968
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 1104 10906 16008 10928
rect 1104 10854 4698 10906
rect 4750 10854 4762 10906
rect 4814 10854 4826 10906
rect 4878 10854 4890 10906
rect 4942 10854 4954 10906
rect 5006 10854 8446 10906
rect 8498 10854 8510 10906
rect 8562 10854 8574 10906
rect 8626 10854 8638 10906
rect 8690 10854 8702 10906
rect 8754 10854 12194 10906
rect 12246 10854 12258 10906
rect 12310 10854 12322 10906
rect 12374 10854 12386 10906
rect 12438 10854 12450 10906
rect 12502 10854 16008 10906
rect 1104 10832 16008 10854
rect 1854 10792 1860 10804
rect 1815 10764 1860 10792
rect 1854 10752 1860 10764
rect 1912 10752 1918 10804
rect 2130 10752 2136 10804
rect 2188 10792 2194 10804
rect 2225 10795 2283 10801
rect 2225 10792 2237 10795
rect 2188 10764 2237 10792
rect 2188 10752 2194 10764
rect 2225 10761 2237 10764
rect 2271 10761 2283 10795
rect 2225 10755 2283 10761
rect 2317 10795 2375 10801
rect 2317 10761 2329 10795
rect 2363 10792 2375 10795
rect 2685 10795 2743 10801
rect 2685 10792 2697 10795
rect 2363 10764 2697 10792
rect 2363 10761 2375 10764
rect 2317 10755 2375 10761
rect 2685 10761 2697 10764
rect 2731 10761 2743 10795
rect 2685 10755 2743 10761
rect 3145 10795 3203 10801
rect 3145 10761 3157 10795
rect 3191 10792 3203 10795
rect 3513 10795 3571 10801
rect 3513 10792 3525 10795
rect 3191 10764 3525 10792
rect 3191 10761 3203 10764
rect 3145 10755 3203 10761
rect 3513 10761 3525 10764
rect 3559 10761 3571 10795
rect 4338 10792 4344 10804
rect 4299 10764 4344 10792
rect 3513 10755 3571 10761
rect 4338 10752 4344 10764
rect 4396 10752 4402 10804
rect 4522 10752 4528 10804
rect 4580 10792 4586 10804
rect 4709 10795 4767 10801
rect 4709 10792 4721 10795
rect 4580 10764 4721 10792
rect 4580 10752 4586 10764
rect 4709 10761 4721 10764
rect 4755 10761 4767 10795
rect 4709 10755 4767 10761
rect 6086 10752 6092 10804
rect 6144 10792 6150 10804
rect 6457 10795 6515 10801
rect 6457 10792 6469 10795
rect 6144 10764 6469 10792
rect 6144 10752 6150 10764
rect 6457 10761 6469 10764
rect 6503 10761 6515 10795
rect 6457 10755 6515 10761
rect 9950 10752 9956 10804
rect 10008 10792 10014 10804
rect 10321 10795 10379 10801
rect 10321 10792 10333 10795
rect 10008 10764 10333 10792
rect 10008 10752 10014 10764
rect 10321 10761 10333 10764
rect 10367 10761 10379 10795
rect 10321 10755 10379 10761
rect 10686 10752 10692 10804
rect 10744 10792 10750 10804
rect 11977 10795 12035 10801
rect 11977 10792 11989 10795
rect 10744 10764 11989 10792
rect 10744 10752 10750 10764
rect 11977 10761 11989 10764
rect 12023 10761 12035 10795
rect 12526 10792 12532 10804
rect 12487 10764 12532 10792
rect 11977 10755 12035 10761
rect 12526 10752 12532 10764
rect 12584 10752 12590 10804
rect 13265 10795 13323 10801
rect 13265 10761 13277 10795
rect 13311 10792 13323 10795
rect 13354 10792 13360 10804
rect 13311 10764 13360 10792
rect 13311 10761 13323 10764
rect 13265 10755 13323 10761
rect 13354 10752 13360 10764
rect 13412 10752 13418 10804
rect 3881 10727 3939 10733
rect 2746 10696 3188 10724
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 2746 10656 2774 10696
rect 1719 10628 2774 10656
rect 3053 10659 3111 10665
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 3053 10625 3065 10659
rect 3099 10625 3111 10659
rect 3160 10656 3188 10696
rect 3881 10693 3893 10727
rect 3927 10724 3939 10727
rect 4062 10724 4068 10736
rect 3927 10696 4068 10724
rect 3927 10693 3939 10696
rect 3881 10687 3939 10693
rect 4062 10684 4068 10696
rect 4120 10724 4126 10736
rect 5626 10724 5632 10736
rect 4120 10696 5632 10724
rect 4120 10684 4126 10696
rect 5626 10684 5632 10696
rect 5684 10684 5690 10736
rect 5810 10684 5816 10736
rect 5868 10733 5874 10736
rect 5868 10724 5880 10733
rect 11054 10724 11060 10736
rect 5868 10696 5913 10724
rect 7024 10696 11060 10724
rect 5868 10687 5880 10696
rect 5868 10684 5874 10687
rect 7024 10656 7052 10696
rect 11054 10684 11060 10696
rect 11112 10684 11118 10736
rect 12069 10727 12127 10733
rect 12069 10693 12081 10727
rect 12115 10724 12127 10727
rect 12802 10724 12808 10736
rect 12115 10696 12808 10724
rect 12115 10693 12127 10696
rect 12069 10687 12127 10693
rect 12802 10684 12808 10696
rect 12860 10684 12866 10736
rect 13173 10727 13231 10733
rect 13173 10693 13185 10727
rect 13219 10724 13231 10727
rect 14090 10724 14096 10736
rect 13219 10696 14096 10724
rect 13219 10693 13231 10696
rect 13173 10687 13231 10693
rect 14090 10684 14096 10696
rect 14148 10684 14154 10736
rect 3160 10628 7052 10656
rect 3053 10619 3111 10625
rect 2501 10591 2559 10597
rect 2501 10557 2513 10591
rect 2547 10588 2559 10591
rect 2590 10588 2596 10600
rect 2547 10560 2596 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 2590 10548 2596 10560
rect 2648 10548 2654 10600
rect 3068 10588 3096 10619
rect 7098 10616 7104 10668
rect 7156 10656 7162 10668
rect 7558 10656 7564 10668
rect 7616 10665 7622 10668
rect 7156 10628 7564 10656
rect 7156 10616 7162 10628
rect 7558 10616 7564 10628
rect 7616 10656 7628 10665
rect 9208 10659 9266 10665
rect 7616 10628 7661 10656
rect 7616 10619 7628 10628
rect 9208 10625 9220 10659
rect 9254 10656 9266 10659
rect 9674 10656 9680 10668
rect 9254 10628 9680 10656
rect 9254 10625 9266 10628
rect 9208 10619 9266 10625
rect 7616 10616 7622 10619
rect 9674 10616 9680 10628
rect 9732 10656 9738 10668
rect 10042 10656 10048 10668
rect 9732 10628 10048 10656
rect 9732 10616 9738 10628
rect 10042 10616 10048 10628
rect 10100 10616 10106 10668
rect 11900 10628 12434 10656
rect 11900 10600 11928 10628
rect 3142 10588 3148 10600
rect 3068 10560 3148 10588
rect 3142 10548 3148 10560
rect 3200 10548 3206 10600
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10588 3387 10591
rect 3510 10588 3516 10600
rect 3375 10560 3516 10588
rect 3375 10557 3387 10560
rect 3329 10551 3387 10557
rect 3510 10548 3516 10560
rect 3568 10548 3574 10600
rect 3973 10591 4031 10597
rect 3973 10557 3985 10591
rect 4019 10557 4031 10591
rect 4154 10588 4160 10600
rect 4115 10560 4160 10588
rect 3973 10551 4031 10557
rect 3988 10520 4016 10551
rect 4154 10548 4160 10560
rect 4212 10548 4218 10600
rect 4338 10548 4344 10600
rect 4396 10588 4402 10600
rect 4614 10588 4620 10600
rect 4396 10560 4620 10588
rect 4396 10548 4402 10560
rect 4614 10548 4620 10560
rect 4672 10548 4678 10600
rect 6089 10591 6147 10597
rect 6089 10557 6101 10591
rect 6135 10557 6147 10591
rect 6089 10551 6147 10557
rect 7837 10591 7895 10597
rect 7837 10557 7849 10591
rect 7883 10588 7895 10591
rect 8938 10588 8944 10600
rect 7883 10560 8064 10588
rect 8851 10560 8944 10588
rect 7883 10557 7895 10560
rect 7837 10551 7895 10557
rect 4430 10520 4436 10532
rect 3988 10492 4436 10520
rect 4430 10480 4436 10492
rect 4488 10480 4494 10532
rect 1489 10455 1547 10461
rect 1489 10421 1501 10455
rect 1535 10452 1547 10455
rect 1670 10452 1676 10464
rect 1535 10424 1676 10452
rect 1535 10421 1547 10424
rect 1489 10415 1547 10421
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 4525 10455 4583 10461
rect 4525 10421 4537 10455
rect 4571 10452 4583 10455
rect 5902 10452 5908 10464
rect 4571 10424 5908 10452
rect 4571 10421 4583 10424
rect 4525 10415 4583 10421
rect 5902 10412 5908 10424
rect 5960 10452 5966 10464
rect 6104 10452 6132 10551
rect 8036 10464 8064 10560
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 11882 10588 11888 10600
rect 11843 10560 11888 10588
rect 11882 10548 11888 10560
rect 11940 10548 11946 10600
rect 12406 10588 12434 10628
rect 13357 10591 13415 10597
rect 13357 10588 13369 10591
rect 12406 10560 13369 10588
rect 13357 10557 13369 10560
rect 13403 10557 13415 10591
rect 13357 10551 13415 10557
rect 8018 10452 8024 10464
rect 5960 10424 6132 10452
rect 7979 10424 8024 10452
rect 5960 10412 5966 10424
rect 8018 10412 8024 10424
rect 8076 10452 8082 10464
rect 8757 10455 8815 10461
rect 8757 10452 8769 10455
rect 8076 10424 8769 10452
rect 8076 10412 8082 10424
rect 8757 10421 8769 10424
rect 8803 10452 8815 10455
rect 8956 10452 8984 10548
rect 12437 10523 12495 10529
rect 12437 10489 12449 10523
rect 12483 10520 12495 10523
rect 12618 10520 12624 10532
rect 12483 10492 12624 10520
rect 12483 10489 12495 10492
rect 12437 10483 12495 10489
rect 12618 10480 12624 10492
rect 12676 10480 12682 10532
rect 12710 10480 12716 10532
rect 12768 10520 12774 10532
rect 12805 10523 12863 10529
rect 12805 10520 12817 10523
rect 12768 10492 12817 10520
rect 12768 10480 12774 10492
rect 12805 10489 12817 10492
rect 12851 10489 12863 10523
rect 12805 10483 12863 10489
rect 10505 10455 10563 10461
rect 10505 10452 10517 10455
rect 8803 10424 10517 10452
rect 8803 10421 8815 10424
rect 8757 10415 8815 10421
rect 10505 10421 10517 10424
rect 10551 10421 10563 10455
rect 10505 10415 10563 10421
rect 10778 10412 10784 10464
rect 10836 10452 10842 10464
rect 15286 10452 15292 10464
rect 10836 10424 15292 10452
rect 10836 10412 10842 10424
rect 15286 10412 15292 10424
rect 15344 10452 15350 10464
rect 15930 10452 15936 10464
rect 15344 10424 15936 10452
rect 15344 10412 15350 10424
rect 15930 10412 15936 10424
rect 15988 10412 15994 10464
rect 1104 10362 16008 10384
rect 1104 10310 2824 10362
rect 2876 10310 2888 10362
rect 2940 10310 2952 10362
rect 3004 10310 3016 10362
rect 3068 10310 3080 10362
rect 3132 10310 6572 10362
rect 6624 10310 6636 10362
rect 6688 10310 6700 10362
rect 6752 10310 6764 10362
rect 6816 10310 6828 10362
rect 6880 10310 10320 10362
rect 10372 10310 10384 10362
rect 10436 10310 10448 10362
rect 10500 10310 10512 10362
rect 10564 10310 10576 10362
rect 10628 10310 14068 10362
rect 14120 10310 14132 10362
rect 14184 10310 14196 10362
rect 14248 10310 14260 10362
rect 14312 10310 14324 10362
rect 14376 10310 16008 10362
rect 1104 10288 16008 10310
rect 1762 10248 1768 10260
rect 1723 10220 1768 10248
rect 1762 10208 1768 10220
rect 1820 10208 1826 10260
rect 8757 10251 8815 10257
rect 1964 10220 8432 10248
rect 1670 10044 1676 10056
rect 1631 10016 1676 10044
rect 1670 10004 1676 10016
rect 1728 10004 1734 10056
rect 1964 10053 1992 10220
rect 2406 10140 2412 10192
rect 2464 10180 2470 10192
rect 2961 10183 3019 10189
rect 2961 10180 2973 10183
rect 2464 10152 2973 10180
rect 2464 10140 2470 10152
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10013 2007 10047
rect 2608 10044 2636 10152
rect 2961 10149 2973 10152
rect 3007 10149 3019 10183
rect 2961 10143 3019 10149
rect 3510 10140 3516 10192
rect 3568 10180 3574 10192
rect 3881 10183 3939 10189
rect 3881 10180 3893 10183
rect 3568 10152 3893 10180
rect 3568 10140 3574 10152
rect 3881 10149 3893 10152
rect 3927 10149 3939 10183
rect 3881 10143 3939 10149
rect 2685 10115 2743 10121
rect 2685 10081 2697 10115
rect 2731 10112 2743 10115
rect 4246 10112 4252 10124
rect 2731 10084 4252 10112
rect 2731 10081 2743 10084
rect 2685 10075 2743 10081
rect 4246 10072 4252 10084
rect 4304 10072 4310 10124
rect 8404 10112 8432 10220
rect 8757 10217 8769 10251
rect 8803 10248 8815 10251
rect 10778 10248 10784 10260
rect 8803 10220 10784 10248
rect 8803 10217 8815 10220
rect 8757 10211 8815 10217
rect 10778 10208 10784 10220
rect 10836 10208 10842 10260
rect 8404 10084 10272 10112
rect 3510 10044 3516 10056
rect 2608 10016 3516 10044
rect 1949 10007 2007 10013
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4994 10047 5052 10053
rect 4994 10044 5006 10047
rect 4212 10016 5006 10044
rect 4212 10004 4218 10016
rect 4994 10013 5006 10016
rect 5040 10044 5052 10047
rect 5261 10047 5319 10053
rect 5040 10016 5120 10044
rect 5040 10013 5052 10016
rect 4994 10007 5052 10013
rect 1486 9908 1492 9920
rect 1447 9880 1492 9908
rect 1486 9868 1492 9880
rect 1544 9868 1550 9920
rect 1946 9868 1952 9920
rect 2004 9908 2010 9920
rect 2041 9911 2099 9917
rect 2041 9908 2053 9911
rect 2004 9880 2053 9908
rect 2004 9868 2010 9880
rect 2041 9877 2053 9880
rect 2087 9877 2099 9911
rect 2041 9871 2099 9877
rect 2314 9868 2320 9920
rect 2372 9908 2378 9920
rect 2409 9911 2467 9917
rect 2409 9908 2421 9911
rect 2372 9880 2421 9908
rect 2372 9868 2378 9880
rect 2409 9877 2421 9880
rect 2455 9877 2467 9911
rect 2409 9871 2467 9877
rect 2498 9868 2504 9920
rect 2556 9908 2562 9920
rect 5092 9908 5120 10016
rect 5261 10013 5273 10047
rect 5307 10044 5319 10047
rect 5445 10047 5503 10053
rect 5445 10044 5457 10047
rect 5307 10016 5457 10044
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 5445 10013 5457 10016
rect 5491 10044 5503 10047
rect 5629 10047 5687 10053
rect 5629 10044 5641 10047
rect 5491 10016 5641 10044
rect 5491 10013 5503 10016
rect 5445 10007 5503 10013
rect 5629 10013 5641 10016
rect 5675 10044 5687 10047
rect 5813 10047 5871 10053
rect 5813 10044 5825 10047
rect 5675 10016 5825 10044
rect 5675 10013 5687 10016
rect 5629 10007 5687 10013
rect 5813 10013 5825 10016
rect 5859 10044 5871 10047
rect 5902 10044 5908 10056
rect 5859 10016 5908 10044
rect 5859 10013 5871 10016
rect 5813 10007 5871 10013
rect 5902 10004 5908 10016
rect 5960 10004 5966 10056
rect 7018 10047 7076 10053
rect 7018 10013 7030 10047
rect 7064 10044 7076 10047
rect 7190 10044 7196 10056
rect 7064 10016 7196 10044
rect 7064 10013 7076 10016
rect 7018 10007 7076 10013
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 7285 10047 7343 10053
rect 7285 10013 7297 10047
rect 7331 10044 7343 10047
rect 7377 10047 7435 10053
rect 7377 10044 7389 10047
rect 7331 10016 7389 10044
rect 7331 10013 7343 10016
rect 7285 10007 7343 10013
rect 7377 10013 7389 10016
rect 7423 10044 7435 10047
rect 10137 10047 10195 10053
rect 7423 10016 8064 10044
rect 7423 10013 7435 10016
rect 7377 10007 7435 10013
rect 8036 9988 8064 10016
rect 10137 10013 10149 10047
rect 10183 10013 10195 10047
rect 10244 10044 10272 10084
rect 11146 10072 11152 10124
rect 11204 10112 11210 10124
rect 13173 10115 13231 10121
rect 13173 10112 13185 10115
rect 11204 10084 13185 10112
rect 11204 10072 11210 10084
rect 13173 10081 13185 10084
rect 13219 10081 13231 10115
rect 15102 10112 15108 10124
rect 15063 10084 15108 10112
rect 13173 10075 13231 10081
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 15010 10044 15016 10056
rect 10244 10016 12434 10044
rect 14971 10016 15016 10044
rect 10137 10007 10195 10013
rect 7622 9979 7680 9985
rect 7622 9976 7634 9979
rect 7300 9948 7634 9976
rect 7300 9920 7328 9948
rect 7622 9945 7634 9948
rect 7668 9945 7680 9979
rect 7622 9939 7680 9945
rect 8018 9936 8024 9988
rect 8076 9976 8082 9988
rect 9953 9979 10011 9985
rect 9953 9976 9965 9979
rect 8076 9948 9965 9976
rect 8076 9936 8082 9948
rect 9953 9945 9965 9948
rect 9999 9976 10011 9979
rect 10152 9976 10180 10007
rect 9999 9948 10180 9976
rect 10404 9979 10462 9985
rect 9999 9945 10011 9948
rect 9953 9939 10011 9945
rect 10404 9945 10416 9979
rect 10450 9976 10462 9979
rect 12066 9976 12072 9988
rect 10450 9948 12072 9976
rect 10450 9945 10462 9948
rect 10404 9939 10462 9945
rect 12066 9936 12072 9948
rect 12124 9936 12130 9988
rect 5905 9911 5963 9917
rect 5905 9908 5917 9911
rect 2556 9880 2601 9908
rect 5092 9880 5917 9908
rect 2556 9868 2562 9880
rect 5905 9877 5917 9880
rect 5951 9877 5963 9911
rect 5905 9871 5963 9877
rect 7282 9868 7288 9920
rect 7340 9868 7346 9920
rect 11517 9911 11575 9917
rect 11517 9877 11529 9911
rect 11563 9908 11575 9911
rect 11606 9908 11612 9920
rect 11563 9880 11612 9908
rect 11563 9877 11575 9880
rect 11517 9871 11575 9877
rect 11606 9868 11612 9880
rect 11664 9868 11670 9920
rect 12406 9908 12434 10016
rect 15010 10004 15016 10016
rect 15068 10004 15074 10056
rect 15381 10047 15439 10053
rect 15381 10013 15393 10047
rect 15427 10044 15439 10047
rect 16206 10044 16212 10056
rect 15427 10016 16212 10044
rect 15427 10013 15439 10016
rect 15381 10007 15439 10013
rect 16206 10004 16212 10016
rect 16264 10004 16270 10056
rect 12989 9979 13047 9985
rect 12989 9945 13001 9979
rect 13035 9976 13047 9979
rect 14274 9976 14280 9988
rect 13035 9948 14280 9976
rect 13035 9945 13047 9948
rect 12989 9939 13047 9945
rect 14274 9936 14280 9948
rect 14332 9936 14338 9988
rect 14458 9936 14464 9988
rect 14516 9976 14522 9988
rect 14826 9976 14832 9988
rect 14516 9948 14832 9976
rect 14516 9936 14522 9948
rect 14826 9936 14832 9948
rect 14884 9976 14890 9988
rect 14921 9979 14979 9985
rect 14921 9976 14933 9979
rect 14884 9948 14933 9976
rect 14884 9936 14890 9948
rect 14921 9945 14933 9948
rect 14967 9945 14979 9979
rect 14921 9939 14979 9945
rect 12621 9911 12679 9917
rect 12621 9908 12633 9911
rect 12406 9880 12633 9908
rect 12621 9877 12633 9880
rect 12667 9877 12679 9911
rect 12621 9871 12679 9877
rect 13078 9868 13084 9920
rect 13136 9908 13142 9920
rect 14550 9908 14556 9920
rect 13136 9880 13181 9908
rect 14511 9880 14556 9908
rect 13136 9868 13142 9880
rect 14550 9868 14556 9880
rect 14608 9868 14614 9920
rect 15562 9908 15568 9920
rect 15523 9880 15568 9908
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 1104 9818 16008 9840
rect 1104 9766 4698 9818
rect 4750 9766 4762 9818
rect 4814 9766 4826 9818
rect 4878 9766 4890 9818
rect 4942 9766 4954 9818
rect 5006 9766 8446 9818
rect 8498 9766 8510 9818
rect 8562 9766 8574 9818
rect 8626 9766 8638 9818
rect 8690 9766 8702 9818
rect 8754 9766 12194 9818
rect 12246 9766 12258 9818
rect 12310 9766 12322 9818
rect 12374 9766 12386 9818
rect 12438 9766 12450 9818
rect 12502 9766 16008 9818
rect 1104 9744 16008 9766
rect 2317 9707 2375 9713
rect 2317 9673 2329 9707
rect 2363 9704 2375 9707
rect 2498 9704 2504 9716
rect 2363 9676 2504 9704
rect 2363 9673 2375 9676
rect 2317 9667 2375 9673
rect 2498 9664 2504 9676
rect 2556 9664 2562 9716
rect 7190 9664 7196 9716
rect 7248 9704 7254 9716
rect 9585 9707 9643 9713
rect 9585 9704 9597 9707
rect 7248 9676 9597 9704
rect 7248 9664 7254 9676
rect 9585 9673 9597 9676
rect 9631 9704 9643 9707
rect 11146 9704 11152 9716
rect 9631 9676 11152 9704
rect 9631 9673 9643 9676
rect 9585 9667 9643 9673
rect 11146 9664 11152 9676
rect 11204 9664 11210 9716
rect 13078 9664 13084 9716
rect 13136 9704 13142 9716
rect 13173 9707 13231 9713
rect 13173 9704 13185 9707
rect 13136 9676 13185 9704
rect 13136 9664 13142 9676
rect 13173 9673 13185 9676
rect 13219 9673 13231 9707
rect 14274 9704 14280 9716
rect 14235 9676 14280 9704
rect 13173 9667 13231 9673
rect 14274 9664 14280 9676
rect 14332 9664 14338 9716
rect 14550 9664 14556 9716
rect 14608 9704 14614 9716
rect 14737 9707 14795 9713
rect 14737 9704 14749 9707
rect 14608 9676 14749 9704
rect 14608 9664 14614 9676
rect 14737 9673 14749 9676
rect 14783 9673 14795 9707
rect 14737 9667 14795 9673
rect 3878 9596 3884 9648
rect 3936 9636 3942 9648
rect 5362 9639 5420 9645
rect 5362 9636 5374 9639
rect 3936 9608 5374 9636
rect 3936 9596 3942 9608
rect 5362 9605 5374 9608
rect 5408 9605 5420 9639
rect 7592 9639 7650 9645
rect 5362 9599 5420 9605
rect 5460 9608 6040 9636
rect 1670 9568 1676 9580
rect 1631 9540 1676 9568
rect 1670 9528 1676 9540
rect 1728 9528 1734 9580
rect 1946 9568 1952 9580
rect 1907 9540 1952 9568
rect 1946 9528 1952 9540
rect 2004 9528 2010 9580
rect 2406 9528 2412 9580
rect 2464 9568 2470 9580
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 2464 9540 2697 9568
rect 2464 9528 2470 9540
rect 2685 9537 2697 9540
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 3326 9528 3332 9580
rect 3384 9568 3390 9580
rect 3510 9568 3516 9580
rect 3384 9540 3516 9568
rect 3384 9528 3390 9540
rect 3510 9528 3516 9540
rect 3568 9568 3574 9580
rect 3568 9540 4016 9568
rect 3568 9528 3574 9540
rect 2498 9460 2504 9512
rect 2556 9500 2562 9512
rect 2777 9503 2835 9509
rect 2777 9500 2789 9503
rect 2556 9472 2789 9500
rect 2556 9460 2562 9472
rect 2777 9469 2789 9472
rect 2823 9469 2835 9503
rect 2777 9463 2835 9469
rect 2961 9503 3019 9509
rect 2961 9469 2973 9503
rect 3007 9500 3019 9503
rect 3007 9472 3041 9500
rect 3007 9469 3019 9472
rect 2961 9463 3019 9469
rect 1854 9392 1860 9444
rect 1912 9432 1918 9444
rect 2976 9432 3004 9463
rect 3786 9460 3792 9512
rect 3844 9500 3850 9512
rect 3881 9503 3939 9509
rect 3881 9500 3893 9503
rect 3844 9472 3893 9500
rect 3844 9460 3850 9472
rect 3881 9469 3893 9472
rect 3927 9469 3939 9503
rect 3988 9500 4016 9540
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 4157 9571 4215 9577
rect 4157 9568 4169 9571
rect 4120 9540 4169 9568
rect 4120 9528 4126 9540
rect 4157 9537 4169 9540
rect 4203 9537 4215 9571
rect 5460 9568 5488 9608
rect 4157 9531 4215 9537
rect 4264 9540 5488 9568
rect 5629 9571 5687 9577
rect 4264 9500 4292 9540
rect 5629 9537 5641 9571
rect 5675 9568 5687 9571
rect 5902 9568 5908 9580
rect 5675 9540 5908 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 5902 9528 5908 9540
rect 5960 9528 5966 9580
rect 6012 9568 6040 9608
rect 7592 9605 7604 9639
rect 7638 9636 7650 9639
rect 7834 9636 7840 9648
rect 7638 9608 7840 9636
rect 7638 9605 7650 9608
rect 7592 9599 7650 9605
rect 7834 9596 7840 9608
rect 7892 9596 7898 9648
rect 8110 9596 8116 9648
rect 8168 9636 8174 9648
rect 8358 9639 8416 9645
rect 8358 9636 8370 9639
rect 8168 9608 8370 9636
rect 8168 9596 8174 9608
rect 8358 9605 8370 9608
rect 8404 9605 8416 9639
rect 10134 9636 10140 9648
rect 8358 9599 8416 9605
rect 8496 9608 10140 9636
rect 8496 9568 8524 9608
rect 10134 9596 10140 9608
rect 10192 9596 10198 9648
rect 11333 9639 11391 9645
rect 11333 9605 11345 9639
rect 11379 9636 11391 9639
rect 12526 9636 12532 9648
rect 11379 9608 12532 9636
rect 11379 9605 11391 9608
rect 11333 9599 11391 9605
rect 6012 9540 8524 9568
rect 10709 9571 10767 9577
rect 10709 9537 10721 9571
rect 10755 9568 10767 9571
rect 10965 9571 11023 9577
rect 10755 9540 10916 9568
rect 10755 9537 10767 9540
rect 10709 9531 10767 9537
rect 3988 9472 4292 9500
rect 7837 9503 7895 9509
rect 3881 9463 3939 9469
rect 7837 9469 7849 9503
rect 7883 9500 7895 9503
rect 8113 9503 8171 9509
rect 8113 9500 8125 9503
rect 7883 9472 8125 9500
rect 7883 9469 7895 9472
rect 7837 9463 7895 9469
rect 1912 9404 4292 9432
rect 1912 9392 1918 9404
rect 4264 9376 4292 9404
rect 8036 9376 8064 9472
rect 8113 9469 8125 9472
rect 8159 9469 8171 9503
rect 10888 9500 10916 9540
rect 10965 9537 10977 9571
rect 11011 9568 11023 9571
rect 11348 9568 11376 9599
rect 12526 9596 12532 9608
rect 12584 9636 12590 9648
rect 12584 9608 12940 9636
rect 12584 9596 12590 9608
rect 11011 9540 11376 9568
rect 12641 9571 12699 9577
rect 11011 9537 11023 9540
rect 10965 9531 11023 9537
rect 12641 9537 12653 9571
rect 12687 9568 12699 9571
rect 12802 9568 12808 9580
rect 12687 9540 12808 9568
rect 12687 9537 12699 9540
rect 12641 9531 12699 9537
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 12912 9577 12940 9608
rect 15010 9596 15016 9648
rect 15068 9636 15074 9648
rect 15197 9639 15255 9645
rect 15197 9636 15209 9639
rect 15068 9608 15209 9636
rect 15068 9596 15074 9608
rect 15197 9605 15209 9608
rect 15243 9636 15255 9639
rect 15378 9636 15384 9648
rect 15243 9608 15384 9636
rect 15243 9605 15255 9608
rect 15197 9599 15255 9605
rect 15378 9596 15384 9608
rect 15436 9596 15442 9648
rect 12897 9571 12955 9577
rect 12897 9537 12909 9571
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 13814 9568 13820 9580
rect 13587 9540 13820 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 13814 9528 13820 9540
rect 13872 9528 13878 9580
rect 14645 9571 14703 9577
rect 14645 9537 14657 9571
rect 14691 9568 14703 9571
rect 14918 9568 14924 9580
rect 14691 9540 14924 9568
rect 14691 9537 14703 9540
rect 14645 9531 14703 9537
rect 14918 9528 14924 9540
rect 14976 9528 14982 9580
rect 13630 9500 13636 9512
rect 10888 9472 11560 9500
rect 13591 9472 13636 9500
rect 8113 9463 8171 9469
rect 11532 9441 11560 9472
rect 13630 9460 13636 9472
rect 13688 9460 13694 9512
rect 13725 9503 13783 9509
rect 13725 9469 13737 9503
rect 13771 9500 13783 9503
rect 14829 9503 14887 9509
rect 14829 9500 14841 9503
rect 13771 9472 14841 9500
rect 13771 9469 13783 9472
rect 13725 9463 13783 9469
rect 14829 9469 14841 9472
rect 14875 9469 14887 9503
rect 15286 9500 15292 9512
rect 15247 9472 15292 9500
rect 14829 9463 14887 9469
rect 11517 9435 11575 9441
rect 11517 9401 11529 9435
rect 11563 9401 11575 9435
rect 11517 9395 11575 9401
rect 1486 9364 1492 9376
rect 1447 9336 1492 9364
rect 1486 9324 1492 9336
rect 1544 9324 1550 9376
rect 1762 9364 1768 9376
rect 1723 9336 1768 9364
rect 1762 9324 1768 9336
rect 1820 9324 1826 9376
rect 4246 9364 4252 9376
rect 4207 9336 4252 9364
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 5813 9367 5871 9373
rect 5813 9333 5825 9367
rect 5859 9364 5871 9367
rect 5902 9364 5908 9376
rect 5859 9336 5908 9364
rect 5859 9333 5871 9336
rect 5813 9327 5871 9333
rect 5902 9324 5908 9336
rect 5960 9364 5966 9376
rect 6089 9367 6147 9373
rect 6089 9364 6101 9367
rect 5960 9336 6101 9364
rect 5960 9324 5966 9336
rect 6089 9333 6101 9336
rect 6135 9333 6147 9367
rect 6089 9327 6147 9333
rect 6457 9367 6515 9373
rect 6457 9333 6469 9367
rect 6503 9364 6515 9367
rect 7558 9364 7564 9376
rect 6503 9336 7564 9364
rect 6503 9333 6515 9336
rect 6457 9327 6515 9333
rect 7558 9324 7564 9336
rect 7616 9324 7622 9376
rect 8018 9364 8024 9376
rect 7979 9336 8024 9364
rect 8018 9324 8024 9336
rect 8076 9324 8082 9376
rect 9493 9367 9551 9373
rect 9493 9333 9505 9367
rect 9539 9364 9551 9367
rect 9582 9364 9588 9376
rect 9539 9336 9588 9364
rect 9539 9333 9551 9336
rect 9493 9327 9551 9333
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 11532 9364 11560 9395
rect 13740 9364 13768 9463
rect 15286 9460 15292 9472
rect 15344 9460 15350 9512
rect 11532 9336 13768 9364
rect 1104 9274 16008 9296
rect 1104 9222 2824 9274
rect 2876 9222 2888 9274
rect 2940 9222 2952 9274
rect 3004 9222 3016 9274
rect 3068 9222 3080 9274
rect 3132 9222 6572 9274
rect 6624 9222 6636 9274
rect 6688 9222 6700 9274
rect 6752 9222 6764 9274
rect 6816 9222 6828 9274
rect 6880 9222 10320 9274
rect 10372 9222 10384 9274
rect 10436 9222 10448 9274
rect 10500 9222 10512 9274
rect 10564 9222 10576 9274
rect 10628 9222 14068 9274
rect 14120 9222 14132 9274
rect 14184 9222 14196 9274
rect 14248 9222 14260 9274
rect 14312 9222 14324 9274
rect 14376 9222 16008 9274
rect 1104 9200 16008 9222
rect 2406 9160 2412 9172
rect 2367 9132 2412 9160
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 2590 9120 2596 9172
rect 2648 9160 2654 9172
rect 9766 9160 9772 9172
rect 2648 9132 9772 9160
rect 2648 9120 2654 9132
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 10042 9160 10048 9172
rect 10003 9132 10048 9160
rect 10042 9120 10048 9132
rect 10100 9120 10106 9172
rect 13630 9120 13636 9172
rect 13688 9160 13694 9172
rect 14093 9163 14151 9169
rect 14093 9160 14105 9163
rect 13688 9132 14105 9160
rect 13688 9120 13694 9132
rect 14093 9129 14105 9132
rect 14139 9129 14151 9163
rect 14918 9160 14924 9172
rect 14879 9132 14924 9160
rect 14093 9123 14151 9129
rect 14918 9120 14924 9132
rect 14976 9120 14982 9172
rect 3878 9092 3884 9104
rect 1872 9064 3884 9092
rect 1872 9033 1900 9064
rect 3878 9052 3884 9064
rect 3936 9052 3942 9104
rect 12802 9052 12808 9104
rect 12860 9092 12866 9104
rect 12897 9095 12955 9101
rect 12897 9092 12909 9095
rect 12860 9064 12909 9092
rect 12860 9052 12866 9064
rect 12897 9061 12909 9064
rect 12943 9092 12955 9095
rect 13906 9092 13912 9104
rect 12943 9064 13912 9092
rect 12943 9061 12955 9064
rect 12897 9055 12955 9061
rect 13906 9052 13912 9064
rect 13964 9092 13970 9104
rect 13964 9064 14780 9092
rect 13964 9052 13970 9064
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 8993 1915 9027
rect 3329 9027 3387 9033
rect 3329 9024 3341 9027
rect 1857 8987 1915 8993
rect 2746 8996 3341 9024
rect 2746 8968 2774 8996
rect 3329 8993 3341 8996
rect 3375 8993 3387 9027
rect 3510 9024 3516 9036
rect 3471 8996 3516 9024
rect 3329 8987 3387 8993
rect 3510 8984 3516 8996
rect 3568 8984 3574 9036
rect 14752 9033 14780 9064
rect 13081 9027 13139 9033
rect 13081 8993 13093 9027
rect 13127 8993 13139 9027
rect 13081 8987 13139 8993
rect 14737 9027 14795 9033
rect 14737 8993 14749 9027
rect 14783 9024 14795 9027
rect 15102 9024 15108 9036
rect 14783 8996 15108 9024
rect 14783 8993 14795 8996
rect 14737 8987 14795 8993
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8956 2007 8959
rect 2682 8956 2688 8968
rect 1995 8928 2688 8956
rect 1995 8925 2007 8928
rect 1949 8919 2007 8925
rect 2682 8916 2688 8928
rect 2740 8928 2774 8968
rect 3053 8959 3111 8965
rect 2740 8916 2746 8928
rect 3053 8925 3065 8959
rect 3099 8956 3111 8959
rect 3694 8956 3700 8968
rect 3099 8928 3700 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 3694 8916 3700 8928
rect 3752 8916 3758 8968
rect 4433 8959 4491 8965
rect 4433 8925 4445 8959
rect 4479 8956 4491 8959
rect 5902 8956 5908 8968
rect 4479 8928 5908 8956
rect 4479 8925 4491 8928
rect 4433 8919 4491 8925
rect 5902 8916 5908 8928
rect 5960 8916 5966 8968
rect 11425 8959 11483 8965
rect 11425 8956 11437 8959
rect 9876 8928 11437 8956
rect 2041 8891 2099 8897
rect 2041 8857 2053 8891
rect 2087 8888 2099 8891
rect 2087 8860 2774 8888
rect 2087 8857 2099 8860
rect 2041 8851 2099 8857
rect 2746 8820 2774 8860
rect 2866 8848 2872 8900
rect 2924 8888 2930 8900
rect 3142 8888 3148 8900
rect 2924 8860 3148 8888
rect 2924 8848 2930 8860
rect 3142 8848 3148 8860
rect 3200 8888 3206 8900
rect 3200 8860 3464 8888
rect 3200 8848 3206 8860
rect 3326 8820 3332 8832
rect 2746 8792 3332 8820
rect 3326 8780 3332 8792
rect 3384 8780 3390 8832
rect 3436 8820 3464 8860
rect 4338 8848 4344 8900
rect 4396 8888 4402 8900
rect 4678 8891 4736 8897
rect 4678 8888 4690 8891
rect 4396 8860 4690 8888
rect 4396 8848 4402 8860
rect 4678 8857 4690 8860
rect 4724 8857 4736 8891
rect 6150 8891 6208 8897
rect 6150 8888 6162 8891
rect 4678 8851 4736 8857
rect 5828 8860 6162 8888
rect 4522 8820 4528 8832
rect 3436 8792 4528 8820
rect 4522 8780 4528 8792
rect 4580 8780 4586 8832
rect 5718 8780 5724 8832
rect 5776 8820 5782 8832
rect 5828 8829 5856 8860
rect 6150 8857 6162 8860
rect 6196 8857 6208 8891
rect 6150 8851 6208 8857
rect 5813 8823 5871 8829
rect 5813 8820 5825 8823
rect 5776 8792 5825 8820
rect 5776 8780 5782 8792
rect 5813 8789 5825 8792
rect 5859 8789 5871 8823
rect 5813 8783 5871 8789
rect 7285 8823 7343 8829
rect 7285 8789 7297 8823
rect 7331 8820 7343 8823
rect 7926 8820 7932 8832
rect 7331 8792 7932 8820
rect 7331 8789 7343 8792
rect 7285 8783 7343 8789
rect 7926 8780 7932 8792
rect 7984 8780 7990 8832
rect 8018 8780 8024 8832
rect 8076 8820 8082 8832
rect 8846 8820 8852 8832
rect 8076 8792 8852 8820
rect 8076 8780 8082 8792
rect 8846 8780 8852 8792
rect 8904 8820 8910 8832
rect 9876 8829 9904 8928
rect 11425 8925 11437 8928
rect 11471 8956 11483 8959
rect 11517 8959 11575 8965
rect 11517 8956 11529 8959
rect 11471 8928 11529 8956
rect 11471 8925 11483 8928
rect 11425 8919 11483 8925
rect 11517 8925 11529 8928
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 11606 8916 11612 8968
rect 11664 8956 11670 8968
rect 11773 8959 11831 8965
rect 11773 8956 11785 8959
rect 11664 8928 11785 8956
rect 11664 8916 11670 8928
rect 11773 8925 11785 8928
rect 11819 8956 11831 8959
rect 13096 8956 13124 8987
rect 15102 8984 15108 8996
rect 15160 9024 15166 9036
rect 15473 9027 15531 9033
rect 15473 9024 15485 9027
rect 15160 8996 15485 9024
rect 15160 8984 15166 8996
rect 15473 8993 15485 8996
rect 15519 8993 15531 9027
rect 15473 8987 15531 8993
rect 14918 8956 14924 8968
rect 11819 8928 14924 8956
rect 11819 8925 11831 8928
rect 11773 8919 11831 8925
rect 14918 8916 14924 8928
rect 14976 8916 14982 8968
rect 15286 8956 15292 8968
rect 15247 8928 15292 8956
rect 15286 8916 15292 8928
rect 15344 8916 15350 8968
rect 15378 8916 15384 8968
rect 15436 8956 15442 8968
rect 15436 8928 15481 8956
rect 15436 8916 15442 8928
rect 11180 8891 11238 8897
rect 11180 8857 11192 8891
rect 11226 8888 11238 8891
rect 11882 8888 11888 8900
rect 11226 8860 11888 8888
rect 11226 8857 11238 8860
rect 11180 8851 11238 8857
rect 11882 8848 11888 8860
rect 11940 8848 11946 8900
rect 12710 8848 12716 8900
rect 12768 8888 12774 8900
rect 13357 8891 13415 8897
rect 13357 8888 13369 8891
rect 12768 8860 13369 8888
rect 12768 8848 12774 8860
rect 13357 8857 13369 8860
rect 13403 8857 13415 8891
rect 13357 8851 13415 8857
rect 9401 8823 9459 8829
rect 9401 8820 9413 8823
rect 8904 8792 9413 8820
rect 8904 8780 8910 8792
rect 9401 8789 9413 8792
rect 9447 8820 9459 8823
rect 9861 8823 9919 8829
rect 9861 8820 9873 8823
rect 9447 8792 9873 8820
rect 9447 8789 9459 8792
rect 9401 8783 9459 8789
rect 9861 8789 9873 8792
rect 9907 8789 9919 8823
rect 9861 8783 9919 8789
rect 13170 8780 13176 8832
rect 13228 8820 13234 8832
rect 13265 8823 13323 8829
rect 13265 8820 13277 8823
rect 13228 8792 13277 8820
rect 13228 8780 13234 8792
rect 13265 8789 13277 8792
rect 13311 8789 13323 8823
rect 13722 8820 13728 8832
rect 13683 8792 13728 8820
rect 13265 8783 13323 8789
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 14458 8820 14464 8832
rect 14419 8792 14464 8820
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 14550 8780 14556 8832
rect 14608 8820 14614 8832
rect 14608 8792 14653 8820
rect 14608 8780 14614 8792
rect 1104 8730 16008 8752
rect 1104 8678 4698 8730
rect 4750 8678 4762 8730
rect 4814 8678 4826 8730
rect 4878 8678 4890 8730
rect 4942 8678 4954 8730
rect 5006 8678 8446 8730
rect 8498 8678 8510 8730
rect 8562 8678 8574 8730
rect 8626 8678 8638 8730
rect 8690 8678 8702 8730
rect 8754 8678 12194 8730
rect 12246 8678 12258 8730
rect 12310 8678 12322 8730
rect 12374 8678 12386 8730
rect 12438 8678 12450 8730
rect 12502 8678 16008 8730
rect 1104 8656 16008 8678
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 2409 8619 2467 8625
rect 2409 8616 2421 8619
rect 2372 8588 2421 8616
rect 2372 8576 2378 8588
rect 2409 8585 2421 8588
rect 2455 8585 2467 8619
rect 2409 8579 2467 8585
rect 2498 8576 2504 8628
rect 2556 8616 2562 8628
rect 2866 8616 2872 8628
rect 2556 8588 2601 8616
rect 2827 8588 2872 8616
rect 2556 8576 2562 8588
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 2961 8619 3019 8625
rect 2961 8585 2973 8619
rect 3007 8616 3019 8619
rect 3329 8619 3387 8625
rect 3329 8616 3341 8619
rect 3007 8588 3341 8616
rect 3007 8585 3019 8588
rect 2961 8579 3019 8585
rect 3329 8585 3341 8588
rect 3375 8585 3387 8619
rect 3329 8579 3387 8585
rect 3697 8619 3755 8625
rect 3697 8585 3709 8619
rect 3743 8616 3755 8619
rect 4062 8616 4068 8628
rect 3743 8588 4068 8616
rect 3743 8585 3755 8588
rect 3697 8579 3755 8585
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 4338 8576 4344 8628
rect 4396 8616 4402 8628
rect 5537 8619 5595 8625
rect 5537 8616 5549 8619
rect 4396 8588 5549 8616
rect 4396 8576 4402 8588
rect 5537 8585 5549 8588
rect 5583 8585 5595 8619
rect 5537 8579 5595 8585
rect 5813 8619 5871 8625
rect 5813 8585 5825 8619
rect 5859 8616 5871 8619
rect 5902 8616 5908 8628
rect 5859 8588 5908 8616
rect 5859 8585 5871 8588
rect 5813 8579 5871 8585
rect 1949 8551 2007 8557
rect 1949 8517 1961 8551
rect 1995 8548 2007 8551
rect 3142 8548 3148 8560
rect 1995 8520 3148 8548
rect 1995 8517 2007 8520
rect 1949 8511 2007 8517
rect 3142 8508 3148 8520
rect 3200 8508 3206 8560
rect 3234 8508 3240 8560
rect 3292 8548 3298 8560
rect 3510 8548 3516 8560
rect 3292 8520 3516 8548
rect 3292 8508 3298 8520
rect 3510 8508 3516 8520
rect 3568 8508 3574 8560
rect 5828 8548 5856 8579
rect 5902 8576 5908 8588
rect 5960 8616 5966 8628
rect 5997 8619 6055 8625
rect 5997 8616 6009 8619
rect 5960 8588 6009 8616
rect 5960 8576 5966 8588
rect 5997 8585 6009 8588
rect 6043 8616 6055 8619
rect 6181 8619 6239 8625
rect 6181 8616 6193 8619
rect 6043 8588 6193 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 6181 8585 6193 8588
rect 6227 8616 6239 8619
rect 7193 8619 7251 8625
rect 7193 8616 7205 8619
rect 6227 8588 7205 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 7193 8585 7205 8588
rect 7239 8616 7251 8619
rect 7377 8619 7435 8625
rect 7377 8616 7389 8619
rect 7239 8588 7389 8616
rect 7239 8585 7251 8588
rect 7193 8579 7251 8585
rect 7377 8585 7389 8588
rect 7423 8616 7435 8619
rect 8018 8616 8024 8628
rect 7423 8588 8024 8616
rect 7423 8585 7435 8588
rect 7377 8579 7435 8585
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 13357 8619 13415 8625
rect 13357 8585 13369 8619
rect 13403 8616 13415 8619
rect 13722 8616 13728 8628
rect 13403 8588 13728 8616
rect 13403 8585 13415 8588
rect 13357 8579 13415 8585
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 13814 8576 13820 8628
rect 13872 8616 13878 8628
rect 14369 8619 14427 8625
rect 13872 8588 13917 8616
rect 13872 8576 13878 8588
rect 14369 8585 14381 8619
rect 14415 8616 14427 8619
rect 14550 8616 14556 8628
rect 14415 8588 14556 8616
rect 14415 8585 14427 8588
rect 14369 8579 14427 8585
rect 14550 8576 14556 8588
rect 14608 8576 14614 8628
rect 14642 8576 14648 8628
rect 14700 8616 14706 8628
rect 14737 8619 14795 8625
rect 14737 8616 14749 8619
rect 14700 8588 14749 8616
rect 14700 8576 14706 8588
rect 14737 8585 14749 8588
rect 14783 8585 14795 8619
rect 15378 8616 15384 8628
rect 15339 8588 15384 8616
rect 14737 8579 14795 8585
rect 4172 8520 5856 8548
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8480 2099 8483
rect 3878 8480 3884 8492
rect 2087 8452 2774 8480
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 1854 8412 1860 8424
rect 1815 8384 1860 8412
rect 1854 8372 1860 8384
rect 1912 8372 1918 8424
rect 2746 8344 2774 8452
rect 3160 8452 3884 8480
rect 3160 8421 3188 8452
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 4172 8489 4200 8520
rect 6270 8508 6276 8560
rect 6328 8548 6334 8560
rect 9186 8551 9244 8557
rect 9186 8548 9198 8551
rect 6328 8520 9198 8548
rect 6328 8508 6334 8520
rect 9186 8517 9198 8520
rect 9232 8517 9244 8551
rect 9186 8511 9244 8517
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8449 4215 8483
rect 4157 8443 4215 8449
rect 4246 8440 4252 8492
rect 4304 8480 4310 8492
rect 4413 8483 4471 8489
rect 4413 8480 4425 8483
rect 4304 8452 4425 8480
rect 4304 8440 4310 8452
rect 4413 8449 4425 8452
rect 4459 8449 4471 8483
rect 4413 8443 4471 8449
rect 7374 8440 7380 8492
rect 7432 8480 7438 8492
rect 8582 8483 8640 8489
rect 8582 8480 8594 8483
rect 7432 8452 8594 8480
rect 7432 8440 7438 8452
rect 8582 8449 8594 8452
rect 8628 8449 8640 8483
rect 8582 8443 8640 8449
rect 13449 8483 13507 8489
rect 13449 8449 13461 8483
rect 13495 8480 13507 8483
rect 13538 8480 13544 8492
rect 13495 8452 13544 8480
rect 13495 8449 13507 8452
rect 13449 8443 13507 8449
rect 13538 8440 13544 8452
rect 13596 8480 13602 8492
rect 14642 8480 14648 8492
rect 13596 8452 14648 8480
rect 13596 8440 13602 8452
rect 14642 8440 14648 8452
rect 14700 8440 14706 8492
rect 3145 8415 3203 8421
rect 3145 8381 3157 8415
rect 3191 8381 3203 8415
rect 3145 8375 3203 8381
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8381 3847 8415
rect 3789 8375 3847 8381
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8412 4031 8415
rect 8846 8412 8852 8424
rect 4019 8384 4200 8412
rect 8807 8384 8852 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 3234 8344 3240 8356
rect 2746 8316 3240 8344
rect 3234 8304 3240 8316
rect 3292 8304 3298 8356
rect 3804 8344 3832 8375
rect 4062 8344 4068 8356
rect 3804 8316 4068 8344
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 4172 8276 4200 8384
rect 8846 8372 8852 8384
rect 8904 8412 8910 8424
rect 8941 8415 8999 8421
rect 8941 8412 8953 8415
rect 8904 8384 8953 8412
rect 8904 8372 8910 8384
rect 8941 8381 8953 8384
rect 8987 8381 8999 8415
rect 8941 8375 8999 8381
rect 13265 8415 13323 8421
rect 13265 8381 13277 8415
rect 13311 8412 13323 8415
rect 13906 8412 13912 8424
rect 13311 8384 13912 8412
rect 13311 8381 13323 8384
rect 13265 8375 13323 8381
rect 13906 8372 13912 8384
rect 13964 8372 13970 8424
rect 14550 8372 14556 8424
rect 14608 8412 14614 8424
rect 14752 8412 14780 8579
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 14829 8551 14887 8557
rect 14829 8517 14841 8551
rect 14875 8548 14887 8551
rect 15470 8548 15476 8560
rect 14875 8520 15476 8548
rect 14875 8517 14887 8520
rect 14829 8511 14887 8517
rect 15470 8508 15476 8520
rect 15528 8508 15534 8560
rect 14608 8384 14780 8412
rect 14608 8372 14614 8384
rect 14918 8372 14924 8424
rect 14976 8412 14982 8424
rect 14976 8384 15021 8412
rect 14976 8372 14982 8384
rect 7466 8344 7472 8356
rect 7427 8316 7472 8344
rect 7466 8304 7472 8316
rect 7524 8304 7530 8356
rect 10321 8347 10379 8353
rect 10321 8313 10333 8347
rect 10367 8344 10379 8347
rect 11606 8344 11612 8356
rect 10367 8316 11612 8344
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 11606 8304 11612 8316
rect 11664 8304 11670 8356
rect 12897 8347 12955 8353
rect 12897 8313 12909 8347
rect 12943 8344 12955 8347
rect 13170 8344 13176 8356
rect 12943 8316 13176 8344
rect 12943 8313 12955 8316
rect 12897 8307 12955 8313
rect 13170 8304 13176 8316
rect 13228 8344 13234 8356
rect 13814 8344 13820 8356
rect 13228 8316 13820 8344
rect 13228 8304 13234 8316
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 15194 8304 15200 8356
rect 15252 8344 15258 8356
rect 15473 8347 15531 8353
rect 15473 8344 15485 8347
rect 15252 8316 15485 8344
rect 15252 8304 15258 8316
rect 15473 8313 15485 8316
rect 15519 8313 15531 8347
rect 15473 8307 15531 8313
rect 5166 8276 5172 8288
rect 4172 8248 5172 8276
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 10689 8279 10747 8285
rect 10689 8245 10701 8279
rect 10735 8276 10747 8279
rect 10778 8276 10784 8288
rect 10735 8248 10784 8276
rect 10735 8245 10747 8248
rect 10689 8239 10747 8245
rect 10778 8236 10784 8248
rect 10836 8276 10842 8288
rect 11517 8279 11575 8285
rect 11517 8276 11529 8279
rect 10836 8248 11529 8276
rect 10836 8236 10842 8248
rect 11517 8245 11529 8248
rect 11563 8276 11575 8279
rect 12069 8279 12127 8285
rect 12069 8276 12081 8279
rect 11563 8248 12081 8276
rect 11563 8245 11575 8248
rect 11517 8239 11575 8245
rect 12069 8245 12081 8248
rect 12115 8245 12127 8279
rect 12710 8276 12716 8288
rect 12671 8248 12716 8276
rect 12069 8239 12127 8245
rect 12710 8236 12716 8248
rect 12768 8236 12774 8288
rect 12986 8236 12992 8288
rect 13044 8276 13050 8288
rect 14550 8276 14556 8288
rect 13044 8248 14556 8276
rect 13044 8236 13050 8248
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 1104 8186 16008 8208
rect 1104 8134 2824 8186
rect 2876 8134 2888 8186
rect 2940 8134 2952 8186
rect 3004 8134 3016 8186
rect 3068 8134 3080 8186
rect 3132 8134 6572 8186
rect 6624 8134 6636 8186
rect 6688 8134 6700 8186
rect 6752 8134 6764 8186
rect 6816 8134 6828 8186
rect 6880 8134 10320 8186
rect 10372 8134 10384 8186
rect 10436 8134 10448 8186
rect 10500 8134 10512 8186
rect 10564 8134 10576 8186
rect 10628 8134 14068 8186
rect 14120 8134 14132 8186
rect 14184 8134 14196 8186
rect 14248 8134 14260 8186
rect 14312 8134 14324 8186
rect 14376 8134 16008 8186
rect 1104 8112 16008 8134
rect 1486 8072 1492 8084
rect 1447 8044 1492 8072
rect 1486 8032 1492 8044
rect 1544 8032 1550 8084
rect 2869 8075 2927 8081
rect 2869 8041 2881 8075
rect 2915 8072 2927 8075
rect 3142 8072 3148 8084
rect 2915 8044 3148 8072
rect 2915 8041 2927 8044
rect 2869 8035 2927 8041
rect 3142 8032 3148 8044
rect 3200 8032 3206 8084
rect 3878 8072 3884 8084
rect 3839 8044 3884 8072
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 11882 8032 11888 8084
rect 11940 8072 11946 8084
rect 12253 8075 12311 8081
rect 12253 8072 12265 8075
rect 11940 8044 12265 8072
rect 11940 8032 11946 8044
rect 12253 8041 12265 8044
rect 12299 8072 12311 8075
rect 12894 8072 12900 8084
rect 12299 8044 12900 8072
rect 12299 8041 12311 8044
rect 12253 8035 12311 8041
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 13446 8032 13452 8084
rect 13504 8072 13510 8084
rect 14458 8072 14464 8084
rect 13504 8044 13952 8072
rect 14419 8044 14464 8072
rect 13504 8032 13510 8044
rect 1765 8007 1823 8013
rect 1765 7973 1777 8007
rect 1811 7973 1823 8007
rect 1765 7967 1823 7973
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 1780 7868 1808 7967
rect 3418 7896 3424 7948
rect 3476 7936 3482 7948
rect 3513 7939 3571 7945
rect 3513 7936 3525 7939
rect 3476 7908 3525 7936
rect 3476 7896 3482 7908
rect 3513 7905 3525 7908
rect 3559 7936 3571 7939
rect 3896 7936 3924 8032
rect 12161 8007 12219 8013
rect 12161 7973 12173 8007
rect 12207 8004 12219 8007
rect 12618 8004 12624 8016
rect 12207 7976 12624 8004
rect 12207 7973 12219 7976
rect 12161 7967 12219 7973
rect 12618 7964 12624 7976
rect 12676 7964 12682 8016
rect 3559 7908 3924 7936
rect 10520 7908 10916 7936
rect 3559 7905 3571 7908
rect 3513 7899 3571 7905
rect 1719 7840 1808 7868
rect 1949 7871 2007 7877
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 1949 7837 1961 7871
rect 1995 7868 2007 7871
rect 4430 7868 4436 7880
rect 1995 7840 4436 7868
rect 1995 7837 2007 7840
rect 1949 7831 2007 7837
rect 4430 7828 4436 7840
rect 4488 7828 4494 7880
rect 5005 7871 5063 7877
rect 5005 7837 5017 7871
rect 5051 7868 5063 7871
rect 5166 7868 5172 7880
rect 5051 7840 5172 7868
rect 5051 7837 5063 7840
rect 5005 7831 5063 7837
rect 5166 7828 5172 7840
rect 5224 7828 5230 7880
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5445 7871 5503 7877
rect 5445 7868 5457 7871
rect 5307 7840 5457 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5445 7837 5457 7840
rect 5491 7868 5503 7871
rect 6917 7871 6975 7877
rect 6917 7868 6929 7871
rect 5491 7840 6929 7868
rect 5491 7837 5503 7840
rect 5445 7831 5503 7837
rect 6917 7837 6929 7840
rect 6963 7868 6975 7871
rect 7193 7871 7251 7877
rect 7193 7868 7205 7871
rect 6963 7840 7205 7868
rect 6963 7837 6975 7840
rect 6917 7831 6975 7837
rect 7193 7837 7205 7840
rect 7239 7868 7251 7871
rect 8665 7871 8723 7877
rect 8665 7868 8677 7871
rect 7239 7840 8677 7868
rect 7239 7837 7251 7840
rect 7193 7831 7251 7837
rect 8665 7837 8677 7840
rect 8711 7868 8723 7871
rect 8846 7868 8852 7880
rect 8711 7840 8852 7868
rect 8711 7837 8723 7840
rect 8665 7831 8723 7837
rect 8846 7828 8852 7840
rect 8904 7868 8910 7880
rect 9033 7871 9091 7877
rect 9033 7868 9045 7871
rect 8904 7840 9045 7868
rect 8904 7828 8910 7840
rect 9033 7837 9045 7840
rect 9079 7868 9091 7871
rect 9217 7871 9275 7877
rect 9217 7868 9229 7871
rect 9079 7840 9229 7868
rect 9079 7837 9091 7840
rect 9033 7831 9091 7837
rect 9217 7837 9229 7840
rect 9263 7868 9275 7871
rect 9309 7871 9367 7877
rect 9309 7868 9321 7871
rect 9263 7840 9321 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 9309 7837 9321 7840
rect 9355 7868 9367 7871
rect 9398 7868 9404 7880
rect 9355 7840 9404 7868
rect 9355 7837 9367 7840
rect 9309 7831 9367 7837
rect 9398 7828 9404 7840
rect 9456 7828 9462 7880
rect 2777 7803 2835 7809
rect 2777 7769 2789 7803
rect 2823 7800 2835 7803
rect 3142 7800 3148 7812
rect 2823 7772 3148 7800
rect 2823 7769 2835 7772
rect 2777 7763 2835 7769
rect 3142 7760 3148 7772
rect 3200 7760 3206 7812
rect 3329 7803 3387 7809
rect 3329 7769 3341 7803
rect 3375 7800 3387 7803
rect 3970 7800 3976 7812
rect 3375 7772 3976 7800
rect 3375 7769 3387 7772
rect 3329 7763 3387 7769
rect 3970 7760 3976 7772
rect 4028 7760 4034 7812
rect 4062 7760 4068 7812
rect 4120 7800 4126 7812
rect 6672 7803 6730 7809
rect 6672 7800 6684 7803
rect 4120 7772 6684 7800
rect 4120 7760 4126 7772
rect 6672 7769 6684 7772
rect 6718 7800 6730 7803
rect 6718 7772 7328 7800
rect 6718 7769 6730 7772
rect 6672 7763 6730 7769
rect 3237 7735 3295 7741
rect 3237 7701 3249 7735
rect 3283 7732 3295 7735
rect 3602 7732 3608 7744
rect 3283 7704 3608 7732
rect 3283 7701 3295 7704
rect 3237 7695 3295 7701
rect 3602 7692 3608 7704
rect 3660 7692 3666 7744
rect 5442 7692 5448 7744
rect 5500 7732 5506 7744
rect 7300 7741 7328 7772
rect 7926 7760 7932 7812
rect 7984 7800 7990 7812
rect 9582 7809 9588 7812
rect 8398 7803 8456 7809
rect 8398 7800 8410 7803
rect 7984 7772 8410 7800
rect 7984 7760 7990 7772
rect 8398 7769 8410 7772
rect 8444 7769 8456 7803
rect 9576 7800 9588 7809
rect 9495 7772 9588 7800
rect 8398 7763 8456 7769
rect 9576 7763 9588 7772
rect 9640 7800 9646 7812
rect 10520 7800 10548 7908
rect 10778 7868 10784 7880
rect 10739 7840 10784 7868
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 10888 7868 10916 7908
rect 13924 7880 13952 8044
rect 14458 8032 14464 8044
rect 14516 8032 14522 8084
rect 14918 7896 14924 7948
rect 14976 7936 14982 7948
rect 15013 7939 15071 7945
rect 15013 7936 15025 7939
rect 14976 7908 15025 7936
rect 14976 7896 14982 7908
rect 15013 7905 15025 7908
rect 15059 7905 15071 7939
rect 15013 7899 15071 7905
rect 13630 7868 13636 7880
rect 10888 7840 13492 7868
rect 13591 7840 13636 7868
rect 11048 7803 11106 7809
rect 11048 7800 11060 7803
rect 9640 7772 10548 7800
rect 10704 7772 11060 7800
rect 9582 7760 9588 7763
rect 9640 7760 9646 7772
rect 10704 7741 10732 7772
rect 11048 7769 11060 7772
rect 11094 7800 11106 7803
rect 11094 7772 12434 7800
rect 11094 7769 11106 7772
rect 11048 7763 11106 7769
rect 5537 7735 5595 7741
rect 5537 7732 5549 7735
rect 5500 7704 5549 7732
rect 5500 7692 5506 7704
rect 5537 7701 5549 7704
rect 5583 7701 5595 7735
rect 5537 7695 5595 7701
rect 7285 7735 7343 7741
rect 7285 7701 7297 7735
rect 7331 7701 7343 7735
rect 7285 7695 7343 7701
rect 10689 7735 10747 7741
rect 10689 7701 10701 7735
rect 10735 7701 10747 7735
rect 12406 7732 12434 7772
rect 12618 7760 12624 7812
rect 12676 7800 12682 7812
rect 13078 7800 13084 7812
rect 12676 7772 13084 7800
rect 12676 7760 12682 7772
rect 13078 7760 13084 7772
rect 13136 7800 13142 7812
rect 13366 7803 13424 7809
rect 13366 7800 13378 7803
rect 13136 7772 13378 7800
rect 13136 7760 13142 7772
rect 13366 7769 13378 7772
rect 13412 7769 13424 7803
rect 13464 7800 13492 7840
rect 13630 7828 13636 7840
rect 13688 7828 13694 7880
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 13964 7840 14964 7868
rect 13964 7828 13970 7840
rect 14366 7800 14372 7812
rect 13464 7772 14372 7800
rect 13366 7763 13424 7769
rect 14366 7760 14372 7772
rect 14424 7760 14430 7812
rect 14936 7809 14964 7840
rect 14921 7803 14979 7809
rect 14921 7769 14933 7803
rect 14967 7769 14979 7803
rect 14921 7763 14979 7769
rect 13446 7732 13452 7744
rect 12406 7704 13452 7732
rect 10689 7695 10747 7701
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 13538 7692 13544 7744
rect 13596 7732 13602 7744
rect 14093 7735 14151 7741
rect 14093 7732 14105 7735
rect 13596 7704 14105 7732
rect 13596 7692 13602 7704
rect 14093 7701 14105 7704
rect 14139 7701 14151 7735
rect 14093 7695 14151 7701
rect 14277 7735 14335 7741
rect 14277 7701 14289 7735
rect 14323 7732 14335 7735
rect 14458 7732 14464 7744
rect 14323 7704 14464 7732
rect 14323 7701 14335 7704
rect 14277 7695 14335 7701
rect 14458 7692 14464 7704
rect 14516 7692 14522 7744
rect 14734 7692 14740 7744
rect 14792 7732 14798 7744
rect 14829 7735 14887 7741
rect 14829 7732 14841 7735
rect 14792 7704 14841 7732
rect 14792 7692 14798 7704
rect 14829 7701 14841 7704
rect 14875 7732 14887 7735
rect 15010 7732 15016 7744
rect 14875 7704 15016 7732
rect 14875 7701 14887 7704
rect 14829 7695 14887 7701
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 15470 7732 15476 7744
rect 15431 7704 15476 7732
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 15654 7732 15660 7744
rect 15615 7704 15660 7732
rect 15654 7692 15660 7704
rect 15712 7692 15718 7744
rect 1104 7642 16008 7664
rect 1104 7590 4698 7642
rect 4750 7590 4762 7642
rect 4814 7590 4826 7642
rect 4878 7590 4890 7642
rect 4942 7590 4954 7642
rect 5006 7590 8446 7642
rect 8498 7590 8510 7642
rect 8562 7590 8574 7642
rect 8626 7590 8638 7642
rect 8690 7590 8702 7642
rect 8754 7590 12194 7642
rect 12246 7590 12258 7642
rect 12310 7590 12322 7642
rect 12374 7590 12386 7642
rect 12438 7590 12450 7642
rect 12502 7590 16008 7642
rect 1104 7568 16008 7590
rect 1670 7488 1676 7540
rect 1728 7528 1734 7540
rect 1765 7531 1823 7537
rect 1765 7528 1777 7531
rect 1728 7500 1777 7528
rect 1728 7488 1734 7500
rect 1765 7497 1777 7500
rect 1811 7497 1823 7531
rect 1765 7491 1823 7497
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 2593 7531 2651 7537
rect 2593 7528 2605 7531
rect 2096 7500 2605 7528
rect 2096 7488 2102 7500
rect 2593 7497 2605 7500
rect 2639 7497 2651 7531
rect 12989 7531 13047 7537
rect 12989 7528 13001 7531
rect 2593 7491 2651 7497
rect 2746 7500 13001 7528
rect 2746 7460 2774 7500
rect 12989 7497 13001 7500
rect 13035 7497 13047 7531
rect 12989 7491 13047 7497
rect 13446 7488 13452 7540
rect 13504 7528 13510 7540
rect 15010 7528 15016 7540
rect 13504 7500 15016 7528
rect 13504 7488 13510 7500
rect 15010 7488 15016 7500
rect 15068 7528 15074 7540
rect 15197 7531 15255 7537
rect 15068 7500 15148 7528
rect 15068 7488 15074 7500
rect 3142 7460 3148 7472
rect 1964 7432 2774 7460
rect 3103 7432 3148 7460
rect 1964 7401 1992 7432
rect 3142 7420 3148 7432
rect 3200 7420 3206 7472
rect 3789 7463 3847 7469
rect 3789 7429 3801 7463
rect 3835 7460 3847 7463
rect 3970 7460 3976 7472
rect 3835 7432 3976 7460
rect 3835 7429 3847 7432
rect 3789 7423 3847 7429
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7361 1731 7395
rect 1673 7355 1731 7361
rect 1949 7395 2007 7401
rect 1949 7361 1961 7395
rect 1995 7361 2007 7395
rect 1949 7355 2007 7361
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7392 2191 7395
rect 2406 7392 2412 7404
rect 2179 7364 2412 7392
rect 2179 7361 2191 7364
rect 2133 7355 2191 7361
rect 1688 7324 1716 7355
rect 2406 7352 2412 7364
rect 2464 7392 2470 7404
rect 3804 7392 3832 7423
rect 3970 7420 3976 7432
rect 4028 7420 4034 7472
rect 5166 7420 5172 7472
rect 5224 7460 5230 7472
rect 9861 7463 9919 7469
rect 5224 7432 8248 7460
rect 5224 7420 5230 7432
rect 2464 7364 3832 7392
rect 2464 7352 2470 7364
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 5442 7392 5448 7404
rect 5500 7401 5506 7404
rect 4212 7364 5448 7392
rect 4212 7352 4218 7364
rect 5442 7352 5448 7364
rect 5500 7355 5512 7401
rect 5500 7352 5506 7355
rect 5810 7352 5816 7404
rect 5868 7392 5874 7404
rect 6989 7395 7047 7401
rect 6989 7392 7001 7395
rect 5868 7364 7001 7392
rect 5868 7352 5874 7364
rect 6989 7361 7001 7364
rect 7035 7361 7047 7395
rect 6989 7355 7047 7361
rect 2222 7324 2228 7336
rect 1688 7296 2228 7324
rect 2222 7284 2228 7296
rect 2280 7284 2286 7336
rect 3237 7327 3295 7333
rect 3237 7293 3249 7327
rect 3283 7293 3295 7327
rect 3418 7324 3424 7336
rect 3379 7296 3424 7324
rect 3237 7287 3295 7293
rect 2314 7256 2320 7268
rect 2275 7228 2320 7256
rect 2314 7216 2320 7228
rect 2372 7216 2378 7268
rect 3252 7256 3280 7287
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7324 5779 7327
rect 6733 7327 6791 7333
rect 6733 7324 6745 7327
rect 5767 7296 5856 7324
rect 5767 7293 5779 7296
rect 5721 7287 5779 7293
rect 3510 7256 3516 7268
rect 3252 7228 3516 7256
rect 3510 7216 3516 7228
rect 3568 7256 3574 7268
rect 4065 7259 4123 7265
rect 4065 7256 4077 7259
rect 3568 7228 4077 7256
rect 3568 7216 3574 7228
rect 4065 7225 4077 7228
rect 4111 7256 4123 7259
rect 4614 7256 4620 7268
rect 4111 7228 4620 7256
rect 4111 7225 4123 7228
rect 4065 7219 4123 7225
rect 4614 7216 4620 7228
rect 4672 7216 4678 7268
rect 1486 7188 1492 7200
rect 1447 7160 1492 7188
rect 1486 7148 1492 7160
rect 1544 7148 1550 7200
rect 2498 7188 2504 7200
rect 2459 7160 2504 7188
rect 2498 7148 2504 7160
rect 2556 7148 2562 7200
rect 2777 7191 2835 7197
rect 2777 7157 2789 7191
rect 2823 7188 2835 7191
rect 3234 7188 3240 7200
rect 2823 7160 3240 7188
rect 2823 7157 2835 7160
rect 2777 7151 2835 7157
rect 3234 7148 3240 7160
rect 3292 7148 3298 7200
rect 3602 7148 3608 7200
rect 3660 7188 3666 7200
rect 3881 7191 3939 7197
rect 3881 7188 3893 7191
rect 3660 7160 3893 7188
rect 3660 7148 3666 7160
rect 3881 7157 3893 7160
rect 3927 7157 3939 7191
rect 4338 7188 4344 7200
rect 4299 7160 4344 7188
rect 3881 7151 3939 7157
rect 4338 7148 4344 7160
rect 4396 7148 4402 7200
rect 4430 7148 4436 7200
rect 4488 7188 4494 7200
rect 5442 7188 5448 7200
rect 4488 7160 5448 7188
rect 4488 7148 4494 7160
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 5828 7197 5856 7296
rect 6564 7296 6745 7324
rect 5813 7191 5871 7197
rect 5813 7157 5825 7191
rect 5859 7188 5871 7191
rect 6089 7191 6147 7197
rect 6089 7188 6101 7191
rect 5859 7160 6101 7188
rect 5859 7157 5871 7160
rect 5813 7151 5871 7157
rect 6089 7157 6101 7160
rect 6135 7188 6147 7191
rect 6454 7188 6460 7200
rect 6135 7160 6460 7188
rect 6135 7157 6147 7160
rect 6089 7151 6147 7157
rect 6454 7148 6460 7160
rect 6512 7188 6518 7200
rect 6564 7197 6592 7296
rect 6733 7293 6745 7296
rect 6779 7293 6791 7327
rect 6733 7287 6791 7293
rect 8220 7265 8248 7432
rect 9861 7429 9873 7463
rect 9907 7460 9919 7463
rect 10778 7460 10784 7472
rect 9907 7432 10784 7460
rect 9907 7429 9919 7432
rect 9861 7423 9919 7429
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 9306 7392 9312 7404
rect 9364 7401 9370 7404
rect 8444 7364 9312 7392
rect 8444 7352 8450 7364
rect 9306 7352 9312 7364
rect 9364 7392 9376 7401
rect 9582 7392 9588 7404
rect 9364 7364 9409 7392
rect 9495 7364 9588 7392
rect 9364 7355 9376 7364
rect 9364 7352 9370 7355
rect 9582 7352 9588 7364
rect 9640 7392 9646 7404
rect 9968 7401 9996 7432
rect 10778 7420 10784 7432
rect 10836 7460 10842 7472
rect 10836 7432 11560 7460
rect 10836 7420 10842 7432
rect 9953 7395 10011 7401
rect 9953 7392 9965 7395
rect 9640 7364 9965 7392
rect 9640 7352 9646 7364
rect 9953 7361 9965 7364
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 10220 7395 10278 7401
rect 10220 7361 10232 7395
rect 10266 7392 10278 7395
rect 11146 7392 11152 7404
rect 10266 7364 11152 7392
rect 10266 7361 10278 7364
rect 10220 7355 10278 7361
rect 11146 7352 11152 7364
rect 11204 7352 11210 7404
rect 11532 7336 11560 7432
rect 11606 7420 11612 7472
rect 11664 7460 11670 7472
rect 11762 7463 11820 7469
rect 11762 7460 11774 7463
rect 11664 7432 11774 7460
rect 11664 7420 11670 7432
rect 11762 7429 11774 7432
rect 11808 7460 11820 7463
rect 12710 7460 12716 7472
rect 11808 7432 12716 7460
rect 11808 7429 11820 7432
rect 11762 7423 11820 7429
rect 12710 7420 12716 7432
rect 12768 7420 12774 7472
rect 12894 7420 12900 7472
rect 12952 7460 12958 7472
rect 14185 7463 14243 7469
rect 12952 7432 13584 7460
rect 12952 7420 12958 7432
rect 13354 7392 13360 7404
rect 13315 7364 13360 7392
rect 13354 7352 13360 7364
rect 13412 7352 13418 7404
rect 11514 7324 11520 7336
rect 11475 7296 11520 7324
rect 11514 7284 11520 7296
rect 11572 7284 11578 7336
rect 13446 7324 13452 7336
rect 13407 7296 13452 7324
rect 13446 7284 13452 7296
rect 13504 7284 13510 7336
rect 13556 7333 13584 7432
rect 14185 7429 14197 7463
rect 14231 7460 14243 7463
rect 14550 7460 14556 7472
rect 14231 7432 14556 7460
rect 14231 7429 14243 7432
rect 14185 7423 14243 7429
rect 14550 7420 14556 7432
rect 14608 7420 14614 7472
rect 15120 7460 15148 7500
rect 15197 7497 15209 7531
rect 15243 7528 15255 7531
rect 15378 7528 15384 7540
rect 15243 7500 15384 7528
rect 15243 7497 15255 7500
rect 15197 7491 15255 7497
rect 15378 7488 15384 7500
rect 15436 7528 15442 7540
rect 15565 7531 15623 7537
rect 15565 7528 15577 7531
rect 15436 7500 15577 7528
rect 15436 7488 15442 7500
rect 15565 7497 15577 7500
rect 15611 7528 15623 7531
rect 15838 7528 15844 7540
rect 15611 7500 15844 7528
rect 15611 7497 15623 7500
rect 15565 7491 15623 7497
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 15120 7432 15240 7460
rect 15102 7392 15108 7404
rect 15063 7364 15108 7392
rect 15102 7352 15108 7364
rect 15160 7352 15166 7404
rect 15212 7392 15240 7432
rect 15212 7364 15332 7392
rect 13541 7327 13599 7333
rect 13541 7293 13553 7327
rect 13587 7293 13599 7327
rect 13541 7287 13599 7293
rect 14277 7327 14335 7333
rect 14277 7293 14289 7327
rect 14323 7293 14335 7327
rect 14277 7287 14335 7293
rect 8205 7259 8263 7265
rect 8205 7225 8217 7259
rect 8251 7225 8263 7259
rect 14292 7256 14320 7287
rect 14366 7284 14372 7336
rect 14424 7324 14430 7336
rect 15304 7333 15332 7364
rect 15289 7327 15347 7333
rect 14424 7296 14469 7324
rect 14424 7284 14430 7296
rect 15289 7293 15301 7327
rect 15335 7293 15347 7327
rect 15289 7287 15347 7293
rect 15562 7256 15568 7268
rect 8205 7219 8263 7225
rect 13648 7228 15568 7256
rect 6549 7191 6607 7197
rect 6549 7188 6561 7191
rect 6512 7160 6561 7188
rect 6512 7148 6518 7160
rect 6549 7157 6561 7160
rect 6595 7157 6607 7191
rect 6549 7151 6607 7157
rect 7006 7148 7012 7200
rect 7064 7188 7070 7200
rect 8110 7188 8116 7200
rect 7064 7160 8116 7188
rect 7064 7148 7070 7160
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 11330 7188 11336 7200
rect 11291 7160 11336 7188
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13170 7148 13176 7200
rect 13228 7188 13234 7200
rect 13648 7188 13676 7228
rect 15562 7216 15568 7228
rect 15620 7216 15626 7268
rect 13814 7188 13820 7200
rect 13228 7160 13676 7188
rect 13775 7160 13820 7188
rect 13228 7148 13234 7160
rect 13814 7148 13820 7160
rect 13872 7148 13878 7200
rect 13998 7148 14004 7200
rect 14056 7188 14062 7200
rect 14550 7188 14556 7200
rect 14056 7160 14556 7188
rect 14056 7148 14062 7160
rect 14550 7148 14556 7160
rect 14608 7148 14614 7200
rect 14734 7188 14740 7200
rect 14695 7160 14740 7188
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 1104 7098 16008 7120
rect 1104 7046 2824 7098
rect 2876 7046 2888 7098
rect 2940 7046 2952 7098
rect 3004 7046 3016 7098
rect 3068 7046 3080 7098
rect 3132 7046 6572 7098
rect 6624 7046 6636 7098
rect 6688 7046 6700 7098
rect 6752 7046 6764 7098
rect 6816 7046 6828 7098
rect 6880 7046 10320 7098
rect 10372 7046 10384 7098
rect 10436 7046 10448 7098
rect 10500 7046 10512 7098
rect 10564 7046 10576 7098
rect 10628 7046 14068 7098
rect 14120 7046 14132 7098
rect 14184 7046 14196 7098
rect 14248 7046 14260 7098
rect 14312 7046 14324 7098
rect 14376 7046 16008 7098
rect 1104 7024 16008 7046
rect 1949 6987 2007 6993
rect 1949 6953 1961 6987
rect 1995 6984 2007 6987
rect 2038 6984 2044 6996
rect 1995 6956 2044 6984
rect 1995 6953 2007 6956
rect 1949 6947 2007 6953
rect 2038 6944 2044 6956
rect 2096 6944 2102 6996
rect 7285 6987 7343 6993
rect 7285 6953 7297 6987
rect 7331 6984 7343 6987
rect 8386 6984 8392 6996
rect 7331 6956 8392 6984
rect 7331 6953 7343 6956
rect 7285 6947 7343 6953
rect 8386 6944 8392 6956
rect 8444 6944 8450 6996
rect 9033 6987 9091 6993
rect 9033 6953 9045 6987
rect 9079 6984 9091 6987
rect 9582 6984 9588 6996
rect 9079 6956 9588 6984
rect 9079 6953 9091 6956
rect 9033 6947 9091 6953
rect 4154 6876 4160 6928
rect 4212 6876 4218 6928
rect 1578 6848 1584 6860
rect 1539 6820 1584 6848
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 1765 6851 1823 6857
rect 1765 6817 1777 6851
rect 1811 6848 1823 6851
rect 1946 6848 1952 6860
rect 1811 6820 1952 6848
rect 1811 6817 1823 6820
rect 1765 6811 1823 6817
rect 1946 6808 1952 6820
rect 2004 6848 2010 6860
rect 2130 6848 2136 6860
rect 2004 6820 2136 6848
rect 2004 6808 2010 6820
rect 2130 6808 2136 6820
rect 2188 6808 2194 6860
rect 3326 6808 3332 6860
rect 3384 6808 3390 6860
rect 3421 6851 3479 6857
rect 3421 6817 3433 6851
rect 3467 6848 3479 6851
rect 4172 6848 4200 6876
rect 3467 6820 4200 6848
rect 8757 6851 8815 6857
rect 3467 6817 3479 6820
rect 3421 6811 3479 6817
rect 8757 6817 8769 6851
rect 8803 6848 8815 6851
rect 9048 6848 9076 6947
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 13078 6944 13084 6996
rect 13136 6984 13142 6996
rect 13909 6987 13967 6993
rect 13136 6956 13768 6984
rect 13136 6944 13142 6956
rect 8803 6820 9076 6848
rect 13357 6851 13415 6857
rect 8803 6817 8815 6820
rect 8757 6811 8815 6817
rect 13357 6817 13369 6851
rect 13403 6848 13415 6851
rect 13630 6848 13636 6860
rect 13403 6820 13636 6848
rect 13403 6817 13415 6820
rect 13357 6811 13415 6817
rect 1394 6740 1400 6792
rect 1452 6780 1458 6792
rect 1854 6780 1860 6792
rect 1452 6752 1860 6780
rect 1452 6740 1458 6752
rect 1854 6740 1860 6752
rect 1912 6780 1918 6792
rect 2590 6780 2596 6792
rect 1912 6752 2596 6780
rect 1912 6740 1918 6752
rect 2590 6740 2596 6752
rect 2648 6740 2654 6792
rect 3344 6780 3372 6808
rect 3878 6780 3884 6792
rect 3344 6752 3884 6780
rect 3878 6740 3884 6752
rect 3936 6740 3942 6792
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6780 4215 6783
rect 5813 6783 5871 6789
rect 5813 6780 5825 6783
rect 4203 6752 5825 6780
rect 4203 6749 4215 6752
rect 4157 6743 4215 6749
rect 5813 6749 5825 6752
rect 5859 6780 5871 6783
rect 5905 6783 5963 6789
rect 5905 6780 5917 6783
rect 5859 6752 5917 6780
rect 5859 6749 5871 6752
rect 5813 6743 5871 6749
rect 5905 6749 5917 6752
rect 5951 6780 5963 6783
rect 6454 6780 6460 6792
rect 5951 6752 6460 6780
rect 5951 6749 5963 6752
rect 5905 6743 5963 6749
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 10413 6783 10471 6789
rect 10413 6749 10425 6783
rect 10459 6780 10471 6783
rect 11885 6783 11943 6789
rect 11885 6780 11897 6783
rect 10459 6752 11897 6780
rect 10459 6749 10471 6752
rect 10413 6743 10471 6749
rect 11885 6749 11897 6752
rect 11931 6780 11943 6783
rect 12066 6780 12072 6792
rect 11931 6752 12072 6780
rect 11931 6749 11943 6752
rect 11885 6743 11943 6749
rect 12066 6740 12072 6752
rect 12124 6780 12130 6792
rect 13372 6780 13400 6811
rect 13630 6808 13636 6820
rect 13688 6808 13694 6860
rect 13740 6848 13768 6956
rect 13909 6953 13921 6987
rect 13955 6984 13967 6987
rect 14550 6984 14556 6996
rect 13955 6956 14556 6984
rect 13955 6953 13967 6956
rect 13909 6947 13967 6953
rect 14550 6944 14556 6956
rect 14608 6944 14614 6996
rect 14568 6916 14596 6944
rect 14568 6888 14872 6916
rect 14645 6851 14703 6857
rect 14645 6848 14657 6851
rect 13740 6820 14657 6848
rect 14645 6817 14657 6820
rect 14691 6817 14703 6851
rect 14645 6811 14703 6817
rect 12124 6752 13400 6780
rect 13725 6783 13783 6789
rect 12124 6740 12130 6752
rect 13725 6749 13737 6783
rect 13771 6780 13783 6783
rect 13906 6780 13912 6792
rect 13771 6752 13912 6780
rect 13771 6749 13783 6752
rect 13725 6743 13783 6749
rect 13906 6740 13912 6752
rect 13964 6740 13970 6792
rect 14461 6783 14519 6789
rect 14461 6749 14473 6783
rect 14507 6780 14519 6783
rect 14734 6780 14740 6792
rect 14507 6752 14740 6780
rect 14507 6749 14519 6752
rect 14461 6743 14519 6749
rect 14734 6740 14740 6752
rect 14792 6740 14798 6792
rect 2317 6715 2375 6721
rect 2317 6681 2329 6715
rect 2363 6712 2375 6715
rect 2682 6712 2688 6724
rect 2363 6684 2688 6712
rect 2363 6681 2375 6684
rect 2317 6675 2375 6681
rect 2682 6672 2688 6684
rect 2740 6672 2746 6724
rect 3326 6672 3332 6724
rect 3384 6712 3390 6724
rect 4402 6715 4460 6721
rect 4402 6712 4414 6715
rect 3384 6684 4414 6712
rect 3384 6672 3390 6684
rect 4402 6681 4414 6684
rect 4448 6681 4460 6715
rect 4402 6675 4460 6681
rect 6172 6715 6230 6721
rect 6172 6681 6184 6715
rect 6218 6712 6230 6715
rect 8512 6715 8570 6721
rect 6218 6684 7972 6712
rect 6218 6681 6230 6684
rect 6172 6675 6230 6681
rect 2130 6644 2136 6656
rect 2091 6616 2136 6644
rect 2130 6604 2136 6616
rect 2188 6604 2194 6656
rect 2498 6644 2504 6656
rect 2459 6616 2504 6644
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 2774 6604 2780 6656
rect 2832 6644 2838 6656
rect 3142 6644 3148 6656
rect 2832 6616 2877 6644
rect 3103 6616 3148 6644
rect 2832 6604 2838 6616
rect 3142 6604 3148 6616
rect 3200 6604 3206 6656
rect 3237 6647 3295 6653
rect 3237 6613 3249 6647
rect 3283 6644 3295 6647
rect 3418 6644 3424 6656
rect 3283 6616 3424 6644
rect 3283 6613 3295 6616
rect 3237 6607 3295 6613
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3786 6644 3792 6656
rect 3747 6616 3792 6644
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 5534 6644 5540 6656
rect 5495 6616 5540 6644
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 7374 6604 7380 6656
rect 7432 6644 7438 6656
rect 7944 6644 7972 6684
rect 8512 6681 8524 6715
rect 8558 6712 8570 6715
rect 11238 6712 11244 6724
rect 8558 6684 11244 6712
rect 8558 6681 8570 6684
rect 8512 6675 8570 6681
rect 11238 6672 11244 6684
rect 11296 6672 11302 6724
rect 11330 6672 11336 6724
rect 11388 6712 11394 6724
rect 11618 6715 11676 6721
rect 11618 6712 11630 6715
rect 11388 6684 11630 6712
rect 11388 6672 11394 6684
rect 11618 6681 11630 6684
rect 11664 6681 11676 6715
rect 11618 6675 11676 6681
rect 12894 6672 12900 6724
rect 12952 6712 12958 6724
rect 13090 6715 13148 6721
rect 13090 6712 13102 6715
rect 12952 6684 13102 6712
rect 12952 6672 12958 6684
rect 13090 6681 13102 6684
rect 13136 6712 13148 6715
rect 13262 6712 13268 6724
rect 13136 6684 13268 6712
rect 13136 6681 13148 6684
rect 13090 6675 13148 6681
rect 13262 6672 13268 6684
rect 13320 6672 13326 6724
rect 13354 6672 13360 6724
rect 13412 6712 13418 6724
rect 14844 6712 14872 6888
rect 15010 6876 15016 6928
rect 15068 6916 15074 6928
rect 15068 6888 15516 6916
rect 15068 6876 15074 6888
rect 15488 6857 15516 6888
rect 15473 6851 15531 6857
rect 15473 6817 15485 6851
rect 15519 6817 15531 6851
rect 15473 6811 15531 6817
rect 14918 6740 14924 6792
rect 14976 6780 14982 6792
rect 15381 6783 15439 6789
rect 15381 6780 15393 6783
rect 14976 6752 15393 6780
rect 14976 6740 14982 6752
rect 15381 6749 15393 6752
rect 15427 6749 15439 6783
rect 15381 6743 15439 6749
rect 15286 6712 15292 6724
rect 13412 6684 14136 6712
rect 14844 6684 15292 6712
rect 13412 6672 13418 6684
rect 9674 6644 9680 6656
rect 7432 6616 7477 6644
rect 7944 6616 9680 6644
rect 7432 6604 7438 6616
rect 9674 6604 9680 6616
rect 9732 6644 9738 6656
rect 10505 6647 10563 6653
rect 10505 6644 10517 6647
rect 9732 6616 10517 6644
rect 9732 6604 9738 6616
rect 10505 6613 10517 6616
rect 10551 6613 10563 6647
rect 11974 6644 11980 6656
rect 11935 6616 11980 6644
rect 10505 6607 10563 6613
rect 11974 6604 11980 6616
rect 12032 6604 12038 6656
rect 13541 6647 13599 6653
rect 13541 6613 13553 6647
rect 13587 6644 13599 6647
rect 13630 6644 13636 6656
rect 13587 6616 13636 6644
rect 13587 6613 13599 6616
rect 13541 6607 13599 6613
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 14108 6653 14136 6684
rect 15286 6672 15292 6684
rect 15344 6672 15350 6724
rect 14093 6647 14151 6653
rect 14093 6613 14105 6647
rect 14139 6613 14151 6647
rect 14093 6607 14151 6613
rect 14550 6604 14556 6656
rect 14608 6644 14614 6656
rect 14608 6616 14653 6644
rect 14608 6604 14614 6616
rect 14734 6604 14740 6656
rect 14792 6644 14798 6656
rect 14921 6647 14979 6653
rect 14921 6644 14933 6647
rect 14792 6616 14933 6644
rect 14792 6604 14798 6616
rect 14921 6613 14933 6616
rect 14967 6613 14979 6647
rect 14921 6607 14979 6613
rect 1104 6554 16008 6576
rect 1104 6502 4698 6554
rect 4750 6502 4762 6554
rect 4814 6502 4826 6554
rect 4878 6502 4890 6554
rect 4942 6502 4954 6554
rect 5006 6502 8446 6554
rect 8498 6502 8510 6554
rect 8562 6502 8574 6554
rect 8626 6502 8638 6554
rect 8690 6502 8702 6554
rect 8754 6502 12194 6554
rect 12246 6502 12258 6554
rect 12310 6502 12322 6554
rect 12374 6502 12386 6554
rect 12438 6502 12450 6554
rect 12502 6502 16008 6554
rect 1104 6480 16008 6502
rect 2041 6443 2099 6449
rect 2041 6440 2053 6443
rect 1688 6412 2053 6440
rect 1688 6313 1716 6412
rect 2041 6409 2053 6412
rect 2087 6409 2099 6443
rect 2041 6403 2099 6409
rect 2869 6443 2927 6449
rect 2869 6409 2881 6443
rect 2915 6440 2927 6443
rect 3786 6440 3792 6452
rect 2915 6412 3792 6440
rect 2915 6409 2927 6412
rect 2869 6403 2927 6409
rect 3786 6400 3792 6412
rect 3844 6400 3850 6452
rect 6181 6443 6239 6449
rect 6181 6409 6193 6443
rect 6227 6440 6239 6443
rect 6270 6440 6276 6452
rect 6227 6412 6276 6440
rect 6227 6409 6239 6412
rect 6181 6403 6239 6409
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 7926 6440 7932 6452
rect 6564 6412 7932 6440
rect 2774 6372 2780 6384
rect 1964 6344 2780 6372
rect 1964 6313 1992 6344
rect 2774 6332 2780 6344
rect 2832 6332 2838 6384
rect 2961 6375 3019 6381
rect 2961 6341 2973 6375
rect 3007 6372 3019 6375
rect 3510 6372 3516 6384
rect 3007 6344 3516 6372
rect 3007 6341 3019 6344
rect 2961 6335 3019 6341
rect 3510 6332 3516 6344
rect 3568 6332 3574 6384
rect 4338 6332 4344 6384
rect 4396 6372 4402 6384
rect 4442 6375 4500 6381
rect 4442 6372 4454 6375
rect 4396 6344 4454 6372
rect 4396 6332 4402 6344
rect 4442 6341 4454 6344
rect 4488 6341 4500 6375
rect 6454 6372 6460 6384
rect 4442 6335 4500 6341
rect 4816 6344 6460 6372
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 2222 6304 2228 6316
rect 2183 6276 2228 6304
rect 1949 6267 2007 6273
rect 2222 6264 2228 6276
rect 2280 6264 2286 6316
rect 2590 6264 2596 6316
rect 2648 6304 2654 6316
rect 4816 6313 4844 6344
rect 6454 6332 6460 6344
rect 6512 6332 6518 6384
rect 4709 6307 4767 6313
rect 2648 6276 4660 6304
rect 2648 6264 2654 6276
rect 2409 6239 2467 6245
rect 2409 6205 2421 6239
rect 2455 6236 2467 6239
rect 2774 6236 2780 6248
rect 2455 6208 2780 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 2774 6196 2780 6208
rect 2832 6196 2838 6248
rect 3145 6239 3203 6245
rect 3145 6205 3157 6239
rect 3191 6236 3203 6239
rect 3234 6236 3240 6248
rect 3191 6208 3240 6236
rect 3191 6205 3203 6208
rect 3145 6199 3203 6205
rect 3234 6196 3240 6208
rect 3292 6196 3298 6248
rect 4632 6236 4660 6276
rect 4709 6273 4721 6307
rect 4755 6304 4767 6307
rect 4801 6307 4859 6313
rect 4801 6304 4813 6307
rect 4755 6276 4813 6304
rect 4755 6273 4767 6276
rect 4709 6267 4767 6273
rect 4801 6273 4813 6276
rect 4847 6273 4859 6307
rect 5057 6307 5115 6313
rect 5057 6304 5069 6307
rect 4801 6267 4859 6273
rect 4908 6276 5069 6304
rect 4908 6236 4936 6276
rect 5057 6273 5069 6276
rect 5103 6304 5115 6307
rect 5534 6304 5540 6316
rect 5103 6276 5540 6304
rect 5103 6273 5115 6276
rect 5057 6267 5115 6273
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 5994 6264 6000 6316
rect 6052 6304 6058 6316
rect 6564 6304 6592 6412
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 9950 6400 9956 6452
rect 10008 6440 10014 6452
rect 11149 6443 11207 6449
rect 11149 6440 11161 6443
rect 10008 6412 11161 6440
rect 10008 6400 10014 6412
rect 11149 6409 11161 6412
rect 11195 6440 11207 6443
rect 11422 6440 11428 6452
rect 11195 6412 11428 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 11422 6400 11428 6412
rect 11480 6400 11486 6452
rect 11514 6400 11520 6452
rect 11572 6440 11578 6452
rect 11609 6443 11667 6449
rect 11609 6440 11621 6443
rect 11572 6412 11621 6440
rect 11572 6400 11578 6412
rect 11609 6409 11621 6412
rect 11655 6440 11667 6443
rect 11885 6443 11943 6449
rect 11885 6440 11897 6443
rect 11655 6412 11897 6440
rect 11655 6409 11667 6412
rect 11609 6403 11667 6409
rect 11885 6409 11897 6412
rect 11931 6440 11943 6443
rect 12066 6440 12072 6452
rect 11931 6412 12072 6440
rect 11931 6409 11943 6412
rect 11885 6403 11943 6409
rect 12066 6400 12072 6412
rect 12124 6400 12130 6452
rect 12158 6400 12164 6452
rect 12216 6440 12222 6452
rect 12345 6443 12403 6449
rect 12345 6440 12357 6443
rect 12216 6412 12357 6440
rect 12216 6400 12222 6412
rect 12345 6409 12357 6412
rect 12391 6409 12403 6443
rect 12345 6403 12403 6409
rect 13173 6443 13231 6449
rect 13173 6409 13185 6443
rect 13219 6440 13231 6443
rect 13725 6443 13783 6449
rect 13725 6440 13737 6443
rect 13219 6412 13737 6440
rect 13219 6409 13231 6412
rect 13173 6403 13231 6409
rect 13725 6409 13737 6412
rect 13771 6409 13783 6443
rect 13725 6403 13783 6409
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 14185 6443 14243 6449
rect 14185 6440 14197 6443
rect 13872 6412 14197 6440
rect 13872 6400 13878 6412
rect 14185 6409 14197 6412
rect 14231 6409 14243 6443
rect 14550 6440 14556 6452
rect 14511 6412 14556 6440
rect 14185 6403 14243 6409
rect 14550 6400 14556 6412
rect 14608 6400 14614 6452
rect 14826 6400 14832 6452
rect 14884 6440 14890 6452
rect 14921 6443 14979 6449
rect 14921 6440 14933 6443
rect 14884 6412 14933 6440
rect 14884 6400 14890 6412
rect 14921 6409 14933 6412
rect 14967 6440 14979 6443
rect 15746 6440 15752 6452
rect 14967 6412 15752 6440
rect 14967 6409 14979 6412
rect 14921 6403 14979 6409
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 7650 6332 7656 6384
rect 7708 6372 7714 6384
rect 7834 6372 7840 6384
rect 7708 6344 7840 6372
rect 7708 6332 7714 6344
rect 7834 6332 7840 6344
rect 7892 6332 7898 6384
rect 8754 6332 8760 6384
rect 8812 6372 8818 6384
rect 10781 6375 10839 6381
rect 10781 6372 10793 6375
rect 8812 6344 10793 6372
rect 8812 6332 8818 6344
rect 10781 6341 10793 6344
rect 10827 6372 10839 6375
rect 10962 6372 10968 6384
rect 10827 6344 10968 6372
rect 10827 6341 10839 6344
rect 10781 6335 10839 6341
rect 10962 6332 10968 6344
rect 11020 6332 11026 6384
rect 11698 6332 11704 6384
rect 11756 6372 11762 6384
rect 11977 6375 12035 6381
rect 11977 6372 11989 6375
rect 11756 6344 11989 6372
rect 11756 6332 11762 6344
rect 11977 6341 11989 6344
rect 12023 6341 12035 6375
rect 11977 6335 12035 6341
rect 13265 6375 13323 6381
rect 13265 6341 13277 6375
rect 13311 6372 13323 6375
rect 14734 6372 14740 6384
rect 13311 6344 14740 6372
rect 13311 6341 13323 6344
rect 13265 6335 13323 6341
rect 14734 6332 14740 6344
rect 14792 6332 14798 6384
rect 15010 6372 15016 6384
rect 14844 6344 15016 6372
rect 6052 6276 6592 6304
rect 7460 6307 7518 6313
rect 6052 6264 6058 6276
rect 7460 6273 7472 6307
rect 7506 6304 7518 6307
rect 7926 6304 7932 6316
rect 7506 6276 7932 6304
rect 7506 6273 7518 6276
rect 7460 6267 7518 6273
rect 7926 6264 7932 6276
rect 7984 6264 7990 6316
rect 8938 6313 8944 6316
rect 8932 6304 8944 6313
rect 8899 6276 8944 6304
rect 8932 6267 8944 6276
rect 8938 6264 8944 6267
rect 8996 6264 9002 6316
rect 9306 6264 9312 6316
rect 9364 6304 9370 6316
rect 9364 6276 12296 6304
rect 9364 6264 9370 6276
rect 6454 6236 6460 6248
rect 4632 6208 4752 6236
rect 4724 6180 4752 6208
rect 4816 6208 4936 6236
rect 6367 6208 6460 6236
rect 1486 6168 1492 6180
rect 1447 6140 1492 6168
rect 1486 6128 1492 6140
rect 1544 6128 1550 6180
rect 2590 6128 2596 6180
rect 2648 6168 2654 6180
rect 2648 6140 2774 6168
rect 2648 6128 2654 6140
rect 1670 6060 1676 6112
rect 1728 6100 1734 6112
rect 1765 6103 1823 6109
rect 1765 6100 1777 6103
rect 1728 6072 1777 6100
rect 1728 6060 1734 6072
rect 1765 6069 1777 6072
rect 1811 6069 1823 6103
rect 1765 6063 1823 6069
rect 2038 6060 2044 6112
rect 2096 6100 2102 6112
rect 2501 6103 2559 6109
rect 2501 6100 2513 6103
rect 2096 6072 2513 6100
rect 2096 6060 2102 6072
rect 2501 6069 2513 6072
rect 2547 6069 2559 6103
rect 2746 6100 2774 6140
rect 3160 6140 3832 6168
rect 3160 6100 3188 6140
rect 2746 6072 3188 6100
rect 2501 6063 2559 6069
rect 3234 6060 3240 6112
rect 3292 6100 3298 6112
rect 3329 6103 3387 6109
rect 3329 6100 3341 6103
rect 3292 6072 3341 6100
rect 3292 6060 3298 6072
rect 3329 6069 3341 6072
rect 3375 6069 3387 6103
rect 3804 6100 3832 6140
rect 4706 6128 4712 6180
rect 4764 6128 4770 6180
rect 4816 6100 4844 6208
rect 6454 6196 6460 6208
rect 6512 6236 6518 6248
rect 6641 6239 6699 6245
rect 6641 6236 6653 6239
rect 6512 6208 6653 6236
rect 6512 6196 6518 6208
rect 6641 6205 6653 6208
rect 6687 6236 6699 6239
rect 7101 6239 7159 6245
rect 7101 6236 7113 6239
rect 6687 6208 7113 6236
rect 6687 6205 6699 6208
rect 6641 6199 6699 6205
rect 7101 6205 7113 6208
rect 7147 6236 7159 6239
rect 7190 6236 7196 6248
rect 7147 6208 7196 6236
rect 7147 6205 7159 6208
rect 7101 6199 7159 6205
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 8662 6236 8668 6248
rect 8623 6208 8668 6236
rect 8662 6196 8668 6208
rect 8720 6196 8726 6248
rect 11882 6196 11888 6248
rect 11940 6236 11946 6248
rect 12158 6236 12164 6248
rect 11940 6208 12164 6236
rect 11940 6196 11946 6208
rect 12158 6196 12164 6208
rect 12216 6196 12222 6248
rect 12268 6236 12296 6276
rect 12342 6264 12348 6316
rect 12400 6304 12406 6316
rect 12529 6307 12587 6313
rect 12529 6304 12541 6307
rect 12400 6276 12541 6304
rect 12400 6264 12406 6276
rect 12529 6273 12541 6276
rect 12575 6273 12587 6307
rect 14090 6304 14096 6316
rect 14051 6276 14096 6304
rect 12529 6267 12587 6273
rect 14090 6264 14096 6276
rect 14148 6264 14154 6316
rect 12618 6236 12624 6248
rect 12268 6208 12624 6236
rect 12618 6196 12624 6208
rect 12676 6196 12682 6248
rect 13078 6236 13084 6248
rect 13039 6208 13084 6236
rect 13078 6196 13084 6208
rect 13136 6196 13142 6248
rect 14369 6239 14427 6245
rect 14369 6205 14381 6239
rect 14415 6236 14427 6239
rect 14844 6236 14872 6344
rect 15010 6332 15016 6344
rect 15068 6332 15074 6384
rect 15028 6304 15056 6332
rect 15378 6304 15384 6316
rect 15028 6276 15148 6304
rect 15339 6276 15384 6304
rect 15120 6245 15148 6276
rect 15378 6264 15384 6276
rect 15436 6264 15442 6316
rect 14415 6208 14872 6236
rect 15013 6239 15071 6245
rect 14415 6205 14427 6208
rect 14369 6199 14427 6205
rect 15013 6205 15025 6239
rect 15059 6205 15071 6239
rect 15013 6199 15071 6205
rect 15105 6239 15163 6245
rect 15105 6205 15117 6239
rect 15151 6205 15163 6239
rect 15105 6199 15163 6205
rect 5736 6140 6868 6168
rect 3804 6072 4844 6100
rect 3329 6063 3387 6069
rect 5166 6060 5172 6112
rect 5224 6100 5230 6112
rect 5736 6100 5764 6140
rect 5224 6072 5764 6100
rect 5224 6060 5230 6072
rect 6362 6060 6368 6112
rect 6420 6100 6426 6112
rect 6733 6103 6791 6109
rect 6733 6100 6745 6103
rect 6420 6072 6745 6100
rect 6420 6060 6426 6072
rect 6733 6069 6745 6072
rect 6779 6069 6791 6103
rect 6840 6100 6868 6140
rect 13446 6128 13452 6180
rect 13504 6168 13510 6180
rect 13633 6171 13691 6177
rect 13633 6168 13645 6171
rect 13504 6140 13645 6168
rect 13504 6128 13510 6140
rect 13633 6137 13645 6140
rect 13679 6137 13691 6171
rect 13633 6131 13691 6137
rect 13722 6128 13728 6180
rect 13780 6168 13786 6180
rect 15028 6168 15056 6199
rect 13780 6140 15056 6168
rect 13780 6128 13786 6140
rect 8110 6100 8116 6112
rect 6840 6072 8116 6100
rect 6733 6063 6791 6069
rect 8110 6060 8116 6072
rect 8168 6060 8174 6112
rect 8573 6103 8631 6109
rect 8573 6069 8585 6103
rect 8619 6100 8631 6103
rect 8938 6100 8944 6112
rect 8619 6072 8944 6100
rect 8619 6069 8631 6072
rect 8573 6063 8631 6069
rect 8938 6060 8944 6072
rect 8996 6060 9002 6112
rect 9766 6060 9772 6112
rect 9824 6100 9830 6112
rect 10045 6103 10103 6109
rect 10045 6100 10057 6103
rect 9824 6072 10057 6100
rect 9824 6060 9830 6072
rect 10045 6069 10057 6072
rect 10091 6069 10103 6103
rect 10045 6063 10103 6069
rect 11333 6103 11391 6109
rect 11333 6069 11345 6103
rect 11379 6100 11391 6103
rect 11606 6100 11612 6112
rect 11379 6072 11612 6100
rect 11379 6069 11391 6072
rect 11333 6063 11391 6069
rect 11606 6060 11612 6072
rect 11664 6060 11670 6112
rect 12158 6100 12164 6112
rect 12119 6072 12164 6100
rect 12158 6060 12164 6072
rect 12216 6060 12222 6112
rect 12805 6103 12863 6109
rect 12805 6069 12817 6103
rect 12851 6100 12863 6103
rect 12986 6100 12992 6112
rect 12851 6072 12992 6100
rect 12851 6069 12863 6072
rect 12805 6063 12863 6069
rect 12986 6060 12992 6072
rect 13044 6060 13050 6112
rect 15562 6100 15568 6112
rect 15523 6072 15568 6100
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 1104 6010 16008 6032
rect 1104 5958 2824 6010
rect 2876 5958 2888 6010
rect 2940 5958 2952 6010
rect 3004 5958 3016 6010
rect 3068 5958 3080 6010
rect 3132 5958 6572 6010
rect 6624 5958 6636 6010
rect 6688 5958 6700 6010
rect 6752 5958 6764 6010
rect 6816 5958 6828 6010
rect 6880 5958 10320 6010
rect 10372 5958 10384 6010
rect 10436 5958 10448 6010
rect 10500 5958 10512 6010
rect 10564 5958 10576 6010
rect 10628 5958 14068 6010
rect 14120 5958 14132 6010
rect 14184 5958 14196 6010
rect 14248 5958 14260 6010
rect 14312 5958 14324 6010
rect 14376 5958 16008 6010
rect 1104 5936 16008 5958
rect 2593 5899 2651 5905
rect 2593 5865 2605 5899
rect 2639 5896 2651 5899
rect 3050 5896 3056 5908
rect 2639 5868 3056 5896
rect 2639 5865 2651 5868
rect 2593 5859 2651 5865
rect 3050 5856 3056 5868
rect 3108 5856 3114 5908
rect 3418 5896 3424 5908
rect 3379 5868 3424 5896
rect 3418 5856 3424 5868
rect 3476 5856 3482 5908
rect 5810 5896 5816 5908
rect 5771 5868 5816 5896
rect 5810 5856 5816 5868
rect 5868 5896 5874 5908
rect 6270 5896 6276 5908
rect 5868 5868 6276 5896
rect 5868 5856 5874 5868
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 7377 5899 7435 5905
rect 7377 5896 7389 5899
rect 7248 5868 7389 5896
rect 7248 5856 7254 5868
rect 7377 5865 7389 5868
rect 7423 5896 7435 5899
rect 8294 5896 8300 5908
rect 7423 5868 8300 5896
rect 7423 5865 7435 5868
rect 7377 5859 7435 5865
rect 1394 5788 1400 5840
rect 1452 5828 1458 5840
rect 1946 5828 1952 5840
rect 1452 5800 1952 5828
rect 1452 5788 1458 5800
rect 1946 5788 1952 5800
rect 2004 5828 2010 5840
rect 3789 5831 3847 5837
rect 3789 5828 3801 5831
rect 2004 5800 3801 5828
rect 2004 5788 2010 5800
rect 2148 5769 2176 5800
rect 3789 5797 3801 5800
rect 3835 5797 3847 5831
rect 3789 5791 3847 5797
rect 2041 5763 2099 5769
rect 2041 5729 2053 5763
rect 2087 5729 2099 5763
rect 2041 5723 2099 5729
rect 2133 5763 2191 5769
rect 2133 5729 2145 5763
rect 2179 5729 2191 5763
rect 2866 5760 2872 5772
rect 2779 5732 2872 5760
rect 2133 5723 2191 5729
rect 1670 5692 1676 5704
rect 1631 5664 1676 5692
rect 1670 5652 1676 5664
rect 1728 5652 1734 5704
rect 2056 5692 2084 5723
rect 2866 5720 2872 5732
rect 2924 5760 2930 5772
rect 4062 5760 4068 5772
rect 2924 5732 4068 5760
rect 2924 5720 2930 5732
rect 4062 5720 4068 5732
rect 4120 5720 4126 5772
rect 7193 5763 7251 5769
rect 7193 5729 7205 5763
rect 7239 5760 7251 5763
rect 7392 5760 7420 5859
rect 8294 5856 8300 5868
rect 8352 5896 8358 5908
rect 8573 5899 8631 5905
rect 8573 5896 8585 5899
rect 8352 5868 8585 5896
rect 8352 5856 8358 5868
rect 8573 5865 8585 5868
rect 8619 5896 8631 5899
rect 8662 5896 8668 5908
rect 8619 5868 8668 5896
rect 8619 5865 8631 5868
rect 8573 5859 8631 5865
rect 8662 5856 8668 5868
rect 8720 5896 8726 5908
rect 9582 5896 9588 5908
rect 8720 5868 9588 5896
rect 8720 5856 8726 5868
rect 9582 5856 9588 5868
rect 9640 5856 9646 5908
rect 10686 5896 10692 5908
rect 9784 5868 10692 5896
rect 7558 5828 7564 5840
rect 7519 5800 7564 5828
rect 7558 5788 7564 5800
rect 7616 5788 7622 5840
rect 7742 5828 7748 5840
rect 7703 5800 7748 5828
rect 7742 5788 7748 5800
rect 7800 5788 7806 5840
rect 7834 5788 7840 5840
rect 7892 5828 7898 5840
rect 8110 5828 8116 5840
rect 7892 5800 7937 5828
rect 8023 5800 8116 5828
rect 7892 5788 7898 5800
rect 8110 5788 8116 5800
rect 8168 5828 8174 5840
rect 9784 5828 9812 5868
rect 10686 5856 10692 5868
rect 10744 5856 10750 5908
rect 11238 5896 11244 5908
rect 11199 5868 11244 5896
rect 11238 5856 11244 5868
rect 11296 5856 11302 5908
rect 12710 5856 12716 5908
rect 12768 5896 12774 5908
rect 12768 5868 13400 5896
rect 12768 5856 12774 5868
rect 11146 5828 11152 5840
rect 8168 5800 9812 5828
rect 11107 5800 11152 5828
rect 8168 5788 8174 5800
rect 11146 5788 11152 5800
rect 11204 5788 11210 5840
rect 12618 5788 12624 5840
rect 12676 5828 12682 5840
rect 12676 5800 13308 5828
rect 12676 5788 12682 5800
rect 7239 5732 7420 5760
rect 7239 5729 7251 5732
rect 7193 5723 7251 5729
rect 8386 5720 8392 5772
rect 8444 5760 8450 5772
rect 9306 5760 9312 5772
rect 8444 5732 9312 5760
rect 8444 5720 8450 5732
rect 9306 5720 9312 5732
rect 9364 5720 9370 5772
rect 9582 5720 9588 5772
rect 9640 5760 9646 5772
rect 9769 5763 9827 5769
rect 9769 5760 9781 5763
rect 9640 5732 9781 5760
rect 9640 5720 9646 5732
rect 9769 5729 9781 5732
rect 9815 5729 9827 5763
rect 9769 5723 9827 5729
rect 2774 5692 2780 5704
rect 2056 5664 2780 5692
rect 2774 5652 2780 5664
rect 2832 5652 2838 5704
rect 3050 5652 3056 5704
rect 3108 5692 3114 5704
rect 4249 5695 4307 5701
rect 3108 5664 3153 5692
rect 3108 5652 3114 5664
rect 4249 5661 4261 5695
rect 4295 5692 4307 5695
rect 4341 5695 4399 5701
rect 4341 5692 4353 5695
rect 4295 5664 4353 5692
rect 4295 5661 4307 5664
rect 4249 5655 4307 5661
rect 4341 5661 4353 5664
rect 4387 5692 4399 5695
rect 6454 5692 6460 5704
rect 4387 5664 6460 5692
rect 4387 5661 4399 5664
rect 4341 5655 4399 5661
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 6937 5695 6995 5701
rect 6937 5661 6949 5695
rect 6983 5692 6995 5695
rect 7466 5692 7472 5704
rect 6983 5664 7472 5692
rect 6983 5661 6995 5664
rect 6937 5655 6995 5661
rect 7466 5652 7472 5664
rect 7524 5652 7530 5704
rect 7926 5652 7932 5704
rect 7984 5692 7990 5704
rect 9858 5692 9864 5704
rect 7984 5664 9864 5692
rect 7984 5652 7990 5664
rect 9858 5652 9864 5664
rect 9916 5652 9922 5704
rect 12066 5652 12072 5704
rect 12124 5692 12130 5704
rect 12621 5695 12679 5701
rect 12621 5692 12633 5695
rect 12124 5664 12633 5692
rect 12124 5652 12130 5664
rect 12621 5661 12633 5664
rect 12667 5661 12679 5695
rect 12621 5655 12679 5661
rect 12710 5652 12716 5704
rect 12768 5692 12774 5704
rect 13173 5695 13231 5701
rect 13173 5692 13185 5695
rect 12768 5664 13185 5692
rect 12768 5652 12774 5664
rect 13173 5661 13185 5664
rect 13219 5661 13231 5695
rect 13280 5692 13308 5800
rect 13372 5772 13400 5868
rect 13722 5856 13728 5908
rect 13780 5896 13786 5908
rect 13817 5899 13875 5905
rect 13817 5896 13829 5899
rect 13780 5868 13829 5896
rect 13780 5856 13786 5868
rect 13817 5865 13829 5868
rect 13863 5896 13875 5899
rect 14369 5899 14427 5905
rect 14369 5896 14381 5899
rect 13863 5868 14381 5896
rect 13863 5865 13875 5868
rect 13817 5859 13875 5865
rect 14369 5865 14381 5868
rect 14415 5865 14427 5899
rect 15378 5896 15384 5908
rect 15339 5868 15384 5896
rect 14369 5859 14427 5865
rect 15378 5856 15384 5868
rect 15436 5856 15442 5908
rect 13354 5720 13360 5772
rect 13412 5760 13418 5772
rect 15102 5760 15108 5772
rect 13412 5732 13505 5760
rect 15063 5732 15108 5760
rect 13412 5720 13418 5732
rect 15102 5720 15108 5732
rect 15160 5720 15166 5772
rect 13633 5695 13691 5701
rect 13633 5692 13645 5695
rect 13280 5664 13645 5692
rect 13173 5655 13231 5661
rect 13633 5661 13645 5664
rect 13679 5692 13691 5695
rect 14182 5692 14188 5704
rect 13679 5664 14188 5692
rect 13679 5661 13691 5664
rect 13633 5655 13691 5661
rect 14182 5652 14188 5664
rect 14240 5652 14246 5704
rect 15562 5692 15568 5704
rect 15523 5664 15568 5692
rect 15562 5652 15568 5664
rect 15620 5652 15626 5704
rect 1578 5584 1584 5636
rect 1636 5624 1642 5636
rect 1946 5624 1952 5636
rect 1636 5596 1952 5624
rect 1636 5584 1642 5596
rect 1946 5584 1952 5596
rect 2004 5624 2010 5636
rect 2004 5596 4108 5624
rect 2004 5584 2010 5596
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 1854 5516 1860 5568
rect 1912 5556 1918 5568
rect 2225 5559 2283 5565
rect 2225 5556 2237 5559
rect 1912 5528 2237 5556
rect 1912 5516 1918 5528
rect 2225 5525 2237 5528
rect 2271 5525 2283 5559
rect 2225 5519 2283 5525
rect 2961 5559 3019 5565
rect 2961 5525 2973 5559
rect 3007 5556 3019 5559
rect 3418 5556 3424 5568
rect 3007 5528 3424 5556
rect 3007 5525 3019 5528
rect 2961 5519 3019 5525
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 3510 5516 3516 5568
rect 3568 5556 3574 5568
rect 3605 5559 3663 5565
rect 3605 5556 3617 5559
rect 3568 5528 3617 5556
rect 3568 5516 3574 5528
rect 3605 5525 3617 5528
rect 3651 5556 3663 5559
rect 3786 5556 3792 5568
rect 3651 5528 3792 5556
rect 3651 5525 3663 5528
rect 3605 5519 3663 5525
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 3878 5516 3884 5568
rect 3936 5556 3942 5568
rect 3973 5559 4031 5565
rect 3973 5556 3985 5559
rect 3936 5528 3985 5556
rect 3936 5516 3942 5528
rect 3973 5525 3985 5528
rect 4019 5525 4031 5559
rect 4080 5556 4108 5596
rect 4154 5584 4160 5636
rect 4212 5624 4218 5636
rect 4586 5627 4644 5633
rect 4586 5624 4598 5627
rect 4212 5596 4598 5624
rect 4212 5584 4218 5596
rect 4586 5593 4598 5596
rect 4632 5593 4644 5627
rect 4586 5587 4644 5593
rect 4706 5584 4712 5636
rect 4764 5624 4770 5636
rect 9306 5624 9312 5636
rect 4764 5596 9312 5624
rect 4764 5584 4770 5596
rect 9306 5584 9312 5596
rect 9364 5584 9370 5636
rect 9766 5584 9772 5636
rect 9824 5624 9830 5636
rect 10014 5627 10072 5633
rect 10014 5624 10026 5627
rect 9824 5596 10026 5624
rect 9824 5584 9830 5596
rect 10014 5593 10026 5596
rect 10060 5593 10072 5627
rect 10014 5587 10072 5593
rect 11790 5584 11796 5636
rect 11848 5624 11854 5636
rect 12158 5624 12164 5636
rect 11848 5596 12164 5624
rect 11848 5584 11854 5596
rect 12158 5584 12164 5596
rect 12216 5584 12222 5636
rect 12354 5627 12412 5633
rect 12354 5593 12366 5627
rect 12400 5593 12412 5627
rect 12354 5587 12412 5593
rect 4430 5556 4436 5568
rect 4080 5528 4436 5556
rect 3973 5519 4031 5525
rect 4430 5516 4436 5528
rect 4488 5516 4494 5568
rect 5721 5559 5779 5565
rect 5721 5525 5733 5559
rect 5767 5556 5779 5559
rect 7098 5556 7104 5568
rect 5767 5528 7104 5556
rect 5767 5525 5779 5528
rect 5721 5519 5779 5525
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 7190 5516 7196 5568
rect 7248 5556 7254 5568
rect 8205 5559 8263 5565
rect 8205 5556 8217 5559
rect 7248 5528 8217 5556
rect 7248 5516 7254 5528
rect 8205 5525 8217 5528
rect 8251 5556 8263 5559
rect 8386 5556 8392 5568
rect 8251 5528 8392 5556
rect 8251 5525 8263 5528
rect 8205 5519 8263 5525
rect 8386 5516 8392 5528
rect 8444 5516 8450 5568
rect 8754 5556 8760 5568
rect 8715 5528 8760 5556
rect 8754 5516 8760 5528
rect 8812 5516 8818 5568
rect 9122 5516 9128 5568
rect 9180 5556 9186 5568
rect 10318 5556 10324 5568
rect 9180 5528 10324 5556
rect 9180 5516 9186 5528
rect 10318 5516 10324 5528
rect 10376 5556 10382 5568
rect 10962 5556 10968 5568
rect 10376 5528 10968 5556
rect 10376 5516 10382 5528
rect 10962 5516 10968 5528
rect 11020 5516 11026 5568
rect 11146 5516 11152 5568
rect 11204 5556 11210 5568
rect 11698 5556 11704 5568
rect 11204 5528 11704 5556
rect 11204 5516 11210 5528
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 11974 5516 11980 5568
rect 12032 5556 12038 5568
rect 12360 5556 12388 5587
rect 13446 5584 13452 5636
rect 13504 5624 13510 5636
rect 14274 5624 14280 5636
rect 13504 5596 14280 5624
rect 13504 5584 13510 5596
rect 14274 5584 14280 5596
rect 14332 5584 14338 5636
rect 14642 5624 14648 5636
rect 14555 5596 14648 5624
rect 14642 5584 14648 5596
rect 14700 5624 14706 5636
rect 15930 5624 15936 5636
rect 14700 5596 15936 5624
rect 14700 5584 14706 5596
rect 15930 5584 15936 5596
rect 15988 5584 15994 5636
rect 12618 5556 12624 5568
rect 12032 5528 12624 5556
rect 12032 5516 12038 5528
rect 12618 5516 12624 5528
rect 12676 5516 12682 5568
rect 12710 5516 12716 5568
rect 12768 5556 12774 5568
rect 12805 5559 12863 5565
rect 12805 5556 12817 5559
rect 12768 5528 12817 5556
rect 12768 5516 12774 5528
rect 12805 5525 12817 5528
rect 12851 5525 12863 5559
rect 13262 5556 13268 5568
rect 13223 5528 13268 5556
rect 12805 5519 12863 5525
rect 13262 5516 13268 5528
rect 13320 5516 13326 5568
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 14093 5559 14151 5565
rect 14093 5556 14105 5559
rect 13872 5528 14105 5556
rect 13872 5516 13878 5528
rect 14093 5525 14105 5528
rect 14139 5525 14151 5559
rect 14734 5556 14740 5568
rect 14695 5528 14740 5556
rect 14093 5519 14151 5525
rect 14734 5516 14740 5528
rect 14792 5516 14798 5568
rect 15013 5559 15071 5565
rect 15013 5525 15025 5559
rect 15059 5556 15071 5559
rect 15378 5556 15384 5568
rect 15059 5528 15384 5556
rect 15059 5525 15071 5528
rect 15013 5519 15071 5525
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 1104 5466 16008 5488
rect 1104 5414 4698 5466
rect 4750 5414 4762 5466
rect 4814 5414 4826 5466
rect 4878 5414 4890 5466
rect 4942 5414 4954 5466
rect 5006 5414 8446 5466
rect 8498 5414 8510 5466
rect 8562 5414 8574 5466
rect 8626 5414 8638 5466
rect 8690 5414 8702 5466
rect 8754 5414 12194 5466
rect 12246 5414 12258 5466
rect 12310 5414 12322 5466
rect 12374 5414 12386 5466
rect 12438 5414 12450 5466
rect 12502 5414 16008 5466
rect 1104 5392 16008 5414
rect 2222 5352 2228 5364
rect 2183 5324 2228 5352
rect 2222 5312 2228 5324
rect 2280 5312 2286 5364
rect 2314 5312 2320 5364
rect 2372 5352 2378 5364
rect 2372 5324 2417 5352
rect 2372 5312 2378 5324
rect 3142 5312 3148 5364
rect 3200 5352 3206 5364
rect 3421 5355 3479 5361
rect 3421 5352 3433 5355
rect 3200 5324 3433 5352
rect 3200 5312 3206 5324
rect 3421 5321 3433 5324
rect 3467 5321 3479 5355
rect 3421 5315 3479 5321
rect 3510 5312 3516 5364
rect 3568 5352 3574 5364
rect 3973 5355 4031 5361
rect 3568 5324 3613 5352
rect 3568 5312 3574 5324
rect 3973 5321 3985 5355
rect 4019 5352 4031 5355
rect 4617 5355 4675 5361
rect 4617 5352 4629 5355
rect 4019 5324 4629 5352
rect 4019 5321 4031 5324
rect 3973 5315 4031 5321
rect 4617 5321 4629 5324
rect 4663 5321 4675 5355
rect 5074 5352 5080 5364
rect 5035 5324 5080 5352
rect 4617 5315 4675 5321
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 5442 5352 5448 5364
rect 5403 5324 5448 5352
rect 5442 5312 5448 5324
rect 5500 5312 5506 5364
rect 6454 5352 6460 5364
rect 6415 5324 6460 5352
rect 6454 5312 6460 5324
rect 6512 5312 6518 5364
rect 6822 5312 6828 5364
rect 6880 5352 6886 5364
rect 7009 5355 7067 5361
rect 7009 5352 7021 5355
rect 6880 5324 7021 5352
rect 6880 5312 6886 5324
rect 7009 5321 7021 5324
rect 7055 5321 7067 5355
rect 8294 5352 8300 5364
rect 8255 5324 8300 5352
rect 7009 5315 7067 5321
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 9861 5355 9919 5361
rect 9861 5321 9873 5355
rect 9907 5352 9919 5355
rect 10042 5352 10048 5364
rect 9907 5324 10048 5352
rect 9907 5321 9919 5324
rect 9861 5315 9919 5321
rect 10042 5312 10048 5324
rect 10100 5312 10106 5364
rect 10226 5312 10232 5364
rect 10284 5352 10290 5364
rect 10778 5352 10784 5364
rect 10284 5324 10784 5352
rect 10284 5312 10290 5324
rect 10778 5312 10784 5324
rect 10836 5312 10842 5364
rect 11149 5355 11207 5361
rect 11149 5321 11161 5355
rect 11195 5352 11207 5355
rect 12066 5352 12072 5364
rect 11195 5324 12072 5352
rect 11195 5321 11207 5324
rect 11149 5315 11207 5321
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 13357 5355 13415 5361
rect 13357 5321 13369 5355
rect 13403 5352 13415 5355
rect 13722 5352 13728 5364
rect 13403 5324 13728 5352
rect 13403 5321 13415 5324
rect 13357 5315 13415 5321
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 14182 5352 14188 5364
rect 14143 5324 14188 5352
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 15102 5312 15108 5364
rect 15160 5352 15166 5364
rect 15197 5355 15255 5361
rect 15197 5352 15209 5355
rect 15160 5324 15209 5352
rect 15160 5312 15166 5324
rect 15197 5321 15209 5324
rect 15243 5321 15255 5355
rect 15197 5315 15255 5321
rect 3053 5287 3111 5293
rect 3053 5253 3065 5287
rect 3099 5284 3111 5287
rect 5166 5284 5172 5296
rect 3099 5256 5172 5284
rect 3099 5253 3111 5256
rect 3053 5247 3111 5253
rect 5166 5244 5172 5256
rect 5224 5244 5230 5296
rect 5534 5244 5540 5296
rect 5592 5284 5598 5296
rect 7190 5284 7196 5296
rect 5592 5256 7196 5284
rect 5592 5244 5598 5256
rect 7190 5244 7196 5256
rect 7248 5244 7254 5296
rect 7300 5256 7880 5284
rect 1854 5216 1860 5228
rect 1815 5188 1860 5216
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 2498 5216 2504 5228
rect 2459 5188 2504 5216
rect 2498 5176 2504 5188
rect 2556 5176 2562 5228
rect 3878 5216 3884 5228
rect 3839 5188 3884 5216
rect 3878 5176 3884 5188
rect 3936 5176 3942 5228
rect 4430 5176 4436 5228
rect 4488 5216 4494 5228
rect 4985 5219 5043 5225
rect 4985 5216 4997 5219
rect 4488 5188 4997 5216
rect 4488 5176 4494 5188
rect 4985 5185 4997 5188
rect 5031 5216 5043 5219
rect 5626 5216 5632 5228
rect 5031 5188 5632 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 5626 5176 5632 5188
rect 5684 5176 5690 5228
rect 5810 5216 5816 5228
rect 5771 5188 5816 5216
rect 5810 5176 5816 5188
rect 5868 5176 5874 5228
rect 6914 5216 6920 5228
rect 6827 5188 6920 5216
rect 6914 5176 6920 5188
rect 6972 5216 6978 5228
rect 7300 5216 7328 5256
rect 6972 5188 7328 5216
rect 6972 5176 6978 5188
rect 7374 5176 7380 5228
rect 7432 5216 7438 5228
rect 7742 5216 7748 5228
rect 7432 5188 7604 5216
rect 7703 5188 7748 5216
rect 7432 5176 7438 5188
rect 1581 5151 1639 5157
rect 1581 5117 1593 5151
rect 1627 5117 1639 5151
rect 1762 5148 1768 5160
rect 1723 5120 1768 5148
rect 1581 5111 1639 5117
rect 1596 5080 1624 5111
rect 1762 5108 1768 5120
rect 1820 5108 1826 5160
rect 2866 5148 2872 5160
rect 2827 5120 2872 5148
rect 2866 5108 2872 5120
rect 2924 5108 2930 5160
rect 2961 5151 3019 5157
rect 2961 5117 2973 5151
rect 3007 5148 3019 5151
rect 3326 5148 3332 5160
rect 3007 5120 3332 5148
rect 3007 5117 3019 5120
rect 2961 5111 3019 5117
rect 3326 5108 3332 5120
rect 3384 5108 3390 5160
rect 4062 5148 4068 5160
rect 4023 5120 4068 5148
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5148 4583 5151
rect 5074 5148 5080 5160
rect 4571 5120 5080 5148
rect 4571 5117 4583 5120
rect 4525 5111 4583 5117
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5148 5319 5151
rect 5718 5148 5724 5160
rect 5307 5120 5724 5148
rect 5307 5117 5319 5120
rect 5261 5111 5319 5117
rect 5718 5108 5724 5120
rect 5776 5108 5782 5160
rect 5902 5148 5908 5160
rect 5863 5120 5908 5148
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 6089 5151 6147 5157
rect 6089 5117 6101 5151
rect 6135 5148 6147 5151
rect 7006 5148 7012 5160
rect 6135 5120 7012 5148
rect 6135 5117 6147 5120
rect 6089 5111 6147 5117
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 7193 5151 7251 5157
rect 7193 5117 7205 5151
rect 7239 5148 7251 5151
rect 7466 5148 7472 5160
rect 7239 5120 7472 5148
rect 7239 5117 7251 5120
rect 7193 5111 7251 5117
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 6178 5080 6184 5092
rect 1596 5052 6184 5080
rect 6178 5040 6184 5052
rect 6236 5040 6242 5092
rect 6270 5040 6276 5092
rect 6328 5080 6334 5092
rect 6328 5052 6776 5080
rect 6328 5040 6334 5052
rect 2774 4972 2780 5024
rect 2832 5012 2838 5024
rect 4062 5012 4068 5024
rect 2832 4984 4068 5012
rect 2832 4972 2838 4984
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 4614 4972 4620 5024
rect 4672 5012 4678 5024
rect 5534 5012 5540 5024
rect 4672 4984 5540 5012
rect 4672 4972 4678 4984
rect 5534 4972 5540 4984
rect 5592 4972 5598 5024
rect 6454 4972 6460 5024
rect 6512 5012 6518 5024
rect 6549 5015 6607 5021
rect 6549 5012 6561 5015
rect 6512 4984 6561 5012
rect 6512 4972 6518 4984
rect 6549 4981 6561 4984
rect 6595 4981 6607 5015
rect 6748 5012 6776 5052
rect 6822 5040 6828 5092
rect 6880 5080 6886 5092
rect 7377 5083 7435 5089
rect 7377 5080 7389 5083
rect 6880 5052 7389 5080
rect 6880 5040 6886 5052
rect 7377 5049 7389 5052
rect 7423 5049 7435 5083
rect 7576 5080 7604 5188
rect 7742 5176 7748 5188
rect 7800 5176 7806 5228
rect 7852 5216 7880 5256
rect 8202 5216 8208 5228
rect 7852 5188 8208 5216
rect 8202 5176 8208 5188
rect 8260 5176 8266 5228
rect 8312 5216 8340 5312
rect 10134 5244 10140 5296
rect 10192 5284 10198 5296
rect 11609 5287 11667 5293
rect 11609 5284 11621 5287
rect 10192 5256 11621 5284
rect 10192 5244 10198 5256
rect 11609 5253 11621 5256
rect 11655 5284 11667 5287
rect 12250 5284 12256 5296
rect 11655 5256 12256 5284
rect 11655 5253 11667 5256
rect 11609 5247 11667 5253
rect 12250 5244 12256 5256
rect 12308 5244 12314 5296
rect 13265 5287 13323 5293
rect 13265 5253 13277 5287
rect 13311 5284 13323 5287
rect 15010 5284 15016 5296
rect 13311 5256 15016 5284
rect 13311 5253 13323 5256
rect 13265 5247 13323 5253
rect 15010 5244 15016 5256
rect 15068 5244 15074 5296
rect 8389 5219 8447 5225
rect 8389 5216 8401 5219
rect 8312 5188 8401 5216
rect 8389 5185 8401 5188
rect 8435 5185 8447 5219
rect 8645 5219 8703 5225
rect 8645 5216 8657 5219
rect 8389 5179 8447 5185
rect 8496 5188 8657 5216
rect 7650 5108 7656 5160
rect 7708 5148 7714 5160
rect 7837 5151 7895 5157
rect 7837 5148 7849 5151
rect 7708 5120 7849 5148
rect 7708 5108 7714 5120
rect 7837 5117 7849 5120
rect 7883 5117 7895 5151
rect 7837 5111 7895 5117
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5117 7987 5151
rect 8496 5148 8524 5188
rect 8645 5185 8657 5188
rect 8691 5185 8703 5219
rect 8645 5179 8703 5185
rect 10229 5219 10287 5225
rect 10229 5185 10241 5219
rect 10275 5216 10287 5219
rect 11514 5216 11520 5228
rect 10275 5188 11520 5216
rect 10275 5185 10287 5188
rect 10229 5179 10287 5185
rect 11514 5176 11520 5188
rect 11572 5176 11578 5228
rect 12437 5219 12495 5225
rect 12437 5185 12449 5219
rect 12483 5216 12495 5219
rect 13170 5216 13176 5228
rect 12483 5188 13176 5216
rect 12483 5185 12495 5188
rect 12437 5179 12495 5185
rect 13170 5176 13176 5188
rect 13228 5176 13234 5228
rect 14090 5216 14096 5228
rect 14051 5188 14096 5216
rect 14090 5176 14096 5188
rect 14148 5216 14154 5228
rect 14829 5219 14887 5225
rect 14829 5216 14841 5219
rect 14148 5188 14841 5216
rect 14148 5176 14154 5188
rect 14829 5185 14841 5188
rect 14875 5216 14887 5219
rect 14918 5216 14924 5228
rect 14875 5188 14924 5216
rect 14875 5185 14887 5188
rect 14829 5179 14887 5185
rect 14918 5176 14924 5188
rect 14976 5176 14982 5228
rect 15470 5216 15476 5228
rect 15431 5188 15476 5216
rect 15470 5176 15476 5188
rect 15528 5176 15534 5228
rect 7929 5111 7987 5117
rect 8404 5120 8524 5148
rect 10321 5151 10379 5157
rect 7944 5080 7972 5111
rect 7576 5052 7972 5080
rect 7377 5043 7435 5049
rect 7006 5012 7012 5024
rect 6748 4984 7012 5012
rect 6549 4975 6607 4981
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 7098 4972 7104 5024
rect 7156 5012 7162 5024
rect 7834 5012 7840 5024
rect 7156 4984 7840 5012
rect 7156 4972 7162 4984
rect 7834 4972 7840 4984
rect 7892 5012 7898 5024
rect 8404 5012 8432 5120
rect 10321 5117 10333 5151
rect 10367 5117 10379 5151
rect 10321 5111 10379 5117
rect 10413 5151 10471 5157
rect 10413 5117 10425 5151
rect 10459 5117 10471 5151
rect 10413 5111 10471 5117
rect 9398 5040 9404 5092
rect 9456 5080 9462 5092
rect 9456 5052 9996 5080
rect 9456 5040 9462 5052
rect 7892 4984 8432 5012
rect 9769 5015 9827 5021
rect 7892 4972 7898 4984
rect 9769 4981 9781 5015
rect 9815 5012 9827 5015
rect 9858 5012 9864 5024
rect 9815 4984 9864 5012
rect 9815 4981 9827 4984
rect 9769 4975 9827 4981
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 9968 5012 9996 5052
rect 10226 5040 10232 5092
rect 10284 5080 10290 5092
rect 10336 5080 10364 5111
rect 10284 5052 10364 5080
rect 10284 5040 10290 5052
rect 10428 5012 10456 5111
rect 11238 5108 11244 5160
rect 11296 5108 11302 5160
rect 11333 5151 11391 5157
rect 11333 5117 11345 5151
rect 11379 5148 11391 5151
rect 11422 5148 11428 5160
rect 11379 5120 11428 5148
rect 11379 5117 11391 5120
rect 11333 5111 11391 5117
rect 11422 5108 11428 5120
rect 11480 5108 11486 5160
rect 11977 5151 12035 5157
rect 11977 5117 11989 5151
rect 12023 5148 12035 5151
rect 12250 5148 12256 5160
rect 12023 5120 12256 5148
rect 12023 5117 12035 5120
rect 11977 5111 12035 5117
rect 12250 5108 12256 5120
rect 12308 5108 12314 5160
rect 12526 5148 12532 5160
rect 12487 5120 12532 5148
rect 12526 5108 12532 5120
rect 12584 5108 12590 5160
rect 12621 5151 12679 5157
rect 12621 5117 12633 5151
rect 12667 5117 12679 5151
rect 13446 5148 13452 5160
rect 13407 5120 13452 5148
rect 12621 5111 12679 5117
rect 11256 5080 11284 5108
rect 12636 5080 12664 5111
rect 13446 5108 13452 5120
rect 13504 5108 13510 5160
rect 14274 5148 14280 5160
rect 14235 5120 14280 5148
rect 14274 5108 14280 5120
rect 14332 5108 14338 5160
rect 14458 5108 14464 5160
rect 14516 5148 14522 5160
rect 14553 5151 14611 5157
rect 14553 5148 14565 5151
rect 14516 5120 14565 5148
rect 14516 5108 14522 5120
rect 14553 5117 14565 5120
rect 14599 5117 14611 5151
rect 14553 5111 14611 5117
rect 11256 5052 12664 5080
rect 14292 5080 14320 5108
rect 14642 5080 14648 5092
rect 14292 5052 14648 5080
rect 14642 5040 14648 5052
rect 14700 5040 14706 5092
rect 10686 5012 10692 5024
rect 9968 4984 10456 5012
rect 10647 4984 10692 5012
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 10870 5012 10876 5024
rect 10831 4984 10876 5012
rect 10870 4972 10876 4984
rect 10928 4972 10934 5024
rect 12066 5012 12072 5024
rect 12027 4984 12072 5012
rect 12066 4972 12072 4984
rect 12124 4972 12130 5024
rect 12158 4972 12164 5024
rect 12216 5012 12222 5024
rect 12897 5015 12955 5021
rect 12897 5012 12909 5015
rect 12216 4984 12909 5012
rect 12216 4972 12222 4984
rect 12897 4981 12909 4984
rect 12943 4981 12955 5015
rect 12897 4975 12955 4981
rect 13630 4972 13636 5024
rect 13688 5012 13694 5024
rect 13725 5015 13783 5021
rect 13725 5012 13737 5015
rect 13688 4984 13737 5012
rect 13688 4972 13694 4984
rect 13725 4981 13737 4984
rect 13771 4981 13783 5015
rect 15102 5012 15108 5024
rect 15063 4984 15108 5012
rect 13725 4975 13783 4981
rect 15102 4972 15108 4984
rect 15160 4972 15166 5024
rect 15657 5015 15715 5021
rect 15657 4981 15669 5015
rect 15703 5012 15715 5015
rect 15930 5012 15936 5024
rect 15703 4984 15936 5012
rect 15703 4981 15715 4984
rect 15657 4975 15715 4981
rect 15930 4972 15936 4984
rect 15988 4972 15994 5024
rect 1104 4922 16008 4944
rect 1104 4870 2824 4922
rect 2876 4870 2888 4922
rect 2940 4870 2952 4922
rect 3004 4870 3016 4922
rect 3068 4870 3080 4922
rect 3132 4870 6572 4922
rect 6624 4870 6636 4922
rect 6688 4870 6700 4922
rect 6752 4870 6764 4922
rect 6816 4870 6828 4922
rect 6880 4870 10320 4922
rect 10372 4870 10384 4922
rect 10436 4870 10448 4922
rect 10500 4870 10512 4922
rect 10564 4870 10576 4922
rect 10628 4870 14068 4922
rect 14120 4870 14132 4922
rect 14184 4870 14196 4922
rect 14248 4870 14260 4922
rect 14312 4870 14324 4922
rect 14376 4870 16008 4922
rect 1104 4848 16008 4870
rect 1762 4768 1768 4820
rect 1820 4808 1826 4820
rect 1857 4811 1915 4817
rect 1857 4808 1869 4811
rect 1820 4780 1869 4808
rect 1820 4768 1826 4780
rect 1857 4777 1869 4780
rect 1903 4777 1915 4811
rect 1857 4771 1915 4777
rect 3973 4811 4031 4817
rect 3973 4777 3985 4811
rect 4019 4808 4031 4811
rect 4154 4808 4160 4820
rect 4019 4780 4160 4808
rect 4019 4777 4031 4780
rect 3973 4771 4031 4777
rect 4154 4768 4160 4780
rect 4212 4768 4218 4820
rect 5626 4808 5632 4820
rect 4264 4780 5488 4808
rect 5587 4780 5632 4808
rect 2130 4700 2136 4752
rect 2188 4740 2194 4752
rect 2869 4743 2927 4749
rect 2869 4740 2881 4743
rect 2188 4712 2881 4740
rect 2188 4700 2194 4712
rect 2869 4709 2881 4712
rect 2915 4709 2927 4743
rect 2869 4703 2927 4709
rect 3878 4700 3884 4752
rect 3936 4740 3942 4752
rect 4264 4740 4292 4780
rect 3936 4712 4292 4740
rect 4341 4743 4399 4749
rect 3936 4700 3942 4712
rect 4341 4709 4353 4743
rect 4387 4740 4399 4743
rect 5460 4740 5488 4780
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 5902 4768 5908 4820
rect 5960 4808 5966 4820
rect 6181 4811 6239 4817
rect 6181 4808 6193 4811
rect 5960 4780 6193 4808
rect 5960 4768 5966 4780
rect 6181 4777 6193 4780
rect 6227 4777 6239 4811
rect 6181 4771 6239 4777
rect 6288 4780 6500 4808
rect 6288 4740 6316 4780
rect 4387 4712 5405 4740
rect 5460 4712 6316 4740
rect 6472 4740 6500 4780
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 8941 4811 8999 4817
rect 8941 4808 8953 4811
rect 7708 4780 8953 4808
rect 7708 4768 7714 4780
rect 8941 4777 8953 4780
rect 8987 4777 8999 4811
rect 8941 4771 8999 4777
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 9493 4811 9551 4817
rect 9493 4808 9505 4811
rect 9272 4780 9505 4808
rect 9272 4768 9278 4780
rect 9493 4777 9505 4780
rect 9539 4777 9551 4811
rect 9493 4771 9551 4777
rect 10226 4768 10232 4820
rect 10284 4808 10290 4820
rect 10321 4811 10379 4817
rect 10321 4808 10333 4811
rect 10284 4780 10333 4808
rect 10284 4768 10290 4780
rect 10321 4777 10333 4780
rect 10367 4777 10379 4811
rect 10321 4771 10379 4777
rect 10410 4768 10416 4820
rect 10468 4808 10474 4820
rect 10778 4808 10784 4820
rect 10468 4780 10784 4808
rect 10468 4768 10474 4780
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 10962 4808 10968 4820
rect 10923 4780 10968 4808
rect 10962 4768 10968 4780
rect 11020 4768 11026 4820
rect 11514 4808 11520 4820
rect 11475 4780 11520 4808
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 14826 4768 14832 4820
rect 14884 4808 14890 4820
rect 14921 4811 14979 4817
rect 14921 4808 14933 4811
rect 14884 4780 14933 4808
rect 14884 4768 14890 4780
rect 14921 4777 14933 4780
rect 14967 4777 14979 4811
rect 14921 4771 14979 4777
rect 8573 4743 8631 4749
rect 6472 4712 7880 4740
rect 4387 4709 4399 4712
rect 4341 4703 4399 4709
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4672 2559 4675
rect 2590 4672 2596 4684
rect 2547 4644 2596 4672
rect 2547 4641 2559 4644
rect 2501 4635 2559 4641
rect 2590 4632 2596 4644
rect 2648 4632 2654 4684
rect 2682 4632 2688 4684
rect 2740 4672 2746 4684
rect 2740 4632 2774 4672
rect 3234 4632 3240 4684
rect 3292 4672 3298 4684
rect 3421 4675 3479 4681
rect 3421 4672 3433 4675
rect 3292 4644 3433 4672
rect 3292 4632 3298 4644
rect 3421 4641 3433 4644
rect 3467 4672 3479 4675
rect 4985 4675 5043 4681
rect 4985 4672 4997 4675
rect 3467 4644 4997 4672
rect 3467 4641 3479 4644
rect 3421 4635 3479 4641
rect 4985 4641 4997 4644
rect 5031 4641 5043 4675
rect 5377 4672 5405 4712
rect 5377 4644 5580 4672
rect 4985 4635 5043 4641
rect 1670 4604 1676 4616
rect 1631 4576 1676 4604
rect 1670 4564 1676 4576
rect 1728 4564 1734 4616
rect 2746 4604 2774 4632
rect 3789 4607 3847 4613
rect 3789 4604 3801 4607
rect 2746 4576 3801 4604
rect 3789 4573 3801 4576
rect 3835 4573 3847 4607
rect 4154 4604 4160 4616
rect 4067 4576 4160 4604
rect 3789 4567 3847 4573
rect 4154 4564 4160 4576
rect 4212 4604 4218 4616
rect 5442 4604 5448 4616
rect 4212 4576 5448 4604
rect 4212 4564 4218 4576
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 2225 4539 2283 4545
rect 2225 4505 2237 4539
rect 2271 4536 2283 4539
rect 5552 4536 5580 4644
rect 5902 4632 5908 4684
rect 5960 4672 5966 4684
rect 6362 4672 6368 4684
rect 5960 4644 6368 4672
rect 5960 4632 5966 4644
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 6454 4632 6460 4684
rect 6512 4672 6518 4684
rect 6641 4675 6699 4681
rect 6641 4672 6653 4675
rect 6512 4644 6653 4672
rect 6512 4632 6518 4644
rect 6641 4641 6653 4644
rect 6687 4641 6699 4675
rect 6641 4635 6699 4641
rect 6825 4675 6883 4681
rect 6825 4641 6837 4675
rect 6871 4641 6883 4675
rect 7098 4672 7104 4684
rect 7059 4644 7104 4672
rect 6825 4635 6883 4641
rect 6086 4604 6092 4616
rect 5999 4576 6092 4604
rect 6086 4564 6092 4576
rect 6144 4604 6150 4616
rect 6840 4604 6868 4635
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 7190 4632 7196 4684
rect 7248 4672 7254 4684
rect 7285 4675 7343 4681
rect 7285 4672 7297 4675
rect 7248 4644 7297 4672
rect 7248 4632 7254 4644
rect 7285 4641 7297 4644
rect 7331 4672 7343 4675
rect 7742 4672 7748 4684
rect 7331 4644 7748 4672
rect 7331 4641 7343 4644
rect 7285 4635 7343 4641
rect 7742 4632 7748 4644
rect 7800 4632 7806 4684
rect 7006 4604 7012 4616
rect 6144 4576 6684 4604
rect 6840 4576 7012 4604
rect 6144 4564 6150 4576
rect 6656 4548 6684 4576
rect 7006 4564 7012 4576
rect 7064 4564 7070 4616
rect 7852 4604 7880 4712
rect 8036 4712 8340 4740
rect 8036 4681 8064 4712
rect 8021 4675 8079 4681
rect 8021 4641 8033 4675
rect 8067 4641 8079 4675
rect 8312 4672 8340 4712
rect 8573 4709 8585 4743
rect 8619 4740 8631 4743
rect 9398 4740 9404 4752
rect 8619 4712 9404 4740
rect 8619 4709 8631 4712
rect 8573 4703 8631 4709
rect 9398 4700 9404 4712
rect 9456 4700 9462 4752
rect 9582 4700 9588 4752
rect 9640 4740 9646 4752
rect 11241 4743 11299 4749
rect 11241 4740 11253 4743
rect 9640 4712 11253 4740
rect 9640 4700 9646 4712
rect 11241 4709 11253 4712
rect 11287 4709 11299 4743
rect 11241 4703 11299 4709
rect 11330 4700 11336 4752
rect 11388 4740 11394 4752
rect 13446 4740 13452 4752
rect 11388 4712 13452 4740
rect 11388 4700 11394 4712
rect 8938 4672 8944 4684
rect 8312 4644 8944 4672
rect 8021 4635 8079 4641
rect 8938 4632 8944 4644
rect 8996 4632 9002 4684
rect 9674 4672 9680 4684
rect 9048 4644 9352 4672
rect 9635 4644 9680 4672
rect 9048 4604 9076 4644
rect 7852 4576 9076 4604
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4604 9183 4607
rect 9324 4604 9352 4644
rect 9674 4632 9680 4644
rect 9732 4672 9738 4684
rect 12069 4675 12127 4681
rect 12069 4672 12081 4675
rect 9732 4644 12081 4672
rect 9732 4632 9738 4644
rect 12069 4641 12081 4644
rect 12115 4641 12127 4675
rect 12802 4672 12808 4684
rect 12069 4635 12127 4641
rect 12176 4644 12808 4672
rect 10226 4604 10232 4616
rect 9171 4576 9205 4604
rect 9324 4576 10232 4604
rect 9171 4573 9183 4576
rect 9125 4567 9183 4573
rect 6178 4536 6184 4548
rect 2271 4508 4476 4536
rect 5552 4508 6184 4536
rect 2271 4505 2283 4508
rect 2225 4499 2283 4505
rect 1486 4468 1492 4480
rect 1447 4440 1492 4468
rect 1486 4428 1492 4440
rect 1544 4428 1550 4480
rect 2314 4468 2320 4480
rect 2275 4440 2320 4468
rect 2314 4428 2320 4440
rect 2372 4428 2378 4480
rect 2498 4428 2504 4480
rect 2556 4468 2562 4480
rect 2682 4468 2688 4480
rect 2556 4440 2688 4468
rect 2556 4428 2562 4440
rect 2682 4428 2688 4440
rect 2740 4428 2746 4480
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 2832 4440 2877 4468
rect 2832 4428 2838 4440
rect 3050 4428 3056 4480
rect 3108 4468 3114 4480
rect 3237 4471 3295 4477
rect 3237 4468 3249 4471
rect 3108 4440 3249 4468
rect 3108 4428 3114 4440
rect 3237 4437 3249 4440
rect 3283 4437 3295 4471
rect 3237 4431 3295 4437
rect 3329 4471 3387 4477
rect 3329 4437 3341 4471
rect 3375 4468 3387 4471
rect 3418 4468 3424 4480
rect 3375 4440 3424 4468
rect 3375 4437 3387 4440
rect 3329 4431 3387 4437
rect 3418 4428 3424 4440
rect 3476 4468 3482 4480
rect 3786 4468 3792 4480
rect 3476 4440 3792 4468
rect 3476 4428 3482 4440
rect 3786 4428 3792 4440
rect 3844 4428 3850 4480
rect 4448 4477 4476 4508
rect 6178 4496 6184 4508
rect 6236 4496 6242 4548
rect 6638 4496 6644 4548
rect 6696 4496 6702 4548
rect 7282 4496 7288 4548
rect 7340 4536 7346 4548
rect 7377 4539 7435 4545
rect 7377 4536 7389 4539
rect 7340 4508 7389 4536
rect 7340 4496 7346 4508
rect 7377 4505 7389 4508
rect 7423 4536 7435 4539
rect 8665 4539 8723 4545
rect 8665 4536 8677 4539
rect 7423 4508 8677 4536
rect 7423 4505 7435 4508
rect 7377 4499 7435 4505
rect 8665 4505 8677 4508
rect 8711 4505 8723 4539
rect 8665 4499 8723 4505
rect 8846 4496 8852 4548
rect 8904 4536 8910 4548
rect 9140 4536 9168 4567
rect 10226 4564 10232 4576
rect 10284 4604 10290 4616
rect 10413 4607 10471 4613
rect 10413 4604 10425 4607
rect 10284 4576 10425 4604
rect 10284 4564 10290 4576
rect 10413 4573 10425 4576
rect 10459 4573 10471 4607
rect 10413 4567 10471 4573
rect 10689 4607 10747 4613
rect 10689 4573 10701 4607
rect 10735 4604 10747 4607
rect 10962 4604 10968 4616
rect 10735 4576 10968 4604
rect 10735 4573 10747 4576
rect 10689 4567 10747 4573
rect 10962 4564 10968 4576
rect 11020 4564 11026 4616
rect 11425 4607 11483 4613
rect 11425 4573 11437 4607
rect 11471 4604 11483 4607
rect 12176 4604 12204 4644
rect 12802 4632 12808 4644
rect 12860 4632 12866 4684
rect 12912 4681 12940 4712
rect 13446 4700 13452 4712
rect 13504 4700 13510 4752
rect 12897 4675 12955 4681
rect 12897 4641 12909 4675
rect 12943 4641 12955 4675
rect 13630 4672 13636 4684
rect 13591 4644 13636 4672
rect 12897 4635 12955 4641
rect 13630 4632 13636 4644
rect 13688 4632 13694 4684
rect 13725 4675 13783 4681
rect 13725 4641 13737 4675
rect 13771 4641 13783 4675
rect 14642 4672 14648 4684
rect 14603 4644 14648 4672
rect 13725 4635 13783 4641
rect 11471 4576 12204 4604
rect 11471 4573 11483 4576
rect 11425 4567 11483 4573
rect 12250 4564 12256 4616
rect 12308 4604 12314 4616
rect 12713 4607 12771 4613
rect 12713 4604 12725 4607
rect 12308 4576 12725 4604
rect 12308 4564 12314 4576
rect 12713 4573 12725 4576
rect 12759 4573 12771 4607
rect 13740 4604 13768 4635
rect 14642 4632 14648 4644
rect 14700 4632 14706 4684
rect 14458 4604 14464 4616
rect 12713 4567 12771 4573
rect 13464 4576 13768 4604
rect 14419 4576 14464 4604
rect 9217 4539 9275 4545
rect 9217 4536 9229 4539
rect 8904 4508 9229 4536
rect 8904 4496 8910 4508
rect 9217 4505 9229 4508
rect 9263 4505 9275 4539
rect 10318 4536 10324 4548
rect 9217 4499 9275 4505
rect 9876 4508 10324 4536
rect 4433 4471 4491 4477
rect 4433 4437 4445 4471
rect 4479 4437 4491 4471
rect 4798 4468 4804 4480
rect 4759 4440 4804 4468
rect 4433 4431 4491 4437
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 4893 4471 4951 4477
rect 4893 4437 4905 4471
rect 4939 4468 4951 4471
rect 5074 4468 5080 4480
rect 4939 4440 5080 4468
rect 4939 4437 4951 4440
rect 4893 4431 4951 4437
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 5445 4471 5503 4477
rect 5445 4437 5457 4471
rect 5491 4468 5503 4471
rect 5534 4468 5540 4480
rect 5491 4440 5540 4468
rect 5491 4437 5503 4440
rect 5445 4431 5503 4437
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 5905 4471 5963 4477
rect 5905 4437 5917 4471
rect 5951 4468 5963 4471
rect 6362 4468 6368 4480
rect 5951 4440 6368 4468
rect 5951 4437 5963 4440
rect 5905 4431 5963 4437
rect 6362 4428 6368 4440
rect 6420 4428 6426 4480
rect 6454 4428 6460 4480
rect 6512 4468 6518 4480
rect 6549 4471 6607 4477
rect 6549 4468 6561 4471
rect 6512 4440 6561 4468
rect 6512 4428 6518 4440
rect 6549 4437 6561 4440
rect 6595 4437 6607 4471
rect 7742 4468 7748 4480
rect 7703 4440 7748 4468
rect 6549 4431 6607 4437
rect 7742 4428 7748 4440
rect 7800 4428 7806 4480
rect 8018 4428 8024 4480
rect 8076 4468 8082 4480
rect 8113 4471 8171 4477
rect 8113 4468 8125 4471
rect 8076 4440 8125 4468
rect 8076 4428 8082 4440
rect 8113 4437 8125 4440
rect 8159 4437 8171 4471
rect 8113 4431 8171 4437
rect 8205 4471 8263 4477
rect 8205 4437 8217 4471
rect 8251 4468 8263 4471
rect 8294 4468 8300 4480
rect 8251 4440 8300 4468
rect 8251 4437 8263 4440
rect 8205 4431 8263 4437
rect 8294 4428 8300 4440
rect 8352 4428 8358 4480
rect 9876 4477 9904 4508
rect 10318 4496 10324 4508
rect 10376 4496 10382 4548
rect 11885 4539 11943 4545
rect 11885 4505 11897 4539
rect 11931 4536 11943 4539
rect 11931 4508 12388 4536
rect 11931 4505 11943 4508
rect 11885 4499 11943 4505
rect 9861 4471 9919 4477
rect 9861 4437 9873 4471
rect 9907 4437 9919 4471
rect 9861 4431 9919 4437
rect 9950 4428 9956 4480
rect 10008 4468 10014 4480
rect 10008 4440 10053 4468
rect 10008 4428 10014 4440
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 11514 4468 11520 4480
rect 11112 4440 11520 4468
rect 11112 4428 11118 4440
rect 11514 4428 11520 4440
rect 11572 4428 11578 4480
rect 11977 4471 12035 4477
rect 11977 4437 11989 4471
rect 12023 4468 12035 4471
rect 12158 4468 12164 4480
rect 12023 4440 12164 4468
rect 12023 4437 12035 4440
rect 11977 4431 12035 4437
rect 12158 4428 12164 4440
rect 12216 4428 12222 4480
rect 12360 4477 12388 4508
rect 12434 4496 12440 4548
rect 12492 4536 12498 4548
rect 12618 4536 12624 4548
rect 12492 4508 12624 4536
rect 12492 4496 12498 4508
rect 12618 4496 12624 4508
rect 12676 4536 12682 4548
rect 13464 4536 13492 4576
rect 14458 4564 14464 4576
rect 14516 4564 14522 4616
rect 15102 4604 15108 4616
rect 15063 4576 15108 4604
rect 15102 4564 15108 4576
rect 15160 4564 15166 4616
rect 15378 4564 15384 4616
rect 15436 4604 15442 4616
rect 15473 4607 15531 4613
rect 15473 4604 15485 4607
rect 15436 4576 15485 4604
rect 15436 4564 15442 4576
rect 15473 4573 15485 4576
rect 15519 4573 15531 4607
rect 15473 4567 15531 4573
rect 12676 4508 13492 4536
rect 13541 4539 13599 4545
rect 12676 4496 12682 4508
rect 13541 4505 13553 4539
rect 13587 4536 13599 4539
rect 13587 4508 14136 4536
rect 13587 4505 13599 4508
rect 13541 4499 13599 4505
rect 12345 4471 12403 4477
rect 12345 4437 12357 4471
rect 12391 4437 12403 4471
rect 12802 4468 12808 4480
rect 12763 4440 12808 4468
rect 12345 4431 12403 4437
rect 12802 4428 12808 4440
rect 12860 4428 12866 4480
rect 13170 4468 13176 4480
rect 13131 4440 13176 4468
rect 13170 4428 13176 4440
rect 13228 4428 13234 4480
rect 14108 4477 14136 4508
rect 14093 4471 14151 4477
rect 14093 4437 14105 4471
rect 14139 4437 14151 4471
rect 14093 4431 14151 4437
rect 14458 4428 14464 4480
rect 14516 4468 14522 4480
rect 14553 4471 14611 4477
rect 14553 4468 14565 4471
rect 14516 4440 14565 4468
rect 14516 4428 14522 4440
rect 14553 4437 14565 4440
rect 14599 4437 14611 4471
rect 15378 4468 15384 4480
rect 15339 4440 15384 4468
rect 14553 4431 14611 4437
rect 15378 4428 15384 4440
rect 15436 4468 15442 4480
rect 16022 4468 16028 4480
rect 15436 4440 16028 4468
rect 15436 4428 15442 4440
rect 16022 4428 16028 4440
rect 16080 4428 16086 4480
rect 1104 4378 16008 4400
rect 1104 4326 4698 4378
rect 4750 4326 4762 4378
rect 4814 4326 4826 4378
rect 4878 4326 4890 4378
rect 4942 4326 4954 4378
rect 5006 4326 8446 4378
rect 8498 4326 8510 4378
rect 8562 4326 8574 4378
rect 8626 4326 8638 4378
rect 8690 4326 8702 4378
rect 8754 4326 12194 4378
rect 12246 4326 12258 4378
rect 12310 4326 12322 4378
rect 12374 4326 12386 4378
rect 12438 4326 12450 4378
rect 12502 4326 16008 4378
rect 1104 4304 16008 4326
rect 1673 4267 1731 4273
rect 1673 4233 1685 4267
rect 1719 4264 1731 4267
rect 1854 4264 1860 4276
rect 1719 4236 1860 4264
rect 1719 4233 1731 4236
rect 1673 4227 1731 4233
rect 1854 4224 1860 4236
rect 1912 4224 1918 4276
rect 2038 4264 2044 4276
rect 1999 4236 2044 4264
rect 2038 4224 2044 4236
rect 2096 4224 2102 4276
rect 2961 4267 3019 4273
rect 2961 4233 2973 4267
rect 3007 4264 3019 4267
rect 3142 4264 3148 4276
rect 3007 4236 3148 4264
rect 3007 4233 3019 4236
rect 2961 4227 3019 4233
rect 3142 4224 3148 4236
rect 3200 4224 3206 4276
rect 3326 4264 3332 4276
rect 3287 4236 3332 4264
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 3694 4224 3700 4276
rect 3752 4264 3758 4276
rect 3789 4267 3847 4273
rect 3789 4264 3801 4267
rect 3752 4236 3801 4264
rect 3752 4224 3758 4236
rect 3789 4233 3801 4236
rect 3835 4233 3847 4267
rect 5166 4264 5172 4276
rect 5127 4236 5172 4264
rect 3789 4227 3847 4233
rect 5166 4224 5172 4236
rect 5224 4224 5230 4276
rect 5534 4264 5540 4276
rect 5495 4236 5540 4264
rect 5534 4224 5540 4236
rect 5592 4224 5598 4276
rect 5718 4224 5724 4276
rect 5776 4264 5782 4276
rect 5997 4267 6055 4273
rect 5997 4264 6009 4267
rect 5776 4236 6009 4264
rect 5776 4224 5782 4236
rect 5997 4233 6009 4236
rect 6043 4233 6055 4267
rect 5997 4227 6055 4233
rect 6178 4224 6184 4276
rect 6236 4264 6242 4276
rect 7006 4264 7012 4276
rect 6236 4236 7012 4264
rect 6236 4224 6242 4236
rect 7006 4224 7012 4236
rect 7064 4224 7070 4276
rect 7742 4224 7748 4276
rect 7800 4264 7806 4276
rect 7929 4267 7987 4273
rect 7929 4264 7941 4267
rect 7800 4236 7941 4264
rect 7800 4224 7806 4236
rect 7929 4233 7941 4236
rect 7975 4233 7987 4267
rect 7929 4227 7987 4233
rect 8021 4267 8079 4273
rect 8021 4233 8033 4267
rect 8067 4233 8079 4267
rect 8021 4227 8079 4233
rect 4062 4196 4068 4208
rect 3252 4168 4068 4196
rect 1578 4128 1584 4140
rect 1539 4100 1584 4128
rect 1578 4088 1584 4100
rect 1636 4088 1642 4140
rect 2130 4088 2136 4140
rect 2188 4128 2194 4140
rect 2188 4100 2233 4128
rect 2188 4088 2194 4100
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 2869 4131 2927 4137
rect 2869 4128 2881 4131
rect 2832 4100 2881 4128
rect 2832 4088 2838 4100
rect 2869 4097 2881 4100
rect 2915 4097 2927 4131
rect 2869 4091 2927 4097
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 2590 4060 2596 4072
rect 2363 4032 2596 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 2590 4020 2596 4032
rect 2648 4020 2654 4072
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4060 2743 4063
rect 3252 4060 3280 4168
rect 4062 4156 4068 4168
rect 4120 4196 4126 4208
rect 4120 4168 4660 4196
rect 4120 4156 4126 4168
rect 4338 4128 4344 4140
rect 4080 4100 4344 4128
rect 4080 4069 4108 4100
rect 4338 4088 4344 4100
rect 4396 4088 4402 4140
rect 4522 4128 4528 4140
rect 4483 4100 4528 4128
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 2731 4032 3280 4060
rect 3881 4063 3939 4069
rect 2731 4029 2743 4032
rect 2685 4023 2743 4029
rect 3881 4029 3893 4063
rect 3927 4029 3939 4063
rect 3881 4023 3939 4029
rect 4065 4063 4123 4069
rect 4065 4029 4077 4063
rect 4111 4029 4123 4063
rect 4065 4023 4123 4029
rect 4249 4063 4307 4069
rect 4249 4029 4261 4063
rect 4295 4029 4307 4063
rect 4632 4060 4660 4168
rect 7374 4156 7380 4208
rect 7432 4196 7438 4208
rect 8036 4196 8064 4227
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 8389 4267 8447 4273
rect 8389 4264 8401 4267
rect 8352 4236 8401 4264
rect 8352 4224 8358 4236
rect 8389 4233 8401 4236
rect 8435 4233 8447 4267
rect 9398 4264 9404 4276
rect 9359 4236 9404 4264
rect 8389 4227 8447 4233
rect 9398 4224 9404 4236
rect 9456 4224 9462 4276
rect 10318 4264 10324 4276
rect 10279 4236 10324 4264
rect 10318 4224 10324 4236
rect 10376 4224 10382 4276
rect 10689 4267 10747 4273
rect 10689 4233 10701 4267
rect 10735 4264 10747 4267
rect 11054 4264 11060 4276
rect 10735 4236 11060 4264
rect 10735 4233 10747 4236
rect 10689 4227 10747 4233
rect 11054 4224 11060 4236
rect 11112 4224 11118 4276
rect 11149 4267 11207 4273
rect 11149 4233 11161 4267
rect 11195 4233 11207 4267
rect 11514 4264 11520 4276
rect 11475 4236 11520 4264
rect 11149 4227 11207 4233
rect 9582 4196 9588 4208
rect 7432 4168 8064 4196
rect 8312 4168 9588 4196
rect 7432 4156 7438 4168
rect 7760 4140 7788 4168
rect 8312 4140 8340 4168
rect 9582 4156 9588 4168
rect 9640 4156 9646 4208
rect 10226 4196 10232 4208
rect 9968 4168 10232 4196
rect 5626 4128 5632 4140
rect 5587 4100 5632 4128
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 5994 4128 6000 4140
rect 5736 4100 6000 4128
rect 5736 4069 5764 4100
rect 5994 4088 6000 4100
rect 6052 4088 6058 4140
rect 6178 4088 6184 4140
rect 6236 4128 6242 4140
rect 6236 4100 6281 4128
rect 6236 4088 6242 4100
rect 6362 4088 6368 4140
rect 6420 4128 6426 4140
rect 6457 4131 6515 4137
rect 6457 4128 6469 4131
rect 6420 4100 6469 4128
rect 6420 4088 6426 4100
rect 6457 4097 6469 4100
rect 6503 4097 6515 4131
rect 6457 4091 6515 4097
rect 6638 4088 6644 4140
rect 6696 4128 6702 4140
rect 7009 4131 7067 4137
rect 7009 4128 7021 4131
rect 6696 4100 7021 4128
rect 6696 4088 6702 4100
rect 7009 4097 7021 4100
rect 7055 4097 7067 4131
rect 7558 4128 7564 4140
rect 7519 4100 7564 4128
rect 7009 4091 7067 4097
rect 7558 4088 7564 4100
rect 7616 4088 7622 4140
rect 7742 4088 7748 4140
rect 7800 4088 7806 4140
rect 8294 4088 8300 4140
rect 8352 4088 8358 4140
rect 8754 4128 8760 4140
rect 8715 4100 8760 4128
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 8849 4131 8907 4137
rect 8849 4097 8861 4131
rect 8895 4128 8907 4131
rect 9214 4128 9220 4140
rect 8895 4100 9220 4128
rect 8895 4097 8907 4100
rect 8849 4091 8907 4097
rect 9214 4088 9220 4100
rect 9272 4088 9278 4140
rect 9490 4128 9496 4140
rect 9451 4100 9496 4128
rect 9490 4088 9496 4100
rect 9548 4088 9554 4140
rect 9674 4088 9680 4140
rect 9732 4128 9738 4140
rect 9858 4128 9864 4140
rect 9732 4100 9864 4128
rect 9732 4088 9738 4100
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 9968 4137 9996 4168
rect 10226 4156 10232 4168
rect 10284 4156 10290 4208
rect 11164 4196 11192 4227
rect 11514 4224 11520 4236
rect 11572 4224 11578 4276
rect 11885 4267 11943 4273
rect 11885 4233 11897 4267
rect 11931 4264 11943 4267
rect 11974 4264 11980 4276
rect 11931 4236 11980 4264
rect 11931 4233 11943 4236
rect 11885 4227 11943 4233
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 12434 4224 12440 4276
rect 12492 4264 12498 4276
rect 12894 4264 12900 4276
rect 12492 4236 12900 4264
rect 12492 4224 12498 4236
rect 12894 4224 12900 4236
rect 12952 4264 12958 4276
rect 13081 4267 13139 4273
rect 13081 4264 13093 4267
rect 12952 4236 13093 4264
rect 12952 4224 12958 4236
rect 13081 4233 13093 4236
rect 13127 4233 13139 4267
rect 13081 4227 13139 4233
rect 13814 4224 13820 4276
rect 13872 4264 13878 4276
rect 13909 4267 13967 4273
rect 13909 4264 13921 4267
rect 13872 4236 13921 4264
rect 13872 4224 13878 4236
rect 13909 4233 13921 4236
rect 13955 4264 13967 4267
rect 14458 4264 14464 4276
rect 13955 4236 14464 4264
rect 13955 4233 13967 4236
rect 13909 4227 13967 4233
rect 14458 4224 14464 4236
rect 14516 4224 14522 4276
rect 10888 4168 11192 4196
rect 9953 4131 10011 4137
rect 9953 4097 9965 4131
rect 9999 4097 10011 4131
rect 9953 4091 10011 4097
rect 5721 4063 5779 4069
rect 5721 4060 5733 4063
rect 4632 4032 5733 4060
rect 4249 4023 4307 4029
rect 5721 4029 5733 4032
rect 5767 4029 5779 4063
rect 6914 4060 6920 4072
rect 5721 4023 5779 4029
rect 5828 4032 6920 4060
rect 3896 3992 3924 4023
rect 4264 3992 4292 4023
rect 5828 3992 5856 4032
rect 6914 4020 6920 4032
rect 6972 4020 6978 4072
rect 7282 4060 7288 4072
rect 7243 4032 7288 4060
rect 7282 4020 7288 4032
rect 7340 4020 7346 4072
rect 7837 4063 7895 4069
rect 7837 4029 7849 4063
rect 7883 4060 7895 4063
rect 7926 4060 7932 4072
rect 7883 4032 7932 4060
rect 7883 4029 7895 4032
rect 7837 4023 7895 4029
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 9309 4063 9367 4069
rect 9309 4029 9321 4063
rect 9355 4060 9367 4063
rect 9766 4060 9772 4072
rect 9355 4032 9772 4060
rect 9355 4029 9367 4032
rect 9309 4023 9367 4029
rect 9766 4020 9772 4032
rect 9824 4020 9830 4072
rect 3896 3964 5856 3992
rect 6641 3995 6699 4001
rect 6641 3961 6653 3995
rect 6687 3992 6699 3995
rect 7190 3992 7196 4004
rect 6687 3964 7196 3992
rect 6687 3961 6699 3964
rect 6641 3955 6699 3961
rect 7190 3952 7196 3964
rect 7248 3952 7254 4004
rect 9858 3992 9864 4004
rect 9819 3964 9864 3992
rect 9858 3952 9864 3964
rect 9916 3952 9922 4004
rect 1394 3924 1400 3936
rect 1355 3896 1400 3924
rect 1394 3884 1400 3896
rect 1452 3884 1458 3936
rect 2222 3884 2228 3936
rect 2280 3924 2286 3936
rect 2682 3924 2688 3936
rect 2280 3896 2688 3924
rect 2280 3884 2286 3896
rect 2682 3884 2688 3896
rect 2740 3884 2746 3936
rect 3418 3884 3424 3936
rect 3476 3924 3482 3936
rect 3476 3896 3521 3924
rect 3476 3884 3482 3896
rect 3694 3884 3700 3936
rect 3752 3924 3758 3936
rect 6086 3924 6092 3936
rect 3752 3896 6092 3924
rect 3752 3884 3758 3896
rect 6086 3884 6092 3896
rect 6144 3884 6150 3936
rect 6178 3884 6184 3936
rect 6236 3924 6242 3936
rect 6825 3927 6883 3933
rect 6825 3924 6837 3927
rect 6236 3896 6837 3924
rect 6236 3884 6242 3896
rect 6825 3893 6837 3896
rect 6871 3893 6883 3927
rect 7374 3924 7380 3936
rect 7335 3896 7380 3924
rect 6825 3887 6883 3893
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 8202 3884 8208 3936
rect 8260 3924 8266 3936
rect 8573 3927 8631 3933
rect 8573 3924 8585 3927
rect 8260 3896 8585 3924
rect 8260 3884 8266 3896
rect 8573 3893 8585 3896
rect 8619 3893 8631 3927
rect 9030 3924 9036 3936
rect 8991 3896 9036 3924
rect 8573 3887 8631 3893
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 9766 3884 9772 3936
rect 9824 3924 9830 3936
rect 9968 3924 9996 4091
rect 10778 4060 10784 4072
rect 10739 4032 10784 4060
rect 10778 4020 10784 4032
rect 10836 4020 10842 4072
rect 10137 3995 10195 4001
rect 10137 3961 10149 3995
rect 10183 3992 10195 3995
rect 10502 3992 10508 4004
rect 10183 3964 10508 3992
rect 10183 3961 10195 3964
rect 10137 3955 10195 3961
rect 10502 3952 10508 3964
rect 10560 3952 10566 4004
rect 10888 3992 10916 4168
rect 11238 4156 11244 4208
rect 11296 4156 11302 4208
rect 11790 4196 11796 4208
rect 11532 4168 11796 4196
rect 11146 4088 11152 4140
rect 11204 4088 11210 4140
rect 11256 4128 11284 4156
rect 11532 4140 11560 4168
rect 11790 4156 11796 4168
rect 11848 4196 11854 4208
rect 12529 4199 12587 4205
rect 12529 4196 12541 4199
rect 11848 4168 12541 4196
rect 11848 4156 11854 4168
rect 12529 4165 12541 4168
rect 12575 4165 12587 4199
rect 12529 4159 12587 4165
rect 11333 4131 11391 4137
rect 11333 4128 11345 4131
rect 11256 4100 11345 4128
rect 11333 4097 11345 4100
rect 11379 4097 11391 4131
rect 11333 4091 11391 4097
rect 11514 4088 11520 4140
rect 11572 4088 11578 4140
rect 11977 4131 12035 4137
rect 11977 4097 11989 4131
rect 12023 4128 12035 4131
rect 12158 4128 12164 4140
rect 12023 4100 12164 4128
rect 12023 4097 12035 4100
rect 11977 4091 12035 4097
rect 12158 4088 12164 4100
rect 12216 4128 12222 4140
rect 13262 4128 13268 4140
rect 12216 4100 13268 4128
rect 12216 4088 12222 4100
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 14461 4131 14519 4137
rect 14461 4097 14473 4131
rect 14507 4128 14519 4131
rect 14826 4128 14832 4140
rect 14507 4100 14832 4128
rect 14507 4097 14519 4100
rect 14461 4091 14519 4097
rect 14826 4088 14832 4100
rect 14884 4088 14890 4140
rect 15654 4128 15660 4140
rect 15615 4100 15660 4128
rect 15654 4088 15660 4100
rect 15712 4088 15718 4140
rect 10965 4063 11023 4069
rect 10965 4029 10977 4063
rect 11011 4060 11023 4063
rect 11164 4060 11192 4088
rect 11011 4032 11192 4060
rect 11011 4029 11023 4032
rect 10965 4023 11023 4029
rect 11698 4020 11704 4072
rect 11756 4060 11762 4072
rect 12066 4060 12072 4072
rect 11756 4032 12072 4060
rect 11756 4020 11762 4032
rect 12066 4020 12072 4032
rect 12124 4060 12130 4072
rect 12342 4060 12348 4072
rect 12124 4032 12217 4060
rect 12303 4032 12348 4060
rect 12124 4020 12130 4032
rect 12342 4020 12348 4032
rect 12400 4020 12406 4072
rect 13170 4060 13176 4072
rect 13131 4032 13176 4060
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 13354 4060 13360 4072
rect 13315 4032 13360 4060
rect 13354 4020 13360 4032
rect 13412 4020 13418 4072
rect 14001 4063 14059 4069
rect 14001 4029 14013 4063
rect 14047 4029 14059 4063
rect 14001 4023 14059 4029
rect 14185 4063 14243 4069
rect 14185 4029 14197 4063
rect 14231 4060 14243 4063
rect 14642 4060 14648 4072
rect 14231 4032 14648 4060
rect 14231 4029 14243 4032
rect 14185 4023 14243 4029
rect 11054 3992 11060 4004
rect 10888 3964 11060 3992
rect 11054 3952 11060 3964
rect 11112 3952 11118 4004
rect 14016 3992 14044 4023
rect 12406 3964 14044 3992
rect 9824 3896 9996 3924
rect 9824 3884 9830 3896
rect 12066 3884 12072 3936
rect 12124 3924 12130 3936
rect 12406 3924 12434 3964
rect 12124 3896 12434 3924
rect 12713 3927 12771 3933
rect 12124 3884 12130 3896
rect 12713 3893 12725 3927
rect 12759 3924 12771 3927
rect 12802 3924 12808 3936
rect 12759 3896 12808 3924
rect 12759 3893 12771 3896
rect 12713 3887 12771 3893
rect 12802 3884 12808 3896
rect 12860 3884 12866 3936
rect 12894 3884 12900 3936
rect 12952 3924 12958 3936
rect 13541 3927 13599 3933
rect 13541 3924 13553 3927
rect 12952 3896 13553 3924
rect 12952 3884 12958 3896
rect 13541 3893 13553 3896
rect 13587 3893 13599 3927
rect 13541 3887 13599 3893
rect 13814 3884 13820 3936
rect 13872 3924 13878 3936
rect 14200 3924 14228 4023
rect 14642 4020 14648 4032
rect 14700 4020 14706 4072
rect 15381 4063 15439 4069
rect 15381 4029 15393 4063
rect 15427 4060 15439 4063
rect 15746 4060 15752 4072
rect 15427 4032 15752 4060
rect 15427 4029 15439 4032
rect 15381 4023 15439 4029
rect 15746 4020 15752 4032
rect 15804 4020 15810 4072
rect 14642 3924 14648 3936
rect 13872 3896 14228 3924
rect 14603 3896 14648 3924
rect 13872 3884 13878 3896
rect 14642 3884 14648 3896
rect 14700 3884 14706 3936
rect 1104 3834 16008 3856
rect 1104 3782 2824 3834
rect 2876 3782 2888 3834
rect 2940 3782 2952 3834
rect 3004 3782 3016 3834
rect 3068 3782 3080 3834
rect 3132 3782 6572 3834
rect 6624 3782 6636 3834
rect 6688 3782 6700 3834
rect 6752 3782 6764 3834
rect 6816 3782 6828 3834
rect 6880 3782 10320 3834
rect 10372 3782 10384 3834
rect 10436 3782 10448 3834
rect 10500 3782 10512 3834
rect 10564 3782 10576 3834
rect 10628 3782 14068 3834
rect 14120 3782 14132 3834
rect 14184 3782 14196 3834
rect 14248 3782 14260 3834
rect 14312 3782 14324 3834
rect 14376 3782 16008 3834
rect 1104 3760 16008 3782
rect 2314 3680 2320 3732
rect 2372 3720 2378 3732
rect 2685 3723 2743 3729
rect 2685 3720 2697 3723
rect 2372 3692 2697 3720
rect 2372 3680 2378 3692
rect 2685 3689 2697 3692
rect 2731 3689 2743 3723
rect 2685 3683 2743 3689
rect 2774 3680 2780 3732
rect 2832 3720 2838 3732
rect 3605 3723 3663 3729
rect 3605 3720 3617 3723
rect 2832 3692 3617 3720
rect 2832 3680 2838 3692
rect 3605 3689 3617 3692
rect 3651 3720 3663 3723
rect 5166 3720 5172 3732
rect 3651 3692 5172 3720
rect 3651 3689 3663 3692
rect 3605 3683 3663 3689
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 5592 3692 5672 3720
rect 5592 3680 5598 3692
rect 1854 3652 1860 3664
rect 1815 3624 1860 3652
rect 1854 3612 1860 3624
rect 1912 3612 1918 3664
rect 3694 3652 3700 3664
rect 3068 3624 3700 3652
rect 3068 3584 3096 3624
rect 3694 3612 3700 3624
rect 3752 3612 3758 3664
rect 5077 3655 5135 3661
rect 5077 3621 5089 3655
rect 5123 3621 5135 3655
rect 5077 3615 5135 3621
rect 3234 3584 3240 3596
rect 2148 3556 3096 3584
rect 3195 3556 3240 3584
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 2148 3525 2176 3556
rect 3234 3544 3240 3556
rect 3292 3544 3298 3596
rect 4522 3544 4528 3596
rect 4580 3584 4586 3596
rect 4985 3587 5043 3593
rect 4985 3584 4997 3587
rect 4580 3556 4997 3584
rect 4580 3544 4586 3556
rect 4985 3553 4997 3556
rect 5031 3553 5043 3587
rect 4985 3547 5043 3553
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3485 2191 3519
rect 2133 3479 2191 3485
rect 2409 3519 2467 3525
rect 2409 3485 2421 3519
rect 2455 3485 2467 3519
rect 2409 3479 2467 3485
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3516 3111 3519
rect 3418 3516 3424 3528
rect 3099 3488 3424 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 1486 3408 1492 3460
rect 1544 3448 1550 3460
rect 2424 3448 2452 3479
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 4062 3516 4068 3528
rect 4023 3488 4068 3516
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 4246 3476 4252 3528
rect 4304 3516 4310 3528
rect 4709 3519 4767 3525
rect 4709 3516 4721 3519
rect 4304 3488 4721 3516
rect 4304 3476 4310 3488
rect 4709 3485 4721 3488
rect 4755 3485 4767 3519
rect 4709 3479 4767 3485
rect 1544 3420 2452 3448
rect 2593 3451 2651 3457
rect 1544 3408 1550 3420
rect 2593 3417 2605 3451
rect 2639 3448 2651 3451
rect 4430 3448 4436 3460
rect 2639 3420 4436 3448
rect 2639 3417 2651 3420
rect 2593 3411 2651 3417
rect 4430 3408 4436 3420
rect 4488 3408 4494 3460
rect 5000 3448 5028 3547
rect 5092 3528 5120 3615
rect 5644 3593 5672 3692
rect 5810 3680 5816 3732
rect 5868 3720 5874 3732
rect 5997 3723 6055 3729
rect 5997 3720 6009 3723
rect 5868 3692 6009 3720
rect 5868 3680 5874 3692
rect 5997 3689 6009 3692
rect 6043 3689 6055 3723
rect 5997 3683 6055 3689
rect 6454 3680 6460 3732
rect 6512 3720 6518 3732
rect 7837 3723 7895 3729
rect 7837 3720 7849 3723
rect 6512 3692 7849 3720
rect 6512 3680 6518 3692
rect 7837 3689 7849 3692
rect 7883 3689 7895 3723
rect 7837 3683 7895 3689
rect 9490 3680 9496 3732
rect 9548 3720 9554 3732
rect 9769 3723 9827 3729
rect 9769 3720 9781 3723
rect 9548 3692 9781 3720
rect 9548 3680 9554 3692
rect 9769 3689 9781 3692
rect 9815 3689 9827 3723
rect 9769 3683 9827 3689
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 10505 3723 10563 3729
rect 10505 3720 10517 3723
rect 10008 3692 10517 3720
rect 10008 3680 10014 3692
rect 10505 3689 10517 3692
rect 10551 3689 10563 3723
rect 10505 3683 10563 3689
rect 10778 3680 10784 3732
rect 10836 3720 10842 3732
rect 11333 3723 11391 3729
rect 11333 3720 11345 3723
rect 10836 3692 11345 3720
rect 10836 3680 10842 3692
rect 11333 3689 11345 3692
rect 11379 3689 11391 3723
rect 11333 3683 11391 3689
rect 12161 3723 12219 3729
rect 12161 3689 12173 3723
rect 12207 3720 12219 3723
rect 12526 3720 12532 3732
rect 12207 3692 12532 3720
rect 12207 3689 12219 3692
rect 12161 3683 12219 3689
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 13078 3680 13084 3732
rect 13136 3720 13142 3732
rect 13136 3692 13308 3720
rect 13136 3680 13142 3692
rect 6362 3612 6368 3664
rect 6420 3652 6426 3664
rect 6420 3624 8524 3652
rect 6420 3612 6426 3624
rect 5629 3587 5687 3593
rect 5629 3553 5641 3587
rect 5675 3553 5687 3587
rect 6638 3584 6644 3596
rect 6599 3556 6644 3584
rect 5629 3547 5687 3553
rect 6638 3544 6644 3556
rect 6696 3544 6702 3596
rect 7466 3584 7472 3596
rect 7427 3556 7472 3584
rect 7466 3544 7472 3556
rect 7524 3584 7530 3596
rect 8389 3587 8447 3593
rect 8389 3584 8401 3587
rect 7524 3556 8401 3584
rect 7524 3544 7530 3556
rect 8389 3553 8401 3556
rect 8435 3553 8447 3587
rect 8389 3547 8447 3553
rect 5074 3476 5080 3528
rect 5132 3476 5138 3528
rect 5534 3516 5540 3528
rect 5495 3488 5540 3516
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 7098 3516 7104 3528
rect 6187 3488 7104 3516
rect 6187 3448 6215 3488
rect 7098 3476 7104 3488
rect 7156 3476 7162 3528
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3516 7251 3519
rect 7282 3516 7288 3528
rect 7239 3488 7288 3516
rect 7239 3485 7251 3488
rect 7193 3479 7251 3485
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 7742 3516 7748 3528
rect 7703 3488 7748 3516
rect 7742 3476 7748 3488
rect 7800 3516 7806 3528
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 7800 3488 8217 3516
rect 7800 3476 7806 3488
rect 8205 3485 8217 3488
rect 8251 3485 8263 3519
rect 8496 3516 8524 3624
rect 9030 3612 9036 3664
rect 9088 3652 9094 3664
rect 9088 3624 13124 3652
rect 9088 3612 9094 3624
rect 8938 3544 8944 3596
rect 8996 3584 9002 3596
rect 9125 3587 9183 3593
rect 9125 3584 9137 3587
rect 8996 3556 9137 3584
rect 8996 3544 9002 3556
rect 9125 3553 9137 3556
rect 9171 3553 9183 3587
rect 9674 3584 9680 3596
rect 9125 3547 9183 3553
rect 9232 3556 9680 3584
rect 9232 3516 9260 3556
rect 9674 3544 9680 3556
rect 9732 3584 9738 3596
rect 10594 3584 10600 3596
rect 9732 3556 10600 3584
rect 9732 3544 9738 3556
rect 10594 3544 10600 3556
rect 10652 3544 10658 3596
rect 11149 3587 11207 3593
rect 10888 3556 11100 3584
rect 8496 3488 9260 3516
rect 8205 3479 8263 3485
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 9364 3488 9720 3516
rect 9364 3476 9370 3488
rect 6457 3451 6515 3457
rect 6457 3448 6469 3451
rect 5000 3420 6215 3448
rect 6288 3420 6469 3448
rect 6288 3392 6316 3420
rect 6457 3417 6469 3420
rect 6503 3417 6515 3451
rect 8754 3448 8760 3460
rect 8667 3420 8760 3448
rect 6457 3411 6515 3417
rect 8754 3408 8760 3420
rect 8812 3448 8818 3460
rect 9582 3448 9588 3460
rect 8812 3420 9588 3448
rect 8812 3408 8818 3420
rect 9582 3408 9588 3420
rect 9640 3408 9646 3460
rect 9692 3448 9720 3488
rect 10134 3476 10140 3528
rect 10192 3516 10198 3528
rect 10888 3525 10916 3556
rect 10873 3519 10931 3525
rect 10873 3516 10885 3519
rect 10192 3488 10885 3516
rect 10192 3476 10198 3488
rect 10873 3485 10885 3488
rect 10919 3485 10931 3519
rect 10873 3479 10931 3485
rect 10962 3476 10968 3528
rect 11020 3476 11026 3528
rect 11072 3516 11100 3556
rect 11149 3553 11161 3587
rect 11195 3584 11207 3587
rect 11238 3584 11244 3596
rect 11195 3556 11244 3584
rect 11195 3553 11207 3556
rect 11149 3547 11207 3553
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 11808 3593 11836 3624
rect 11793 3587 11851 3593
rect 11793 3553 11805 3587
rect 11839 3553 11851 3587
rect 11974 3584 11980 3596
rect 11935 3556 11980 3584
rect 11793 3547 11851 3553
rect 11974 3544 11980 3556
rect 12032 3544 12038 3596
rect 12618 3544 12624 3596
rect 12676 3584 12682 3596
rect 13096 3593 13124 3624
rect 12713 3587 12771 3593
rect 12713 3584 12725 3587
rect 12676 3556 12725 3584
rect 12676 3544 12682 3556
rect 12713 3553 12725 3556
rect 12759 3553 12771 3587
rect 12713 3547 12771 3553
rect 13081 3587 13139 3593
rect 13081 3553 13093 3587
rect 13127 3584 13139 3587
rect 13170 3584 13176 3596
rect 13127 3556 13176 3584
rect 13127 3553 13139 3556
rect 13081 3547 13139 3553
rect 13170 3544 13176 3556
rect 13228 3544 13234 3596
rect 13280 3584 13308 3692
rect 13354 3680 13360 3732
rect 13412 3720 13418 3732
rect 15102 3720 15108 3732
rect 13412 3692 15108 3720
rect 13412 3680 13418 3692
rect 15102 3680 15108 3692
rect 15160 3680 15166 3732
rect 13722 3612 13728 3664
rect 13780 3652 13786 3664
rect 14093 3655 14151 3661
rect 14093 3652 14105 3655
rect 13780 3624 14105 3652
rect 13780 3612 13786 3624
rect 14093 3621 14105 3624
rect 14139 3621 14151 3655
rect 14093 3615 14151 3621
rect 14737 3655 14795 3661
rect 14737 3621 14749 3655
rect 14783 3652 14795 3655
rect 14918 3652 14924 3664
rect 14783 3624 14924 3652
rect 14783 3621 14795 3624
rect 14737 3615 14795 3621
rect 14918 3612 14924 3624
rect 14976 3612 14982 3664
rect 13357 3587 13415 3593
rect 13357 3584 13369 3587
rect 13280 3556 13369 3584
rect 13357 3553 13369 3556
rect 13403 3553 13415 3587
rect 14826 3584 14832 3596
rect 14739 3556 14832 3584
rect 13357 3547 13415 3553
rect 14826 3544 14832 3556
rect 14884 3584 14890 3596
rect 15562 3584 15568 3596
rect 14884 3556 15568 3584
rect 14884 3544 14890 3556
rect 15562 3544 15568 3556
rect 15620 3544 15626 3596
rect 12529 3519 12587 3525
rect 11072 3488 11284 3516
rect 10321 3451 10379 3457
rect 9692 3420 10272 3448
rect 1578 3380 1584 3392
rect 1539 3352 1584 3380
rect 1578 3340 1584 3352
rect 1636 3340 1642 3392
rect 1854 3340 1860 3392
rect 1912 3380 1918 3392
rect 1949 3383 2007 3389
rect 1949 3380 1961 3383
rect 1912 3352 1961 3380
rect 1912 3340 1918 3352
rect 1949 3349 1961 3352
rect 1995 3349 2007 3383
rect 2222 3380 2228 3392
rect 2183 3352 2228 3380
rect 1949 3343 2007 3349
rect 2222 3340 2228 3352
rect 2280 3340 2286 3392
rect 3142 3380 3148 3392
rect 3103 3352 3148 3380
rect 3142 3340 3148 3352
rect 3200 3340 3206 3392
rect 3878 3380 3884 3392
rect 3839 3352 3884 3380
rect 3878 3340 3884 3352
rect 3936 3340 3942 3392
rect 5166 3340 5172 3392
rect 5224 3380 5230 3392
rect 5445 3383 5503 3389
rect 5445 3380 5457 3383
rect 5224 3352 5457 3380
rect 5224 3340 5230 3352
rect 5445 3349 5457 3352
rect 5491 3380 5503 3383
rect 5534 3380 5540 3392
rect 5491 3352 5540 3380
rect 5491 3349 5503 3352
rect 5445 3343 5503 3349
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 6270 3340 6276 3392
rect 6328 3340 6334 3392
rect 6365 3383 6423 3389
rect 6365 3349 6377 3383
rect 6411 3380 6423 3383
rect 6825 3383 6883 3389
rect 6825 3380 6837 3383
rect 6411 3352 6837 3380
rect 6411 3349 6423 3352
rect 6365 3343 6423 3349
rect 6825 3349 6837 3352
rect 6871 3349 6883 3383
rect 6825 3343 6883 3349
rect 7006 3340 7012 3392
rect 7064 3380 7070 3392
rect 7285 3383 7343 3389
rect 7285 3380 7297 3383
rect 7064 3352 7297 3380
rect 7064 3340 7070 3352
rect 7285 3349 7297 3352
rect 7331 3380 7343 3383
rect 7558 3380 7564 3392
rect 7331 3352 7564 3380
rect 7331 3349 7343 3352
rect 7285 3343 7343 3349
rect 7558 3340 7564 3352
rect 7616 3340 7622 3392
rect 7926 3340 7932 3392
rect 7984 3380 7990 3392
rect 8297 3383 8355 3389
rect 8297 3380 8309 3383
rect 7984 3352 8309 3380
rect 7984 3340 7990 3352
rect 8297 3349 8309 3352
rect 8343 3380 8355 3383
rect 8938 3380 8944 3392
rect 8343 3352 8944 3380
rect 8343 3349 8355 3352
rect 8297 3343 8355 3349
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 9306 3380 9312 3392
rect 9267 3352 9312 3380
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 9398 3340 9404 3392
rect 9456 3380 9462 3392
rect 10042 3380 10048 3392
rect 9456 3352 9501 3380
rect 10003 3352 10048 3380
rect 9456 3340 9462 3352
rect 10042 3340 10048 3352
rect 10100 3340 10106 3392
rect 10244 3389 10272 3420
rect 10321 3417 10333 3451
rect 10367 3448 10379 3451
rect 10980 3448 11008 3476
rect 11256 3460 11284 3488
rect 12529 3485 12541 3519
rect 12575 3516 12587 3519
rect 12894 3516 12900 3528
rect 12575 3488 12900 3516
rect 12575 3485 12587 3488
rect 12529 3479 12587 3485
rect 12894 3476 12900 3488
rect 12952 3476 12958 3528
rect 13722 3476 13728 3528
rect 13780 3516 13786 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 13780 3488 14289 3516
rect 13780 3476 13786 3488
rect 14277 3485 14289 3488
rect 14323 3516 14335 3519
rect 14734 3516 14740 3528
rect 14323 3488 14740 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 14734 3476 14740 3488
rect 14792 3476 14798 3528
rect 15010 3476 15016 3528
rect 15068 3516 15074 3528
rect 15105 3519 15163 3525
rect 15105 3516 15117 3519
rect 15068 3488 15117 3516
rect 15068 3476 15074 3488
rect 15105 3485 15117 3488
rect 15151 3485 15163 3519
rect 15105 3479 15163 3485
rect 11146 3448 11152 3460
rect 10367 3420 11152 3448
rect 10367 3417 10379 3420
rect 10321 3411 10379 3417
rect 11146 3408 11152 3420
rect 11204 3408 11210 3460
rect 11238 3408 11244 3460
rect 11296 3408 11302 3460
rect 11701 3451 11759 3457
rect 11701 3417 11713 3451
rect 11747 3448 11759 3451
rect 12434 3448 12440 3460
rect 11747 3420 12440 3448
rect 11747 3417 11759 3420
rect 11701 3411 11759 3417
rect 12434 3408 12440 3420
rect 12492 3408 12498 3460
rect 13906 3408 13912 3460
rect 13964 3448 13970 3460
rect 14553 3451 14611 3457
rect 14553 3448 14565 3451
rect 13964 3420 14565 3448
rect 13964 3408 13970 3420
rect 14553 3417 14565 3420
rect 14599 3417 14611 3451
rect 14553 3411 14611 3417
rect 10229 3383 10287 3389
rect 10229 3349 10241 3383
rect 10275 3349 10287 3383
rect 10229 3343 10287 3349
rect 10962 3340 10968 3392
rect 11020 3380 11026 3392
rect 11020 3352 11065 3380
rect 11020 3340 11026 3352
rect 12618 3340 12624 3392
rect 12676 3380 12682 3392
rect 12676 3352 12721 3380
rect 12676 3340 12682 3352
rect 13170 3340 13176 3392
rect 13228 3380 13234 3392
rect 13630 3380 13636 3392
rect 13228 3352 13636 3380
rect 13228 3340 13234 3352
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 14458 3340 14464 3392
rect 14516 3380 14522 3392
rect 15010 3380 15016 3392
rect 14516 3352 15016 3380
rect 14516 3340 14522 3352
rect 15010 3340 15016 3352
rect 15068 3340 15074 3392
rect 1104 3290 16008 3312
rect 1104 3238 4698 3290
rect 4750 3238 4762 3290
rect 4814 3238 4826 3290
rect 4878 3238 4890 3290
rect 4942 3238 4954 3290
rect 5006 3238 8446 3290
rect 8498 3238 8510 3290
rect 8562 3238 8574 3290
rect 8626 3238 8638 3290
rect 8690 3238 8702 3290
rect 8754 3238 12194 3290
rect 12246 3238 12258 3290
rect 12310 3238 12322 3290
rect 12374 3238 12386 3290
rect 12438 3238 12450 3290
rect 12502 3238 16008 3290
rect 1104 3216 16008 3238
rect 1964 3148 3096 3176
rect 1964 3049 1992 3148
rect 2682 3068 2688 3120
rect 2740 3108 2746 3120
rect 3068 3108 3096 3148
rect 3142 3136 3148 3188
rect 3200 3176 3206 3188
rect 3697 3179 3755 3185
rect 3697 3176 3709 3179
rect 3200 3148 3709 3176
rect 3200 3136 3206 3148
rect 3697 3145 3709 3148
rect 3743 3145 3755 3179
rect 3697 3139 3755 3145
rect 4157 3179 4215 3185
rect 4157 3145 4169 3179
rect 4203 3176 4215 3179
rect 4522 3176 4528 3188
rect 4203 3148 4528 3176
rect 4203 3145 4215 3148
rect 4157 3139 4215 3145
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 5077 3179 5135 3185
rect 5077 3145 5089 3179
rect 5123 3145 5135 3179
rect 5077 3139 5135 3145
rect 3970 3108 3976 3120
rect 2740 3080 2912 3108
rect 3068 3080 3976 3108
rect 2740 3068 2746 3080
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 1949 3043 2007 3049
rect 1719 3012 1808 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 1780 2913 1808 3012
rect 1949 3009 1961 3043
rect 1995 3009 2007 3043
rect 1949 3003 2007 3009
rect 2038 3000 2044 3052
rect 2096 3040 2102 3052
rect 2225 3043 2283 3049
rect 2225 3040 2237 3043
rect 2096 3012 2237 3040
rect 2096 3000 2102 3012
rect 2225 3009 2237 3012
rect 2271 3009 2283 3043
rect 2225 3003 2283 3009
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3040 2375 3043
rect 2406 3040 2412 3052
rect 2363 3012 2412 3040
rect 2363 3009 2375 3012
rect 2317 3003 2375 3009
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 2774 3040 2780 3052
rect 2735 3012 2780 3040
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 2884 3049 2912 3080
rect 3970 3068 3976 3080
rect 4028 3108 4034 3120
rect 4065 3111 4123 3117
rect 4065 3108 4077 3111
rect 4028 3080 4077 3108
rect 4028 3068 4034 3080
rect 4065 3077 4077 3080
rect 4111 3077 4123 3111
rect 5092 3108 5120 3139
rect 5166 3136 5172 3188
rect 5224 3176 5230 3188
rect 5442 3176 5448 3188
rect 5224 3148 5448 3176
rect 5224 3136 5230 3148
rect 5442 3136 5448 3148
rect 5500 3136 5506 3188
rect 5629 3179 5687 3185
rect 5629 3145 5641 3179
rect 5675 3176 5687 3179
rect 6086 3176 6092 3188
rect 5675 3148 6092 3176
rect 5675 3145 5687 3148
rect 5629 3139 5687 3145
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 6270 3136 6276 3188
rect 6328 3176 6334 3188
rect 6365 3179 6423 3185
rect 6365 3176 6377 3179
rect 6328 3148 6377 3176
rect 6328 3136 6334 3148
rect 6365 3145 6377 3148
rect 6411 3145 6423 3179
rect 6365 3139 6423 3145
rect 6733 3179 6791 3185
rect 6733 3145 6745 3179
rect 6779 3176 6791 3179
rect 6822 3176 6828 3188
rect 6779 3148 6828 3176
rect 6779 3145 6791 3148
rect 6733 3139 6791 3145
rect 5092 3080 5764 3108
rect 4065 3071 4123 3077
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3009 2927 3043
rect 2869 3003 2927 3009
rect 3421 3043 3479 3049
rect 3421 3009 3433 3043
rect 3467 3040 3479 3043
rect 3878 3040 3884 3052
rect 3467 3012 3884 3040
rect 3467 3009 3479 3012
rect 3421 3003 3479 3009
rect 3878 3000 3884 3012
rect 3936 3000 3942 3052
rect 4614 3000 4620 3052
rect 4672 3040 4678 3052
rect 4801 3043 4859 3049
rect 4801 3040 4813 3043
rect 4672 3012 4813 3040
rect 4672 3000 4678 3012
rect 4801 3009 4813 3012
rect 4847 3009 4859 3043
rect 4801 3003 4859 3009
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3040 4951 3043
rect 5258 3040 5264 3052
rect 4939 3012 5264 3040
rect 4939 3009 4951 3012
rect 4893 3003 4951 3009
rect 5258 3000 5264 3012
rect 5316 3000 5322 3052
rect 5353 3043 5411 3049
rect 5353 3009 5365 3043
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 5445 3043 5503 3049
rect 5445 3009 5457 3043
rect 5491 3040 5503 3043
rect 5626 3040 5632 3052
rect 5491 3012 5632 3040
rect 5491 3009 5503 3012
rect 5445 3003 5503 3009
rect 4338 2972 4344 2984
rect 4299 2944 4344 2972
rect 4338 2932 4344 2944
rect 4396 2972 4402 2984
rect 5166 2972 5172 2984
rect 4396 2944 5172 2972
rect 4396 2932 4402 2944
rect 5166 2932 5172 2944
rect 5224 2932 5230 2984
rect 5368 2972 5396 3003
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 5736 3049 5764 3080
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3009 5779 3043
rect 5721 3003 5779 3009
rect 5902 2972 5908 2984
rect 5368 2944 5908 2972
rect 5902 2932 5908 2944
rect 5960 2932 5966 2984
rect 1765 2907 1823 2913
rect 1765 2873 1777 2907
rect 1811 2873 1823 2907
rect 1765 2867 1823 2873
rect 2501 2907 2559 2913
rect 2501 2873 2513 2907
rect 2547 2904 2559 2907
rect 2682 2904 2688 2916
rect 2547 2876 2688 2904
rect 2547 2873 2559 2876
rect 2501 2867 2559 2873
rect 2682 2864 2688 2876
rect 2740 2864 2746 2916
rect 3053 2907 3111 2913
rect 3053 2873 3065 2907
rect 3099 2904 3111 2907
rect 3142 2904 3148 2916
rect 3099 2876 3148 2904
rect 3099 2873 3111 2876
rect 3053 2867 3111 2873
rect 3142 2864 3148 2876
rect 3200 2864 3206 2916
rect 3605 2907 3663 2913
rect 3605 2873 3617 2907
rect 3651 2904 3663 2907
rect 6748 2904 6776 3139
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7098 3136 7104 3188
rect 7156 3176 7162 3188
rect 7650 3176 7656 3188
rect 7156 3148 7656 3176
rect 7156 3136 7162 3148
rect 7650 3136 7656 3148
rect 7708 3176 7714 3188
rect 8021 3179 8079 3185
rect 8021 3176 8033 3179
rect 7708 3148 8033 3176
rect 7708 3136 7714 3148
rect 8021 3145 8033 3148
rect 8067 3145 8079 3179
rect 8938 3176 8944 3188
rect 8899 3148 8944 3176
rect 8021 3139 8079 3145
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 9306 3136 9312 3188
rect 9364 3176 9370 3188
rect 9401 3179 9459 3185
rect 9401 3176 9413 3179
rect 9364 3148 9413 3176
rect 9364 3136 9370 3148
rect 9401 3145 9413 3148
rect 9447 3145 9459 3179
rect 9401 3139 9459 3145
rect 9769 3179 9827 3185
rect 9769 3145 9781 3179
rect 9815 3176 9827 3179
rect 9815 3148 9996 3176
rect 9815 3145 9827 3148
rect 9769 3139 9827 3145
rect 7834 3068 7840 3120
rect 7892 3108 7898 3120
rect 9968 3108 9996 3148
rect 10042 3136 10048 3188
rect 10100 3176 10106 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 10100 3148 10609 3176
rect 10100 3136 10106 3148
rect 10597 3145 10609 3148
rect 10643 3145 10655 3179
rect 10597 3139 10655 3145
rect 10689 3179 10747 3185
rect 10689 3145 10701 3179
rect 10735 3145 10747 3179
rect 10689 3139 10747 3145
rect 11149 3179 11207 3185
rect 11149 3145 11161 3179
rect 11195 3176 11207 3179
rect 11330 3176 11336 3188
rect 11195 3148 11336 3176
rect 11195 3145 11207 3148
rect 11149 3139 11207 3145
rect 10226 3108 10232 3120
rect 7892 3080 9168 3108
rect 9968 3080 10232 3108
rect 7892 3068 7898 3080
rect 7190 3040 7196 3052
rect 7151 3012 7196 3040
rect 7190 3000 7196 3012
rect 7248 3000 7254 3052
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3040 7711 3043
rect 7742 3040 7748 3052
rect 7699 3012 7748 3040
rect 7699 3009 7711 3012
rect 7653 3003 7711 3009
rect 7742 3000 7748 3012
rect 7800 3000 7806 3052
rect 8110 3040 8116 3052
rect 8071 3012 8116 3040
rect 8110 3000 8116 3012
rect 8168 3000 8174 3052
rect 8202 3000 8208 3052
rect 8260 3040 8266 3052
rect 9033 3043 9091 3049
rect 9033 3040 9045 3043
rect 8260 3012 9045 3040
rect 8260 3000 8266 3012
rect 9033 3009 9045 3012
rect 9079 3009 9091 3043
rect 9033 3003 9091 3009
rect 6825 2975 6883 2981
rect 6825 2941 6837 2975
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 7009 2975 7067 2981
rect 7009 2941 7021 2975
rect 7055 2972 7067 2975
rect 7466 2972 7472 2984
rect 7055 2944 7472 2972
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 3651 2876 6776 2904
rect 6840 2904 6868 2935
rect 7466 2932 7472 2944
rect 7524 2932 7530 2984
rect 7834 2972 7840 2984
rect 7795 2944 7840 2972
rect 7834 2932 7840 2944
rect 7892 2932 7898 2984
rect 9140 2981 9168 3080
rect 10226 3068 10232 3080
rect 10284 3068 10290 3120
rect 9306 3000 9312 3052
rect 9364 3040 9370 3052
rect 9582 3040 9588 3052
rect 9364 3012 9588 3040
rect 9364 3000 9370 3012
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 9858 3040 9864 3052
rect 9819 3012 9864 3040
rect 9858 3000 9864 3012
rect 9916 3000 9922 3052
rect 9125 2975 9183 2981
rect 9125 2941 9137 2975
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 9674 2932 9680 2984
rect 9732 2972 9738 2984
rect 9950 2972 9956 2984
rect 9732 2944 9956 2972
rect 9732 2932 9738 2944
rect 9950 2932 9956 2944
rect 10008 2972 10014 2984
rect 10008 2944 10548 2972
rect 10008 2932 10014 2944
rect 6914 2904 6920 2916
rect 6840 2876 6920 2904
rect 3651 2873 3663 2876
rect 3605 2867 3663 2873
rect 6914 2864 6920 2876
rect 6972 2904 6978 2916
rect 7190 2904 7196 2916
rect 6972 2876 7196 2904
rect 6972 2864 6978 2876
rect 7190 2864 7196 2876
rect 7248 2864 7254 2916
rect 8386 2864 8392 2916
rect 8444 2904 8450 2916
rect 8573 2907 8631 2913
rect 8573 2904 8585 2907
rect 8444 2876 8585 2904
rect 8444 2864 8450 2876
rect 8573 2873 8585 2876
rect 8619 2873 8631 2907
rect 8573 2867 8631 2873
rect 9398 2864 9404 2916
rect 9456 2904 9462 2916
rect 10229 2907 10287 2913
rect 10229 2904 10241 2907
rect 9456 2876 10241 2904
rect 9456 2864 9462 2876
rect 10229 2873 10241 2876
rect 10275 2873 10287 2907
rect 10229 2867 10287 2873
rect 1210 2796 1216 2848
rect 1268 2836 1274 2848
rect 1489 2839 1547 2845
rect 1489 2836 1501 2839
rect 1268 2808 1501 2836
rect 1268 2796 1274 2808
rect 1489 2805 1501 2808
rect 1535 2805 1547 2839
rect 2038 2836 2044 2848
rect 1999 2808 2044 2836
rect 1489 2799 1547 2805
rect 2038 2796 2044 2808
rect 2096 2796 2102 2848
rect 2590 2796 2596 2848
rect 2648 2836 2654 2848
rect 3234 2836 3240 2848
rect 2648 2808 2693 2836
rect 3195 2808 3240 2836
rect 2648 2796 2654 2808
rect 3234 2796 3240 2808
rect 3292 2796 3298 2848
rect 4617 2839 4675 2845
rect 4617 2805 4629 2839
rect 4663 2836 4675 2839
rect 4706 2836 4712 2848
rect 4663 2808 4712 2836
rect 4663 2805 4675 2808
rect 4617 2799 4675 2805
rect 4706 2796 4712 2808
rect 4764 2796 4770 2848
rect 5166 2796 5172 2848
rect 5224 2836 5230 2848
rect 5224 2808 5269 2836
rect 5224 2796 5230 2808
rect 5718 2796 5724 2848
rect 5776 2836 5782 2848
rect 5905 2839 5963 2845
rect 5905 2836 5917 2839
rect 5776 2808 5917 2836
rect 5776 2796 5782 2808
rect 5905 2805 5917 2808
rect 5951 2805 5963 2839
rect 5905 2799 5963 2805
rect 6181 2839 6239 2845
rect 6181 2805 6193 2839
rect 6227 2836 6239 2839
rect 7006 2836 7012 2848
rect 6227 2808 7012 2836
rect 6227 2805 6239 2808
rect 6181 2799 6239 2805
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 7098 2796 7104 2848
rect 7156 2836 7162 2848
rect 7377 2839 7435 2845
rect 7377 2836 7389 2839
rect 7156 2808 7389 2836
rect 7156 2796 7162 2808
rect 7377 2805 7389 2808
rect 7423 2805 7435 2839
rect 8478 2836 8484 2848
rect 8439 2808 8484 2836
rect 7377 2799 7435 2805
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 10520 2836 10548 2944
rect 10594 2864 10600 2916
rect 10652 2904 10658 2916
rect 10704 2904 10732 3139
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 12066 3136 12072 3188
rect 12124 3176 12130 3188
rect 12253 3179 12311 3185
rect 12253 3176 12265 3179
rect 12124 3148 12265 3176
rect 12124 3136 12130 3148
rect 12253 3145 12265 3148
rect 12299 3145 12311 3179
rect 12253 3139 12311 3145
rect 12345 3179 12403 3185
rect 12345 3145 12357 3179
rect 12391 3176 12403 3179
rect 12618 3176 12624 3188
rect 12391 3148 12624 3176
rect 12391 3145 12403 3148
rect 12345 3139 12403 3145
rect 12618 3136 12624 3148
rect 12676 3136 12682 3188
rect 12802 3176 12808 3188
rect 12763 3148 12808 3176
rect 12802 3136 12808 3148
rect 12860 3136 12866 3188
rect 10870 3068 10876 3120
rect 10928 3108 10934 3120
rect 11241 3111 11299 3117
rect 11241 3108 11253 3111
rect 10928 3080 11253 3108
rect 10928 3068 10934 3080
rect 11241 3077 11253 3080
rect 11287 3077 11299 3111
rect 11241 3071 11299 3077
rect 11422 3068 11428 3120
rect 11480 3108 11486 3120
rect 11793 3111 11851 3117
rect 11793 3108 11805 3111
rect 11480 3080 11805 3108
rect 11480 3068 11486 3080
rect 11793 3077 11805 3080
rect 11839 3077 11851 3111
rect 12710 3108 12716 3120
rect 12671 3080 12716 3108
rect 11793 3071 11851 3077
rect 12710 3068 12716 3080
rect 12768 3068 12774 3120
rect 11885 3043 11943 3049
rect 11885 3009 11897 3043
rect 11931 3009 11943 3043
rect 13814 3040 13820 3052
rect 11885 3003 11943 3009
rect 13096 3012 13820 3040
rect 10781 2975 10839 2981
rect 10781 2941 10793 2975
rect 10827 2941 10839 2975
rect 10781 2935 10839 2941
rect 11701 2975 11759 2981
rect 11701 2941 11713 2975
rect 11747 2941 11759 2975
rect 11900 2972 11928 3003
rect 11974 2972 11980 2984
rect 11900 2944 11980 2972
rect 11701 2935 11759 2941
rect 10652 2876 10732 2904
rect 10652 2864 10658 2876
rect 10796 2836 10824 2935
rect 11716 2904 11744 2935
rect 11974 2932 11980 2944
rect 12032 2932 12038 2984
rect 12989 2975 13047 2981
rect 12989 2941 13001 2975
rect 13035 2972 13047 2975
rect 13096 2972 13124 3012
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 14090 3040 14096 3052
rect 14051 3012 14096 3040
rect 14090 3000 14096 3012
rect 14148 3000 14154 3052
rect 14277 3043 14335 3049
rect 14277 3009 14289 3043
rect 14323 3009 14335 3043
rect 14550 3040 14556 3052
rect 14511 3012 14556 3040
rect 14277 3003 14335 3009
rect 13035 2944 13124 2972
rect 13173 2975 13231 2981
rect 13035 2941 13047 2944
rect 12989 2935 13047 2941
rect 13173 2941 13185 2975
rect 13219 2972 13231 2975
rect 13262 2972 13268 2984
rect 13219 2944 13268 2972
rect 13219 2941 13231 2944
rect 13173 2935 13231 2941
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 13449 2975 13507 2981
rect 13449 2941 13461 2975
rect 13495 2972 13507 2975
rect 13495 2944 13584 2972
rect 13495 2941 13507 2944
rect 13449 2935 13507 2941
rect 13556 2904 13584 2944
rect 13630 2932 13636 2984
rect 13688 2972 13694 2984
rect 14292 2972 14320 3003
rect 14550 3000 14556 3012
rect 14608 3000 14614 3052
rect 15657 3043 15715 3049
rect 15657 3009 15669 3043
rect 15703 3040 15715 3043
rect 15838 3040 15844 3052
rect 15703 3012 15844 3040
rect 15703 3009 15715 3012
rect 15657 3003 15715 3009
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 13688 2944 14320 2972
rect 13688 2932 13694 2944
rect 14366 2932 14372 2984
rect 14424 2972 14430 2984
rect 14829 2975 14887 2981
rect 14829 2972 14841 2975
rect 14424 2944 14841 2972
rect 14424 2932 14430 2944
rect 14829 2941 14841 2944
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 13814 2904 13820 2916
rect 11716 2876 13492 2904
rect 13556 2876 13820 2904
rect 13464 2848 13492 2876
rect 13814 2864 13820 2876
rect 13872 2864 13878 2916
rect 10520 2808 10824 2836
rect 11606 2796 11612 2848
rect 11664 2836 11670 2848
rect 11790 2836 11796 2848
rect 11664 2808 11796 2836
rect 11664 2796 11670 2808
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 12066 2796 12072 2848
rect 12124 2836 12130 2848
rect 13170 2836 13176 2848
rect 12124 2808 13176 2836
rect 12124 2796 12130 2808
rect 13170 2796 13176 2808
rect 13228 2796 13234 2848
rect 13446 2796 13452 2848
rect 13504 2796 13510 2848
rect 15378 2796 15384 2848
rect 15436 2836 15442 2848
rect 15473 2839 15531 2845
rect 15473 2836 15485 2839
rect 15436 2808 15485 2836
rect 15436 2796 15442 2808
rect 15473 2805 15485 2808
rect 15519 2805 15531 2839
rect 15473 2799 15531 2805
rect 1104 2746 16008 2768
rect 1104 2694 2824 2746
rect 2876 2694 2888 2746
rect 2940 2694 2952 2746
rect 3004 2694 3016 2746
rect 3068 2694 3080 2746
rect 3132 2694 6572 2746
rect 6624 2694 6636 2746
rect 6688 2694 6700 2746
rect 6752 2694 6764 2746
rect 6816 2694 6828 2746
rect 6880 2694 10320 2746
rect 10372 2694 10384 2746
rect 10436 2694 10448 2746
rect 10500 2694 10512 2746
rect 10564 2694 10576 2746
rect 10628 2694 14068 2746
rect 14120 2694 14132 2746
rect 14184 2694 14196 2746
rect 14248 2694 14260 2746
rect 14312 2694 14324 2746
rect 14376 2694 16008 2746
rect 1104 2672 16008 2694
rect 7745 2635 7803 2641
rect 7745 2601 7757 2635
rect 7791 2632 7803 2635
rect 8202 2632 8208 2644
rect 7791 2604 8208 2632
rect 7791 2601 7803 2604
rect 7745 2595 7803 2601
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 9030 2632 9036 2644
rect 8991 2604 9036 2632
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 9401 2635 9459 2641
rect 9401 2601 9413 2635
rect 9447 2632 9459 2635
rect 9766 2632 9772 2644
rect 9447 2604 9772 2632
rect 9447 2601 9459 2604
rect 9401 2595 9459 2601
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 10413 2635 10471 2641
rect 10413 2601 10425 2635
rect 10459 2632 10471 2635
rect 10962 2632 10968 2644
rect 10459 2604 10968 2632
rect 10459 2601 10471 2604
rect 10413 2595 10471 2601
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 12207 2635 12265 2641
rect 12207 2601 12219 2635
rect 12253 2632 12265 2635
rect 15010 2632 15016 2644
rect 12253 2604 15016 2632
rect 12253 2601 12265 2604
rect 12207 2595 12265 2601
rect 15010 2592 15016 2604
rect 15068 2592 15074 2644
rect 3973 2567 4031 2573
rect 3973 2533 3985 2567
rect 4019 2533 4031 2567
rect 3973 2527 4031 2533
rect 7469 2567 7527 2573
rect 7469 2533 7481 2567
rect 7515 2564 7527 2567
rect 7834 2564 7840 2576
rect 7515 2536 7840 2564
rect 7515 2533 7527 2536
rect 7469 2527 7527 2533
rect 2038 2496 2044 2508
rect 1780 2468 2044 2496
rect 1780 2437 1808 2468
rect 2038 2456 2044 2468
rect 2096 2456 2102 2508
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 1854 2388 1860 2440
rect 1912 2428 1918 2440
rect 2222 2428 2228 2440
rect 1912 2400 1957 2428
rect 2183 2400 2228 2428
rect 1912 2388 1918 2400
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 2590 2428 2596 2440
rect 2551 2400 2596 2428
rect 2590 2388 2596 2400
rect 2648 2388 2654 2440
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 2961 2431 3019 2437
rect 2961 2428 2973 2431
rect 2832 2400 2973 2428
rect 2832 2388 2838 2400
rect 2961 2397 2973 2400
rect 3007 2397 3019 2431
rect 2961 2391 3019 2397
rect 3142 2388 3148 2440
rect 3200 2428 3206 2440
rect 3329 2431 3387 2437
rect 3329 2428 3341 2431
rect 3200 2400 3341 2428
rect 3200 2388 3206 2400
rect 3329 2397 3341 2400
rect 3375 2397 3387 2431
rect 3786 2428 3792 2440
rect 3747 2400 3792 2428
rect 3329 2391 3387 2397
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 3988 2428 4016 2527
rect 7834 2524 7840 2536
rect 7892 2524 7898 2576
rect 8018 2564 8024 2576
rect 7979 2536 8024 2564
rect 8018 2524 8024 2536
rect 8076 2524 8082 2576
rect 9490 2524 9496 2576
rect 9548 2564 9554 2576
rect 11517 2567 11575 2573
rect 11517 2564 11529 2567
rect 9548 2536 11529 2564
rect 9548 2524 9554 2536
rect 11517 2533 11529 2536
rect 11563 2533 11575 2567
rect 11517 2527 11575 2533
rect 5994 2496 6000 2508
rect 5092 2468 6000 2496
rect 4065 2431 4123 2437
rect 4065 2428 4077 2431
rect 3988 2400 4077 2428
rect 4065 2397 4077 2400
rect 4111 2397 4123 2431
rect 4706 2428 4712 2440
rect 4667 2400 4712 2428
rect 4065 2391 4123 2397
rect 4706 2388 4712 2400
rect 4764 2388 4770 2440
rect 5092 2437 5120 2468
rect 5994 2456 6000 2468
rect 6052 2456 6058 2508
rect 6086 2456 6092 2508
rect 6144 2496 6150 2508
rect 8294 2496 8300 2508
rect 6144 2468 6592 2496
rect 6144 2456 6150 2468
rect 5077 2431 5135 2437
rect 5077 2397 5089 2431
rect 5123 2397 5135 2431
rect 5077 2391 5135 2397
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 5810 2428 5816 2440
rect 5224 2400 5269 2428
rect 5771 2400 5816 2428
rect 5224 2388 5230 2400
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 6178 2428 6184 2440
rect 6139 2400 6184 2428
rect 6178 2388 6184 2400
rect 6236 2388 6242 2440
rect 6564 2437 6592 2468
rect 7208 2468 8300 2496
rect 7208 2437 7236 2468
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 8478 2496 8484 2508
rect 8439 2468 8484 2496
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 8665 2499 8723 2505
rect 8665 2465 8677 2499
rect 8711 2496 8723 2499
rect 9582 2496 9588 2508
rect 8711 2468 9588 2496
rect 8711 2465 8723 2468
rect 8665 2459 8723 2465
rect 9582 2456 9588 2468
rect 9640 2456 9646 2508
rect 9858 2496 9864 2508
rect 9819 2468 9864 2496
rect 9858 2456 9864 2468
rect 9916 2456 9922 2508
rect 9953 2499 10011 2505
rect 9953 2465 9965 2499
rect 9999 2496 10011 2499
rect 10318 2496 10324 2508
rect 9999 2468 10324 2496
rect 9999 2465 10011 2468
rect 9953 2459 10011 2465
rect 10318 2456 10324 2468
rect 10376 2456 10382 2508
rect 15194 2496 15200 2508
rect 10428 2468 15200 2496
rect 6549 2431 6607 2437
rect 6549 2397 6561 2431
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 7193 2431 7251 2437
rect 7193 2397 7205 2431
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2428 7343 2431
rect 7374 2428 7380 2440
rect 7331 2400 7380 2428
rect 7331 2397 7343 2400
rect 7285 2391 7343 2397
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 7926 2428 7932 2440
rect 7887 2400 7932 2428
rect 7926 2388 7932 2400
rect 7984 2388 7990 2440
rect 8386 2428 8392 2440
rect 8347 2400 8392 2428
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 10428 2428 10456 2468
rect 9048 2400 10456 2428
rect 10505 2431 10563 2437
rect 3602 2320 3608 2372
rect 3660 2360 3666 2372
rect 9048 2360 9076 2400
rect 10505 2397 10517 2431
rect 10551 2428 10563 2431
rect 10686 2428 10692 2440
rect 10551 2400 10692 2428
rect 10551 2397 10563 2400
rect 10505 2391 10563 2397
rect 3660 2332 9076 2360
rect 9125 2363 9183 2369
rect 3660 2320 3666 2332
rect 9125 2329 9137 2363
rect 9171 2329 9183 2363
rect 9125 2323 9183 2329
rect 9493 2363 9551 2369
rect 9493 2329 9505 2363
rect 9539 2360 9551 2363
rect 9674 2360 9680 2372
rect 9539 2332 9680 2360
rect 9539 2329 9551 2332
rect 9493 2323 9551 2329
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 1946 2252 1952 2304
rect 2004 2292 2010 2304
rect 2041 2295 2099 2301
rect 2041 2292 2053 2295
rect 2004 2264 2053 2292
rect 2004 2252 2010 2264
rect 2041 2261 2053 2264
rect 2087 2261 2099 2295
rect 2041 2255 2099 2261
rect 2314 2252 2320 2304
rect 2372 2292 2378 2304
rect 2409 2295 2467 2301
rect 2409 2292 2421 2295
rect 2372 2264 2421 2292
rect 2372 2252 2378 2264
rect 2409 2261 2421 2264
rect 2455 2261 2467 2295
rect 2409 2255 2467 2261
rect 2682 2252 2688 2304
rect 2740 2292 2746 2304
rect 2777 2295 2835 2301
rect 2777 2292 2789 2295
rect 2740 2264 2789 2292
rect 2740 2252 2746 2264
rect 2777 2261 2789 2264
rect 2823 2261 2835 2295
rect 2777 2255 2835 2261
rect 3145 2295 3203 2301
rect 3145 2261 3157 2295
rect 3191 2292 3203 2295
rect 3418 2292 3424 2304
rect 3191 2264 3424 2292
rect 3191 2261 3203 2264
rect 3145 2255 3203 2261
rect 3418 2252 3424 2264
rect 3476 2252 3482 2304
rect 3513 2295 3571 2301
rect 3513 2261 3525 2295
rect 3559 2292 3571 2295
rect 3786 2292 3792 2304
rect 3559 2264 3792 2292
rect 3559 2261 3571 2264
rect 3513 2255 3571 2261
rect 3786 2252 3792 2264
rect 3844 2252 3850 2304
rect 4154 2252 4160 2304
rect 4212 2292 4218 2304
rect 4249 2295 4307 2301
rect 4249 2292 4261 2295
rect 4212 2264 4261 2292
rect 4212 2252 4218 2264
rect 4249 2261 4261 2264
rect 4295 2261 4307 2295
rect 4522 2292 4528 2304
rect 4483 2264 4528 2292
rect 4249 2255 4307 2261
rect 4522 2252 4528 2264
rect 4580 2252 4586 2304
rect 4893 2295 4951 2301
rect 4893 2261 4905 2295
rect 4939 2292 4951 2295
rect 5074 2292 5080 2304
rect 4939 2264 5080 2292
rect 4939 2261 4951 2264
rect 4893 2255 4951 2261
rect 5074 2252 5080 2264
rect 5132 2252 5138 2304
rect 5258 2252 5264 2304
rect 5316 2292 5322 2304
rect 5353 2295 5411 2301
rect 5353 2292 5365 2295
rect 5316 2264 5365 2292
rect 5316 2252 5322 2264
rect 5353 2261 5365 2264
rect 5399 2261 5411 2295
rect 5353 2255 5411 2261
rect 5629 2295 5687 2301
rect 5629 2261 5641 2295
rect 5675 2292 5687 2295
rect 5902 2292 5908 2304
rect 5675 2264 5908 2292
rect 5675 2261 5687 2264
rect 5629 2255 5687 2261
rect 5902 2252 5908 2264
rect 5960 2252 5966 2304
rect 5997 2295 6055 2301
rect 5997 2261 6009 2295
rect 6043 2292 6055 2295
rect 6270 2292 6276 2304
rect 6043 2264 6276 2292
rect 6043 2261 6055 2264
rect 5997 2255 6055 2261
rect 6270 2252 6276 2264
rect 6328 2252 6334 2304
rect 6454 2292 6460 2304
rect 6415 2264 6460 2292
rect 6454 2252 6460 2264
rect 6512 2252 6518 2304
rect 6730 2292 6736 2304
rect 6691 2264 6736 2292
rect 6730 2252 6736 2264
rect 6788 2252 6794 2304
rect 7009 2295 7067 2301
rect 7009 2261 7021 2295
rect 7055 2292 7067 2295
rect 7466 2292 7472 2304
rect 7055 2264 7472 2292
rect 7055 2261 7067 2264
rect 7009 2255 7067 2261
rect 7466 2252 7472 2264
rect 7524 2252 7530 2304
rect 8938 2252 8944 2304
rect 8996 2292 9002 2304
rect 9140 2292 9168 2323
rect 9674 2320 9680 2332
rect 9732 2320 9738 2372
rect 9784 2332 10364 2360
rect 9784 2292 9812 2332
rect 8996 2264 9812 2292
rect 10045 2295 10103 2301
rect 8996 2252 9002 2264
rect 10045 2261 10057 2295
rect 10091 2292 10103 2295
rect 10226 2292 10232 2304
rect 10091 2264 10232 2292
rect 10091 2261 10103 2264
rect 10045 2255 10103 2261
rect 10226 2252 10232 2264
rect 10284 2252 10290 2304
rect 10336 2292 10364 2332
rect 10410 2320 10416 2372
rect 10468 2360 10474 2372
rect 10520 2360 10548 2391
rect 10686 2388 10692 2400
rect 10744 2388 10750 2440
rect 10781 2431 10839 2437
rect 10781 2397 10793 2431
rect 10827 2428 10839 2431
rect 11422 2428 11428 2440
rect 10827 2400 11428 2428
rect 10827 2397 10839 2400
rect 10781 2391 10839 2397
rect 10468 2332 10548 2360
rect 10468 2320 10474 2332
rect 10594 2320 10600 2372
rect 10652 2360 10658 2372
rect 10796 2360 10824 2391
rect 11422 2388 11428 2400
rect 11480 2388 11486 2440
rect 11698 2428 11704 2440
rect 11659 2400 11704 2428
rect 11698 2388 11704 2400
rect 11756 2388 11762 2440
rect 11974 2428 11980 2440
rect 11935 2400 11980 2428
rect 11974 2388 11980 2400
rect 12032 2388 12038 2440
rect 12618 2388 12624 2440
rect 12676 2428 12682 2440
rect 12894 2428 12900 2440
rect 12676 2400 12900 2428
rect 12676 2388 12682 2400
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 13173 2431 13231 2437
rect 13173 2428 13185 2431
rect 13004 2400 13185 2428
rect 10652 2332 10824 2360
rect 10652 2320 10658 2332
rect 11238 2320 11244 2372
rect 11296 2360 11302 2372
rect 13004 2360 13032 2400
rect 13173 2397 13185 2400
rect 13219 2397 13231 2431
rect 13173 2391 13231 2397
rect 13538 2388 13544 2440
rect 13596 2428 13602 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 13596 2400 14105 2428
rect 13596 2388 13602 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14366 2428 14372 2440
rect 14327 2400 14372 2428
rect 14093 2391 14151 2397
rect 14366 2388 14372 2400
rect 14424 2388 14430 2440
rect 15120 2437 15148 2468
rect 15194 2456 15200 2468
rect 15252 2456 15258 2508
rect 15381 2499 15439 2505
rect 15381 2465 15393 2499
rect 15427 2496 15439 2499
rect 15470 2496 15476 2508
rect 15427 2468 15476 2496
rect 15427 2465 15439 2468
rect 15381 2459 15439 2465
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 15105 2431 15163 2437
rect 15105 2397 15117 2431
rect 15151 2397 15163 2431
rect 15105 2391 15163 2397
rect 11296 2332 13032 2360
rect 11296 2320 11302 2332
rect 13078 2320 13084 2372
rect 13136 2360 13142 2372
rect 13556 2360 13584 2388
rect 13136 2332 13584 2360
rect 13136 2320 13142 2332
rect 13817 2295 13875 2301
rect 13817 2292 13829 2295
rect 10336 2264 13829 2292
rect 13817 2261 13829 2264
rect 13863 2261 13875 2295
rect 13817 2255 13875 2261
rect 1104 2202 16008 2224
rect 1104 2150 4698 2202
rect 4750 2150 4762 2202
rect 4814 2150 4826 2202
rect 4878 2150 4890 2202
rect 4942 2150 4954 2202
rect 5006 2150 8446 2202
rect 8498 2150 8510 2202
rect 8562 2150 8574 2202
rect 8626 2150 8638 2202
rect 8690 2150 8702 2202
rect 8754 2150 12194 2202
rect 12246 2150 12258 2202
rect 12310 2150 12322 2202
rect 12374 2150 12386 2202
rect 12438 2150 12450 2202
rect 12502 2150 16008 2202
rect 1104 2128 16008 2150
rect 6454 2048 6460 2100
rect 6512 2088 6518 2100
rect 6512 2060 7880 2088
rect 6512 2048 6518 2060
rect 5810 1980 5816 2032
rect 5868 2020 5874 2032
rect 7852 2020 7880 2060
rect 7926 2048 7932 2100
rect 7984 2088 7990 2100
rect 15378 2088 15384 2100
rect 7984 2060 15384 2088
rect 7984 2048 7990 2060
rect 15378 2048 15384 2060
rect 15436 2048 15442 2100
rect 9674 2020 9680 2032
rect 5868 1992 6914 2020
rect 7852 1992 9680 2020
rect 5868 1980 5874 1992
rect 6886 1952 6914 1992
rect 9674 1980 9680 1992
rect 9732 1980 9738 2032
rect 9858 1980 9864 2032
rect 9916 2020 9922 2032
rect 11606 2020 11612 2032
rect 9916 1992 11612 2020
rect 9916 1980 9922 1992
rect 11606 1980 11612 1992
rect 11664 1980 11670 2032
rect 11054 1952 11060 1964
rect 6886 1924 11060 1952
rect 11054 1912 11060 1924
rect 11112 1912 11118 1964
rect 10042 1504 10048 1556
rect 10100 1544 10106 1556
rect 11698 1544 11704 1556
rect 10100 1516 11704 1544
rect 10100 1504 10106 1516
rect 11698 1504 11704 1516
rect 11756 1504 11762 1556
<< via1 >>
rect 4068 17756 4120 17808
rect 15292 17756 15344 17808
rect 5356 17688 5408 17740
rect 13544 17688 13596 17740
rect 7472 17620 7524 17672
rect 10140 17620 10192 17672
rect 7012 17552 7064 17604
rect 8208 17552 8260 17604
rect 13452 17552 13504 17604
rect 7380 17484 7432 17536
rect 8024 17484 8076 17536
rect 4698 17382 4750 17434
rect 4762 17382 4814 17434
rect 4826 17382 4878 17434
rect 4890 17382 4942 17434
rect 4954 17382 5006 17434
rect 8446 17382 8498 17434
rect 8510 17382 8562 17434
rect 8574 17382 8626 17434
rect 8638 17382 8690 17434
rect 8702 17382 8754 17434
rect 12194 17382 12246 17434
rect 12258 17382 12310 17434
rect 12322 17382 12374 17434
rect 12386 17382 12438 17434
rect 12450 17382 12502 17434
rect 1768 17280 1820 17332
rect 2136 17280 2188 17332
rect 2504 17280 2556 17332
rect 2872 17280 2924 17332
rect 3240 17280 3292 17332
rect 3608 17280 3660 17332
rect 4068 17280 4120 17332
rect 4344 17280 4396 17332
rect 4620 17280 4672 17332
rect 5448 17280 5500 17332
rect 1768 17187 1820 17196
rect 1768 17153 1777 17187
rect 1777 17153 1811 17187
rect 1811 17153 1820 17187
rect 1768 17144 1820 17153
rect 2412 17144 2464 17196
rect 4436 17212 4488 17264
rect 6920 17280 6972 17332
rect 7380 17280 7432 17332
rect 7564 17323 7616 17332
rect 7564 17289 7573 17323
rect 7573 17289 7607 17323
rect 7607 17289 7616 17323
rect 7564 17280 7616 17289
rect 8024 17323 8076 17332
rect 8024 17289 8033 17323
rect 8033 17289 8067 17323
rect 8067 17289 8076 17323
rect 8024 17280 8076 17289
rect 8300 17280 8352 17332
rect 13452 17323 13504 17332
rect 13452 17289 13461 17323
rect 13461 17289 13495 17323
rect 13495 17289 13504 17323
rect 13452 17280 13504 17289
rect 6552 17212 6604 17264
rect 3240 17187 3292 17196
rect 3240 17153 3249 17187
rect 3249 17153 3283 17187
rect 3283 17153 3292 17187
rect 3240 17144 3292 17153
rect 3332 17187 3384 17196
rect 3332 17153 3341 17187
rect 3341 17153 3375 17187
rect 3375 17153 3384 17187
rect 3332 17144 3384 17153
rect 3148 17076 3200 17128
rect 1032 17008 1084 17060
rect 4252 17144 4304 17196
rect 4712 17187 4764 17196
rect 4712 17153 4721 17187
rect 4721 17153 4755 17187
rect 4755 17153 4764 17187
rect 4712 17144 4764 17153
rect 5356 17144 5408 17196
rect 5448 17187 5500 17196
rect 5448 17153 5457 17187
rect 5457 17153 5491 17187
rect 5491 17153 5500 17187
rect 5816 17187 5868 17196
rect 5448 17144 5500 17153
rect 5816 17153 5825 17187
rect 5825 17153 5859 17187
rect 5859 17153 5868 17187
rect 5816 17144 5868 17153
rect 5172 17076 5224 17128
rect 6460 17144 6512 17196
rect 7932 17187 7984 17196
rect 6184 17008 6236 17060
rect 7288 17076 7340 17128
rect 7932 17153 7941 17187
rect 7941 17153 7975 17187
rect 7975 17153 7984 17187
rect 7932 17144 7984 17153
rect 8208 17119 8260 17128
rect 7656 17008 7708 17060
rect 8208 17085 8217 17119
rect 8217 17085 8251 17119
rect 8251 17085 8260 17119
rect 8208 17076 8260 17085
rect 8300 17008 8352 17060
rect 9680 17144 9732 17196
rect 9956 17144 10008 17196
rect 10140 17144 10192 17196
rect 10692 17144 10744 17196
rect 10876 17144 10928 17196
rect 11704 17144 11756 17196
rect 12532 17144 12584 17196
rect 13084 17144 13136 17196
rect 9404 17076 9456 17128
rect 10048 17076 10100 17128
rect 10232 17076 10284 17128
rect 11796 17119 11848 17128
rect 11796 17085 11805 17119
rect 11805 17085 11839 17119
rect 11839 17085 11848 17119
rect 11796 17076 11848 17085
rect 12716 17119 12768 17128
rect 12716 17085 12725 17119
rect 12725 17085 12759 17119
rect 12759 17085 12768 17119
rect 12716 17076 12768 17085
rect 13176 17076 13228 17128
rect 11060 17008 11112 17060
rect 14464 17144 14516 17196
rect 15384 17144 15436 17196
rect 14372 17119 14424 17128
rect 14372 17085 14381 17119
rect 14381 17085 14415 17119
rect 14415 17085 14424 17119
rect 14372 17076 14424 17085
rect 15200 17076 15252 17128
rect 15108 17008 15160 17060
rect 5448 16940 5500 16992
rect 8024 16940 8076 16992
rect 9036 16983 9088 16992
rect 9036 16949 9045 16983
rect 9045 16949 9079 16983
rect 9079 16949 9088 16983
rect 9036 16940 9088 16949
rect 9588 16940 9640 16992
rect 10140 16940 10192 16992
rect 10692 16940 10744 16992
rect 13820 16940 13872 16992
rect 15844 16940 15896 16992
rect 16028 16940 16080 16992
rect 2824 16838 2876 16890
rect 2888 16838 2940 16890
rect 2952 16838 3004 16890
rect 3016 16838 3068 16890
rect 3080 16838 3132 16890
rect 6572 16838 6624 16890
rect 6636 16838 6688 16890
rect 6700 16838 6752 16890
rect 6764 16838 6816 16890
rect 6828 16838 6880 16890
rect 10320 16838 10372 16890
rect 10384 16838 10436 16890
rect 10448 16838 10500 16890
rect 10512 16838 10564 16890
rect 10576 16838 10628 16890
rect 14068 16838 14120 16890
rect 14132 16838 14184 16890
rect 14196 16838 14248 16890
rect 14260 16838 14312 16890
rect 14324 16838 14376 16890
rect 1768 16736 1820 16788
rect 3148 16736 3200 16788
rect 3332 16779 3384 16788
rect 3332 16745 3341 16779
rect 3341 16745 3375 16779
rect 3375 16745 3384 16779
rect 3332 16736 3384 16745
rect 5172 16736 5224 16788
rect 6276 16736 6328 16788
rect 7932 16736 7984 16788
rect 8024 16736 8076 16788
rect 11612 16736 11664 16788
rect 13636 16736 13688 16788
rect 1952 16711 2004 16720
rect 1952 16677 1961 16711
rect 1961 16677 1995 16711
rect 1995 16677 2004 16711
rect 1952 16668 2004 16677
rect 2320 16668 2372 16720
rect 3240 16668 3292 16720
rect 7748 16711 7800 16720
rect 2504 16600 2556 16652
rect 7748 16677 7757 16711
rect 7757 16677 7791 16711
rect 7791 16677 7800 16711
rect 7748 16668 7800 16677
rect 8944 16711 8996 16720
rect 8944 16677 8953 16711
rect 8953 16677 8987 16711
rect 8987 16677 8996 16711
rect 8944 16668 8996 16677
rect 9312 16668 9364 16720
rect 9588 16668 9640 16720
rect 2136 16575 2188 16584
rect 2136 16541 2145 16575
rect 2145 16541 2179 16575
rect 2179 16541 2188 16575
rect 2136 16532 2188 16541
rect 2228 16575 2280 16584
rect 2228 16541 2237 16575
rect 2237 16541 2271 16575
rect 2271 16541 2280 16575
rect 2228 16532 2280 16541
rect 2688 16464 2740 16516
rect 1400 16396 1452 16448
rect 3240 16532 3292 16584
rect 3608 16575 3660 16584
rect 3608 16541 3617 16575
rect 3617 16541 3651 16575
rect 3651 16541 3660 16575
rect 3608 16532 3660 16541
rect 3884 16532 3936 16584
rect 4068 16575 4120 16584
rect 4068 16541 4077 16575
rect 4077 16541 4111 16575
rect 4111 16541 4120 16575
rect 4068 16532 4120 16541
rect 4528 16532 4580 16584
rect 4160 16464 4212 16516
rect 7196 16600 7248 16652
rect 7288 16643 7340 16652
rect 7288 16609 7297 16643
rect 7297 16609 7331 16643
rect 7331 16609 7340 16643
rect 7288 16600 7340 16609
rect 8208 16600 8260 16652
rect 10140 16643 10192 16652
rect 7104 16575 7156 16584
rect 3700 16396 3752 16448
rect 3976 16396 4028 16448
rect 5632 16464 5684 16516
rect 5172 16396 5224 16448
rect 5724 16439 5776 16448
rect 5724 16405 5733 16439
rect 5733 16405 5767 16439
rect 5767 16405 5776 16439
rect 5724 16396 5776 16405
rect 6368 16439 6420 16448
rect 6368 16405 6377 16439
rect 6377 16405 6411 16439
rect 6411 16405 6420 16439
rect 6368 16396 6420 16405
rect 7104 16541 7113 16575
rect 7113 16541 7147 16575
rect 7147 16541 7156 16575
rect 7104 16532 7156 16541
rect 7380 16532 7432 16584
rect 7656 16464 7708 16516
rect 8852 16532 8904 16584
rect 7932 16464 7984 16516
rect 8116 16439 8168 16448
rect 8116 16405 8125 16439
rect 8125 16405 8159 16439
rect 8159 16405 8168 16439
rect 8116 16396 8168 16405
rect 8392 16396 8444 16448
rect 8852 16396 8904 16448
rect 10140 16609 10149 16643
rect 10149 16609 10183 16643
rect 10183 16609 10192 16643
rect 10140 16600 10192 16609
rect 10784 16668 10836 16720
rect 10324 16600 10376 16652
rect 12716 16643 12768 16652
rect 9128 16575 9180 16584
rect 9128 16541 9137 16575
rect 9137 16541 9171 16575
rect 9171 16541 9180 16575
rect 9128 16532 9180 16541
rect 9220 16532 9272 16584
rect 9312 16464 9364 16516
rect 9680 16532 9732 16584
rect 10600 16532 10652 16584
rect 10968 16532 11020 16584
rect 12716 16609 12725 16643
rect 12725 16609 12759 16643
rect 12759 16609 12768 16643
rect 12716 16600 12768 16609
rect 11520 16532 11572 16584
rect 12072 16532 12124 16584
rect 13268 16600 13320 16652
rect 13452 16600 13504 16652
rect 13820 16600 13872 16652
rect 14648 16643 14700 16652
rect 14648 16609 14657 16643
rect 14657 16609 14691 16643
rect 14691 16609 14700 16643
rect 14648 16600 14700 16609
rect 16304 16736 16356 16788
rect 15292 16600 15344 16652
rect 11244 16464 11296 16516
rect 15568 16464 15620 16516
rect 9496 16396 9548 16448
rect 9680 16439 9732 16448
rect 9680 16405 9689 16439
rect 9689 16405 9723 16439
rect 9723 16405 9732 16439
rect 9680 16396 9732 16405
rect 10048 16439 10100 16448
rect 10048 16405 10057 16439
rect 10057 16405 10091 16439
rect 10091 16405 10100 16439
rect 10048 16396 10100 16405
rect 10968 16396 11020 16448
rect 15476 16439 15528 16448
rect 15476 16405 15485 16439
rect 15485 16405 15519 16439
rect 15519 16405 15528 16439
rect 15476 16396 15528 16405
rect 4698 16294 4750 16346
rect 4762 16294 4814 16346
rect 4826 16294 4878 16346
rect 4890 16294 4942 16346
rect 4954 16294 5006 16346
rect 8446 16294 8498 16346
rect 8510 16294 8562 16346
rect 8574 16294 8626 16346
rect 8638 16294 8690 16346
rect 8702 16294 8754 16346
rect 12194 16294 12246 16346
rect 12258 16294 12310 16346
rect 12322 16294 12374 16346
rect 12386 16294 12438 16346
rect 12450 16294 12502 16346
rect 2136 16235 2188 16244
rect 2136 16201 2145 16235
rect 2145 16201 2179 16235
rect 2179 16201 2188 16235
rect 2136 16192 2188 16201
rect 4068 16192 4120 16244
rect 4252 16235 4304 16244
rect 4252 16201 4261 16235
rect 4261 16201 4295 16235
rect 4295 16201 4304 16235
rect 4252 16192 4304 16201
rect 6000 16192 6052 16244
rect 6828 16235 6880 16244
rect 6828 16201 6837 16235
rect 6837 16201 6871 16235
rect 6871 16201 6880 16235
rect 6828 16192 6880 16201
rect 7748 16235 7800 16244
rect 7748 16201 7757 16235
rect 7757 16201 7791 16235
rect 7791 16201 7800 16235
rect 7748 16192 7800 16201
rect 8116 16192 8168 16244
rect 10048 16192 10100 16244
rect 11612 16192 11664 16244
rect 12072 16192 12124 16244
rect 13544 16235 13596 16244
rect 13544 16201 13553 16235
rect 13553 16201 13587 16235
rect 13587 16201 13596 16235
rect 13544 16192 13596 16201
rect 14464 16192 14516 16244
rect 16396 16192 16448 16244
rect 3976 16124 4028 16176
rect 6920 16124 6972 16176
rect 2320 16099 2372 16108
rect 2320 16065 2329 16099
rect 2329 16065 2363 16099
rect 2363 16065 2372 16099
rect 2320 16056 2372 16065
rect 2596 16099 2648 16108
rect 2596 16065 2605 16099
rect 2605 16065 2639 16099
rect 2639 16065 2648 16099
rect 2596 16056 2648 16065
rect 2688 16056 2740 16108
rect 3516 16099 3568 16108
rect 3516 16065 3525 16099
rect 3525 16065 3559 16099
rect 3559 16065 3568 16099
rect 3516 16056 3568 16065
rect 4344 16056 4396 16108
rect 5264 16056 5316 16108
rect 5724 16099 5776 16108
rect 5724 16065 5733 16099
rect 5733 16065 5767 16099
rect 5767 16065 5776 16099
rect 5724 16056 5776 16065
rect 6092 16056 6144 16108
rect 7012 16056 7064 16108
rect 7932 16124 7984 16176
rect 9128 16124 9180 16176
rect 9864 16124 9916 16176
rect 8116 16056 8168 16108
rect 8944 16056 8996 16108
rect 9496 16056 9548 16108
rect 10508 16124 10560 16176
rect 10600 16124 10652 16176
rect 12808 16124 12860 16176
rect 13452 16124 13504 16176
rect 15660 16167 15712 16176
rect 15660 16133 15669 16167
rect 15669 16133 15703 16167
rect 15703 16133 15712 16167
rect 15660 16124 15712 16133
rect 3424 15988 3476 16040
rect 4068 15988 4120 16040
rect 5172 16031 5224 16040
rect 2780 15920 2832 15972
rect 4160 15920 4212 15972
rect 5172 15997 5181 16031
rect 5181 15997 5215 16031
rect 5215 15997 5224 16031
rect 5172 15988 5224 15997
rect 5908 15988 5960 16040
rect 7656 16031 7708 16040
rect 7656 15997 7665 16031
rect 7665 15997 7699 16031
rect 7699 15997 7708 16031
rect 7656 15988 7708 15997
rect 8484 16031 8536 16040
rect 8484 15997 8493 16031
rect 8493 15997 8527 16031
rect 8527 15997 8536 16031
rect 8484 15988 8536 15997
rect 8852 15988 8904 16040
rect 9588 15988 9640 16040
rect 9956 15988 10008 16040
rect 11336 16056 11388 16108
rect 12992 16056 13044 16108
rect 10416 16031 10468 16040
rect 10416 15997 10425 16031
rect 10425 15997 10459 16031
rect 10459 15997 10468 16031
rect 10416 15988 10468 15997
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 4344 15852 4396 15904
rect 4528 15895 4580 15904
rect 4528 15861 4537 15895
rect 4537 15861 4571 15895
rect 4571 15861 4580 15895
rect 4528 15852 4580 15861
rect 5540 15852 5592 15904
rect 7564 15852 7616 15904
rect 8392 15852 8444 15904
rect 8484 15852 8536 15904
rect 9496 15852 9548 15904
rect 9956 15852 10008 15904
rect 10508 15920 10560 15972
rect 12624 15988 12676 16040
rect 13820 16031 13872 16040
rect 12532 15920 12584 15972
rect 13820 15997 13829 16031
rect 13829 15997 13863 16031
rect 13863 15997 13872 16031
rect 13820 15988 13872 15997
rect 15476 15988 15528 16040
rect 13176 15963 13228 15972
rect 13176 15929 13185 15963
rect 13185 15929 13219 15963
rect 13219 15929 13228 15963
rect 13176 15920 13228 15929
rect 10692 15852 10744 15904
rect 11244 15895 11296 15904
rect 11244 15861 11253 15895
rect 11253 15861 11287 15895
rect 11287 15861 11296 15895
rect 11244 15852 11296 15861
rect 12348 15895 12400 15904
rect 12348 15861 12357 15895
rect 12357 15861 12391 15895
rect 12391 15861 12400 15895
rect 12348 15852 12400 15861
rect 2824 15750 2876 15802
rect 2888 15750 2940 15802
rect 2952 15750 3004 15802
rect 3016 15750 3068 15802
rect 3080 15750 3132 15802
rect 6572 15750 6624 15802
rect 6636 15750 6688 15802
rect 6700 15750 6752 15802
rect 6764 15750 6816 15802
rect 6828 15750 6880 15802
rect 10320 15750 10372 15802
rect 10384 15750 10436 15802
rect 10448 15750 10500 15802
rect 10512 15750 10564 15802
rect 10576 15750 10628 15802
rect 14068 15750 14120 15802
rect 14132 15750 14184 15802
rect 14196 15750 14248 15802
rect 14260 15750 14312 15802
rect 14324 15750 14376 15802
rect 1400 15691 1452 15700
rect 1400 15657 1409 15691
rect 1409 15657 1443 15691
rect 1443 15657 1452 15691
rect 1400 15648 1452 15657
rect 2228 15648 2280 15700
rect 2412 15648 2464 15700
rect 3424 15691 3476 15700
rect 3424 15657 3433 15691
rect 3433 15657 3467 15691
rect 3467 15657 3476 15691
rect 3424 15648 3476 15657
rect 2136 15580 2188 15632
rect 2596 15580 2648 15632
rect 2780 15512 2832 15564
rect 3332 15512 3384 15564
rect 3884 15512 3936 15564
rect 4436 15648 4488 15700
rect 5448 15691 5500 15700
rect 5448 15657 5457 15691
rect 5457 15657 5491 15691
rect 5491 15657 5500 15691
rect 5448 15648 5500 15657
rect 5816 15691 5868 15700
rect 5816 15657 5825 15691
rect 5825 15657 5859 15691
rect 5859 15657 5868 15691
rect 5816 15648 5868 15657
rect 6368 15691 6420 15700
rect 6368 15657 6377 15691
rect 6377 15657 6411 15691
rect 6411 15657 6420 15691
rect 6368 15648 6420 15657
rect 5356 15580 5408 15632
rect 7472 15648 7524 15700
rect 8944 15691 8996 15700
rect 8944 15657 8953 15691
rect 8953 15657 8987 15691
rect 8987 15657 8996 15691
rect 8944 15648 8996 15657
rect 10232 15691 10284 15700
rect 10232 15657 10241 15691
rect 10241 15657 10275 15691
rect 10275 15657 10284 15691
rect 10232 15648 10284 15657
rect 11060 15648 11112 15700
rect 12624 15691 12676 15700
rect 4252 15512 4304 15564
rect 4528 15487 4580 15496
rect 4528 15453 4537 15487
rect 4537 15453 4571 15487
rect 4571 15453 4580 15487
rect 4528 15444 4580 15453
rect 5448 15512 5500 15564
rect 5724 15555 5776 15564
rect 5724 15521 5733 15555
rect 5733 15521 5767 15555
rect 5767 15521 5776 15555
rect 5724 15512 5776 15521
rect 6276 15555 6328 15564
rect 6276 15521 6285 15555
rect 6285 15521 6319 15555
rect 6319 15521 6328 15555
rect 6276 15512 6328 15521
rect 5816 15444 5868 15496
rect 5632 15376 5684 15428
rect 6092 15376 6144 15428
rect 7288 15512 7340 15564
rect 7840 15512 7892 15564
rect 8392 15580 8444 15632
rect 7104 15444 7156 15496
rect 8208 15444 8260 15496
rect 9404 15512 9456 15564
rect 9036 15444 9088 15496
rect 9864 15444 9916 15496
rect 12348 15580 12400 15632
rect 12624 15657 12633 15691
rect 12633 15657 12667 15691
rect 12667 15657 12676 15691
rect 12624 15648 12676 15657
rect 10968 15444 11020 15496
rect 11060 15444 11112 15496
rect 11796 15512 11848 15564
rect 12072 15512 12124 15564
rect 11888 15444 11940 15496
rect 12900 15512 12952 15564
rect 12716 15444 12768 15496
rect 14280 15512 14332 15564
rect 15016 15512 15068 15564
rect 15292 15512 15344 15564
rect 7380 15376 7432 15428
rect 2044 15351 2096 15360
rect 2044 15317 2053 15351
rect 2053 15317 2087 15351
rect 2087 15317 2096 15351
rect 2044 15308 2096 15317
rect 2136 15351 2188 15360
rect 2136 15317 2145 15351
rect 2145 15317 2179 15351
rect 2179 15317 2188 15351
rect 2412 15351 2464 15360
rect 2136 15308 2188 15317
rect 2412 15317 2421 15351
rect 2421 15317 2455 15351
rect 2455 15317 2464 15351
rect 2412 15308 2464 15317
rect 2780 15308 2832 15360
rect 3056 15351 3108 15360
rect 3056 15317 3065 15351
rect 3065 15317 3099 15351
rect 3099 15317 3108 15351
rect 3056 15308 3108 15317
rect 3424 15308 3476 15360
rect 3792 15351 3844 15360
rect 3792 15317 3801 15351
rect 3801 15317 3835 15351
rect 3835 15317 3844 15351
rect 3792 15308 3844 15317
rect 4620 15351 4672 15360
rect 4620 15317 4629 15351
rect 4629 15317 4663 15351
rect 4663 15317 4672 15351
rect 4620 15308 4672 15317
rect 6828 15351 6880 15360
rect 6828 15317 6837 15351
rect 6837 15317 6871 15351
rect 6871 15317 6880 15351
rect 7472 15351 7524 15360
rect 6828 15308 6880 15317
rect 7472 15317 7481 15351
rect 7481 15317 7515 15351
rect 7515 15317 7524 15351
rect 7472 15308 7524 15317
rect 8208 15308 8260 15360
rect 8392 15351 8444 15360
rect 8392 15317 8401 15351
rect 8401 15317 8435 15351
rect 8435 15317 8444 15351
rect 8392 15308 8444 15317
rect 8944 15308 8996 15360
rect 10508 15376 10560 15428
rect 10232 15308 10284 15360
rect 10784 15376 10836 15428
rect 11980 15376 12032 15428
rect 13544 15376 13596 15428
rect 14556 15444 14608 15496
rect 14004 15376 14056 15428
rect 14464 15376 14516 15428
rect 14740 15444 14792 15496
rect 14924 15376 14976 15428
rect 11152 15308 11204 15360
rect 11428 15351 11480 15360
rect 11428 15317 11437 15351
rect 11437 15317 11471 15351
rect 11471 15317 11480 15351
rect 11428 15308 11480 15317
rect 12072 15308 12124 15360
rect 12808 15351 12860 15360
rect 12808 15317 12817 15351
rect 12817 15317 12851 15351
rect 12851 15317 12860 15351
rect 12808 15308 12860 15317
rect 13636 15351 13688 15360
rect 13636 15317 13645 15351
rect 13645 15317 13679 15351
rect 13679 15317 13688 15351
rect 13636 15308 13688 15317
rect 13820 15308 13872 15360
rect 13912 15308 13964 15360
rect 14556 15351 14608 15360
rect 14556 15317 14565 15351
rect 14565 15317 14599 15351
rect 14599 15317 14608 15351
rect 14556 15308 14608 15317
rect 4698 15206 4750 15258
rect 4762 15206 4814 15258
rect 4826 15206 4878 15258
rect 4890 15206 4942 15258
rect 4954 15206 5006 15258
rect 8446 15206 8498 15258
rect 8510 15206 8562 15258
rect 8574 15206 8626 15258
rect 8638 15206 8690 15258
rect 8702 15206 8754 15258
rect 12194 15206 12246 15258
rect 12258 15206 12310 15258
rect 12322 15206 12374 15258
rect 12386 15206 12438 15258
rect 12450 15206 12502 15258
rect 3424 15104 3476 15156
rect 3792 15104 3844 15156
rect 1584 14968 1636 15020
rect 1952 15011 2004 15020
rect 1952 14977 1961 15011
rect 1961 14977 1995 15011
rect 1995 14977 2004 15011
rect 1952 14968 2004 14977
rect 3148 15036 3200 15088
rect 4620 15104 4672 15156
rect 5356 15104 5408 15156
rect 3700 14968 3752 15020
rect 4252 14968 4304 15020
rect 4436 14968 4488 15020
rect 3424 14900 3476 14952
rect 3608 14943 3660 14952
rect 3608 14909 3617 14943
rect 3617 14909 3651 14943
rect 3651 14909 3660 14943
rect 3608 14900 3660 14909
rect 3792 14943 3844 14952
rect 3792 14909 3801 14943
rect 3801 14909 3835 14943
rect 3835 14909 3844 14943
rect 3792 14900 3844 14909
rect 3976 14900 4028 14952
rect 6000 15104 6052 15156
rect 6828 15104 6880 15156
rect 7564 15104 7616 15156
rect 7748 15147 7800 15156
rect 7748 15113 7757 15147
rect 7757 15113 7791 15147
rect 7791 15113 7800 15147
rect 7748 15104 7800 15113
rect 8852 15104 8904 15156
rect 6184 15079 6236 15088
rect 5080 14968 5132 15020
rect 6184 15045 6193 15079
rect 6193 15045 6227 15079
rect 6227 15045 6236 15079
rect 6184 15036 6236 15045
rect 6460 15036 6512 15088
rect 7656 15036 7708 15088
rect 8116 15036 8168 15088
rect 8760 15036 8812 15088
rect 6828 14968 6880 15020
rect 7288 14968 7340 15020
rect 7748 14968 7800 15020
rect 8208 14968 8260 15020
rect 9404 15104 9456 15156
rect 9680 15104 9732 15156
rect 9956 15147 10008 15156
rect 9956 15113 9965 15147
rect 9965 15113 9999 15147
rect 9999 15113 10008 15147
rect 9956 15104 10008 15113
rect 10140 15104 10192 15156
rect 10416 15104 10468 15156
rect 11336 15147 11388 15156
rect 10968 15079 11020 15088
rect 10968 15045 10977 15079
rect 10977 15045 11011 15079
rect 11011 15045 11020 15079
rect 10968 15036 11020 15045
rect 11336 15113 11345 15147
rect 11345 15113 11379 15147
rect 11379 15113 11388 15147
rect 11336 15104 11388 15113
rect 12072 15104 12124 15156
rect 11796 15036 11848 15088
rect 13636 15104 13688 15156
rect 14556 15104 14608 15156
rect 15568 15147 15620 15156
rect 15568 15113 15577 15147
rect 15577 15113 15611 15147
rect 15611 15113 15620 15147
rect 15568 15104 15620 15113
rect 14832 15036 14884 15088
rect 15844 15036 15896 15088
rect 11244 14968 11296 15020
rect 12440 14968 12492 15020
rect 14280 15011 14332 15020
rect 5172 14900 5224 14952
rect 5724 14943 5776 14952
rect 5724 14909 5733 14943
rect 5733 14909 5767 14943
rect 5767 14909 5776 14943
rect 5724 14900 5776 14909
rect 5908 14943 5960 14952
rect 5908 14909 5917 14943
rect 5917 14909 5951 14943
rect 5951 14909 5960 14943
rect 5908 14900 5960 14909
rect 7104 14943 7156 14952
rect 7104 14909 7113 14943
rect 7113 14909 7147 14943
rect 7147 14909 7156 14943
rect 7104 14900 7156 14909
rect 7564 14900 7616 14952
rect 2412 14832 2464 14884
rect 3240 14832 3292 14884
rect 5540 14832 5592 14884
rect 5632 14832 5684 14884
rect 7748 14832 7800 14884
rect 7932 14832 7984 14884
rect 8116 14900 8168 14952
rect 9312 14943 9364 14952
rect 9312 14909 9321 14943
rect 9321 14909 9355 14943
rect 9355 14909 9364 14943
rect 9312 14900 9364 14909
rect 10140 14943 10192 14952
rect 10140 14909 10149 14943
rect 10149 14909 10183 14943
rect 10183 14909 10192 14943
rect 10140 14900 10192 14909
rect 8668 14832 8720 14884
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 1676 14764 1728 14816
rect 2504 14764 2556 14816
rect 3148 14807 3200 14816
rect 3148 14773 3157 14807
rect 3157 14773 3191 14807
rect 3191 14773 3200 14807
rect 3148 14764 3200 14773
rect 3608 14764 3660 14816
rect 4344 14764 4396 14816
rect 6460 14764 6512 14816
rect 8392 14764 8444 14816
rect 8576 14764 8628 14816
rect 9956 14832 10008 14884
rect 10784 14900 10836 14952
rect 11612 14943 11664 14952
rect 11612 14909 11621 14943
rect 11621 14909 11655 14943
rect 11655 14909 11664 14943
rect 11612 14900 11664 14909
rect 11796 14943 11848 14952
rect 11796 14909 11805 14943
rect 11805 14909 11839 14943
rect 11839 14909 11848 14943
rect 11796 14900 11848 14909
rect 12072 14900 12124 14952
rect 11980 14832 12032 14884
rect 12624 14900 12676 14952
rect 12992 14900 13044 14952
rect 13728 14900 13780 14952
rect 14280 14977 14289 15011
rect 14289 14977 14323 15011
rect 14323 14977 14332 15011
rect 14280 14968 14332 14977
rect 15660 14968 15712 15020
rect 9680 14764 9732 14816
rect 10416 14807 10468 14816
rect 10416 14773 10425 14807
rect 10425 14773 10459 14807
rect 10459 14773 10468 14807
rect 10416 14764 10468 14773
rect 10508 14764 10560 14816
rect 12440 14764 12492 14816
rect 14832 14900 14884 14952
rect 2824 14662 2876 14714
rect 2888 14662 2940 14714
rect 2952 14662 3004 14714
rect 3016 14662 3068 14714
rect 3080 14662 3132 14714
rect 6572 14662 6624 14714
rect 6636 14662 6688 14714
rect 6700 14662 6752 14714
rect 6764 14662 6816 14714
rect 6828 14662 6880 14714
rect 10320 14662 10372 14714
rect 10384 14662 10436 14714
rect 10448 14662 10500 14714
rect 10512 14662 10564 14714
rect 10576 14662 10628 14714
rect 14068 14662 14120 14714
rect 14132 14662 14184 14714
rect 14196 14662 14248 14714
rect 14260 14662 14312 14714
rect 14324 14662 14376 14714
rect 1584 14560 1636 14612
rect 5080 14603 5132 14612
rect 5080 14569 5089 14603
rect 5089 14569 5123 14603
rect 5123 14569 5132 14603
rect 5080 14560 5132 14569
rect 5724 14560 5776 14612
rect 7012 14603 7064 14612
rect 7012 14569 7021 14603
rect 7021 14569 7055 14603
rect 7055 14569 7064 14603
rect 7012 14560 7064 14569
rect 7288 14603 7340 14612
rect 7288 14569 7297 14603
rect 7297 14569 7331 14603
rect 7331 14569 7340 14603
rect 7288 14560 7340 14569
rect 7656 14560 7708 14612
rect 2596 14492 2648 14544
rect 3056 14424 3108 14476
rect 3792 14424 3844 14476
rect 8300 14560 8352 14612
rect 8760 14560 8812 14612
rect 9220 14560 9272 14612
rect 11428 14560 11480 14612
rect 12440 14560 12492 14612
rect 5908 14424 5960 14476
rect 6368 14424 6420 14476
rect 7840 14467 7892 14476
rect 7840 14433 7849 14467
rect 7849 14433 7883 14467
rect 7883 14433 7892 14467
rect 7840 14424 7892 14433
rect 2688 14356 2740 14408
rect 3148 14399 3200 14408
rect 3148 14365 3157 14399
rect 3157 14365 3191 14399
rect 3191 14365 3200 14399
rect 3148 14356 3200 14365
rect 4436 14356 4488 14408
rect 5356 14356 5408 14408
rect 5632 14356 5684 14408
rect 6276 14399 6328 14408
rect 6276 14365 6285 14399
rect 6285 14365 6319 14399
rect 6319 14365 6328 14399
rect 6276 14356 6328 14365
rect 9036 14424 9088 14476
rect 9128 14424 9180 14476
rect 8852 14356 8904 14408
rect 3516 14263 3568 14272
rect 3516 14229 3525 14263
rect 3525 14229 3559 14263
rect 3559 14229 3568 14263
rect 3516 14220 3568 14229
rect 5724 14288 5776 14340
rect 6000 14288 6052 14340
rect 6184 14288 6236 14340
rect 4160 14263 4212 14272
rect 4160 14229 4169 14263
rect 4169 14229 4203 14263
rect 4203 14229 4212 14263
rect 4160 14220 4212 14229
rect 4252 14263 4304 14272
rect 4252 14229 4261 14263
rect 4261 14229 4295 14263
rect 4295 14229 4304 14263
rect 6828 14288 6880 14340
rect 6920 14288 6972 14340
rect 11520 14492 11572 14544
rect 11980 14492 12032 14544
rect 13360 14560 13412 14612
rect 14372 14492 14424 14544
rect 9404 14424 9456 14476
rect 9956 14424 10008 14476
rect 11244 14424 11296 14476
rect 4252 14220 4304 14229
rect 6460 14220 6512 14272
rect 7472 14220 7524 14272
rect 10692 14288 10744 14340
rect 12532 14356 12584 14408
rect 12900 14331 12952 14340
rect 12900 14297 12918 14331
rect 12918 14297 12952 14331
rect 12900 14288 12952 14297
rect 13084 14288 13136 14340
rect 13636 14356 13688 14408
rect 15016 14356 15068 14408
rect 15476 14356 15528 14408
rect 16212 14356 16264 14408
rect 15752 14288 15804 14340
rect 15936 14288 15988 14340
rect 8944 14220 8996 14272
rect 9772 14263 9824 14272
rect 9772 14229 9781 14263
rect 9781 14229 9815 14263
rect 9815 14229 9824 14263
rect 9772 14220 9824 14229
rect 9956 14263 10008 14272
rect 9956 14229 9965 14263
rect 9965 14229 9999 14263
rect 9999 14229 10008 14263
rect 9956 14220 10008 14229
rect 10784 14220 10836 14272
rect 11796 14263 11848 14272
rect 11796 14229 11805 14263
rect 11805 14229 11839 14263
rect 11839 14229 11848 14263
rect 11796 14220 11848 14229
rect 11980 14220 12032 14272
rect 14280 14263 14332 14272
rect 14280 14229 14289 14263
rect 14289 14229 14323 14263
rect 14323 14229 14332 14263
rect 14280 14220 14332 14229
rect 15476 14220 15528 14272
rect 4698 14118 4750 14170
rect 4762 14118 4814 14170
rect 4826 14118 4878 14170
rect 4890 14118 4942 14170
rect 4954 14118 5006 14170
rect 8446 14118 8498 14170
rect 8510 14118 8562 14170
rect 8574 14118 8626 14170
rect 8638 14118 8690 14170
rect 8702 14118 8754 14170
rect 12194 14118 12246 14170
rect 12258 14118 12310 14170
rect 12322 14118 12374 14170
rect 12386 14118 12438 14170
rect 12450 14118 12502 14170
rect 1032 14016 1084 14068
rect 2780 13948 2832 14000
rect 2872 13948 2924 14000
rect 3424 13991 3476 14000
rect 3424 13957 3433 13991
rect 3433 13957 3467 13991
rect 3467 13957 3476 13991
rect 3424 13948 3476 13957
rect 4252 13991 4304 14000
rect 4252 13957 4261 13991
rect 4261 13957 4295 13991
rect 4295 13957 4304 13991
rect 4252 13948 4304 13957
rect 5448 14016 5500 14068
rect 7656 14016 7708 14068
rect 8024 14059 8076 14068
rect 8024 14025 8033 14059
rect 8033 14025 8067 14059
rect 8067 14025 8076 14059
rect 8024 14016 8076 14025
rect 8208 14016 8260 14068
rect 5172 13948 5224 14000
rect 6828 13948 6880 14000
rect 7564 13948 7616 14000
rect 8116 13948 8168 14000
rect 9036 14016 9088 14068
rect 10692 14016 10744 14068
rect 13728 14059 13780 14068
rect 13728 14025 13737 14059
rect 13737 14025 13771 14059
rect 13771 14025 13780 14059
rect 13728 14016 13780 14025
rect 10968 13991 11020 14000
rect 10968 13957 10977 13991
rect 10977 13957 11011 13991
rect 11011 13957 11020 13991
rect 10968 13948 11020 13957
rect 1676 13923 1728 13932
rect 1676 13889 1685 13923
rect 1685 13889 1719 13923
rect 1719 13889 1728 13923
rect 1676 13880 1728 13889
rect 1400 13812 1452 13864
rect 5816 13923 5868 13932
rect 5816 13889 5834 13923
rect 5834 13889 5868 13923
rect 5816 13880 5868 13889
rect 6000 13880 6052 13932
rect 6460 13880 6512 13932
rect 8944 13880 8996 13932
rect 9956 13880 10008 13932
rect 13084 13948 13136 14000
rect 13820 13991 13872 14000
rect 13820 13957 13829 13991
rect 13829 13957 13863 13991
rect 13863 13957 13872 13991
rect 13820 13948 13872 13957
rect 15476 13991 15528 14000
rect 15476 13957 15485 13991
rect 15485 13957 15519 13991
rect 15519 13957 15528 13991
rect 15476 13948 15528 13957
rect 2228 13812 2280 13864
rect 2872 13812 2924 13864
rect 3792 13812 3844 13864
rect 4160 13812 4212 13864
rect 12808 13880 12860 13932
rect 13360 13923 13412 13932
rect 13360 13889 13369 13923
rect 13369 13889 13403 13923
rect 13403 13889 13412 13923
rect 13360 13880 13412 13889
rect 13176 13855 13228 13864
rect 1492 13787 1544 13796
rect 1492 13753 1501 13787
rect 1501 13753 1535 13787
rect 1535 13753 1544 13787
rect 1492 13744 1544 13753
rect 2320 13719 2372 13728
rect 2320 13685 2329 13719
rect 2329 13685 2363 13719
rect 2363 13685 2372 13719
rect 2320 13676 2372 13685
rect 4528 13719 4580 13728
rect 4528 13685 4537 13719
rect 4537 13685 4571 13719
rect 4571 13685 4580 13719
rect 4528 13676 4580 13685
rect 9956 13744 10008 13796
rect 9864 13676 9916 13728
rect 13176 13821 13185 13855
rect 13185 13821 13219 13855
rect 13219 13821 13228 13855
rect 13176 13812 13228 13821
rect 13728 13812 13780 13864
rect 15660 13855 15712 13864
rect 15660 13821 15669 13855
rect 15669 13821 15703 13855
rect 15703 13821 15712 13855
rect 15660 13812 15712 13821
rect 11428 13744 11480 13796
rect 11336 13719 11388 13728
rect 11336 13685 11345 13719
rect 11345 13685 11379 13719
rect 11379 13685 11388 13719
rect 11336 13676 11388 13685
rect 11796 13676 11848 13728
rect 14648 13744 14700 13796
rect 12900 13719 12952 13728
rect 12900 13685 12909 13719
rect 12909 13685 12943 13719
rect 12943 13685 12952 13719
rect 12900 13676 12952 13685
rect 14372 13676 14424 13728
rect 15476 13676 15528 13728
rect 2824 13574 2876 13626
rect 2888 13574 2940 13626
rect 2952 13574 3004 13626
rect 3016 13574 3068 13626
rect 3080 13574 3132 13626
rect 6572 13574 6624 13626
rect 6636 13574 6688 13626
rect 6700 13574 6752 13626
rect 6764 13574 6816 13626
rect 6828 13574 6880 13626
rect 10320 13574 10372 13626
rect 10384 13574 10436 13626
rect 10448 13574 10500 13626
rect 10512 13574 10564 13626
rect 10576 13574 10628 13626
rect 14068 13574 14120 13626
rect 14132 13574 14184 13626
rect 14196 13574 14248 13626
rect 14260 13574 14312 13626
rect 14324 13574 14376 13626
rect 3148 13472 3200 13524
rect 4068 13472 4120 13524
rect 5908 13472 5960 13524
rect 6276 13472 6328 13524
rect 9128 13515 9180 13524
rect 9128 13481 9137 13515
rect 9137 13481 9171 13515
rect 9171 13481 9180 13515
rect 9128 13472 9180 13481
rect 9772 13515 9824 13524
rect 9772 13481 9781 13515
rect 9781 13481 9815 13515
rect 9815 13481 9824 13515
rect 9772 13472 9824 13481
rect 11612 13472 11664 13524
rect 11980 13472 12032 13524
rect 12808 13472 12860 13524
rect 13084 13515 13136 13524
rect 9036 13404 9088 13456
rect 9680 13404 9732 13456
rect 3148 13336 3200 13388
rect 3424 13379 3476 13388
rect 3424 13345 3433 13379
rect 3433 13345 3467 13379
rect 3467 13345 3476 13379
rect 3424 13336 3476 13345
rect 11152 13404 11204 13456
rect 13084 13481 13093 13515
rect 13093 13481 13127 13515
rect 13127 13481 13136 13515
rect 13084 13472 13136 13481
rect 13360 13472 13412 13524
rect 13728 13472 13780 13524
rect 14648 13379 14700 13388
rect 2320 13268 2372 13320
rect 3516 13268 3568 13320
rect 4528 13268 4580 13320
rect 6000 13268 6052 13320
rect 7656 13311 7708 13320
rect 7656 13277 7690 13311
rect 7690 13277 7708 13311
rect 7656 13268 7708 13277
rect 10140 13311 10192 13320
rect 10140 13277 10174 13311
rect 10174 13277 10192 13311
rect 10140 13268 10192 13277
rect 11612 13268 11664 13320
rect 14648 13345 14657 13379
rect 14657 13345 14691 13379
rect 14691 13345 14700 13379
rect 14648 13336 14700 13345
rect 14556 13311 14608 13320
rect 14556 13277 14565 13311
rect 14565 13277 14599 13311
rect 14599 13277 14608 13311
rect 14556 13268 14608 13277
rect 15752 13268 15804 13320
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 2320 13175 2372 13184
rect 2320 13141 2329 13175
rect 2329 13141 2363 13175
rect 2363 13141 2372 13175
rect 2320 13132 2372 13141
rect 3792 13200 3844 13252
rect 6644 13200 6696 13252
rect 6368 13132 6420 13184
rect 12624 13200 12676 13252
rect 12808 13200 12860 13252
rect 13360 13200 13412 13252
rect 14372 13200 14424 13252
rect 15108 13200 15160 13252
rect 15476 13200 15528 13252
rect 10048 13132 10100 13184
rect 10784 13132 10836 13184
rect 10968 13132 11020 13184
rect 12072 13132 12124 13184
rect 14096 13175 14148 13184
rect 14096 13141 14105 13175
rect 14105 13141 14139 13175
rect 14139 13141 14148 13175
rect 14096 13132 14148 13141
rect 14188 13132 14240 13184
rect 4698 13030 4750 13082
rect 4762 13030 4814 13082
rect 4826 13030 4878 13082
rect 4890 13030 4942 13082
rect 4954 13030 5006 13082
rect 8446 13030 8498 13082
rect 8510 13030 8562 13082
rect 8574 13030 8626 13082
rect 8638 13030 8690 13082
rect 8702 13030 8754 13082
rect 12194 13030 12246 13082
rect 12258 13030 12310 13082
rect 12322 13030 12374 13082
rect 12386 13030 12438 13082
rect 12450 13030 12502 13082
rect 2320 12928 2372 12980
rect 3424 12928 3476 12980
rect 2504 12792 2556 12844
rect 3148 12792 3200 12844
rect 3792 12860 3844 12912
rect 4068 12860 4120 12912
rect 4160 12792 4212 12844
rect 4804 12767 4856 12776
rect 4804 12733 4813 12767
rect 4813 12733 4847 12767
rect 4847 12733 4856 12767
rect 4804 12724 4856 12733
rect 6644 12928 6696 12980
rect 9128 12928 9180 12980
rect 10048 12928 10100 12980
rect 10600 12928 10652 12980
rect 10784 12928 10836 12980
rect 11152 12928 11204 12980
rect 12348 12928 12400 12980
rect 12716 12928 12768 12980
rect 13268 12971 13320 12980
rect 13268 12937 13277 12971
rect 13277 12937 13311 12971
rect 13311 12937 13320 12971
rect 13268 12928 13320 12937
rect 14740 12971 14792 12980
rect 14740 12937 14749 12971
rect 14749 12937 14783 12971
rect 14783 12937 14792 12971
rect 14740 12928 14792 12937
rect 15108 12928 15160 12980
rect 16120 12928 16172 12980
rect 9772 12860 9824 12912
rect 9312 12792 9364 12844
rect 10968 12860 11020 12912
rect 13084 12860 13136 12912
rect 14372 12860 14424 12912
rect 11612 12792 11664 12844
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 14740 12792 14792 12844
rect 14924 12792 14976 12844
rect 15200 12835 15252 12844
rect 15200 12801 15209 12835
rect 15209 12801 15243 12835
rect 15243 12801 15252 12835
rect 15200 12792 15252 12801
rect 15568 12792 15620 12844
rect 11428 12724 11480 12776
rect 12900 12724 12952 12776
rect 3424 12656 3476 12708
rect 8852 12656 8904 12708
rect 9312 12656 9364 12708
rect 10784 12656 10836 12708
rect 14188 12699 14240 12708
rect 14188 12665 14197 12699
rect 14197 12665 14231 12699
rect 14231 12665 14240 12699
rect 14188 12656 14240 12665
rect 14924 12656 14976 12708
rect 15660 12699 15712 12708
rect 15660 12665 15669 12699
rect 15669 12665 15703 12699
rect 15703 12665 15712 12699
rect 15660 12656 15712 12665
rect 9036 12631 9088 12640
rect 9036 12597 9045 12631
rect 9045 12597 9079 12631
rect 9079 12597 9088 12631
rect 9036 12588 9088 12597
rect 9496 12588 9548 12640
rect 9772 12588 9824 12640
rect 13176 12588 13228 12640
rect 2824 12486 2876 12538
rect 2888 12486 2940 12538
rect 2952 12486 3004 12538
rect 3016 12486 3068 12538
rect 3080 12486 3132 12538
rect 6572 12486 6624 12538
rect 6636 12486 6688 12538
rect 6700 12486 6752 12538
rect 6764 12486 6816 12538
rect 6828 12486 6880 12538
rect 10320 12486 10372 12538
rect 10384 12486 10436 12538
rect 10448 12486 10500 12538
rect 10512 12486 10564 12538
rect 10576 12486 10628 12538
rect 14068 12486 14120 12538
rect 14132 12486 14184 12538
rect 14196 12486 14248 12538
rect 14260 12486 14312 12538
rect 14324 12486 14376 12538
rect 3148 12384 3200 12436
rect 6368 12384 6420 12436
rect 7840 12384 7892 12436
rect 10876 12427 10928 12436
rect 10876 12393 10885 12427
rect 10885 12393 10919 12427
rect 10919 12393 10928 12427
rect 10876 12384 10928 12393
rect 13820 12384 13872 12436
rect 15568 12427 15620 12436
rect 15568 12393 15577 12427
rect 15577 12393 15611 12427
rect 15611 12393 15620 12427
rect 15568 12384 15620 12393
rect 3700 12316 3752 12368
rect 5264 12316 5316 12368
rect 11060 12316 11112 12368
rect 12900 12316 12952 12368
rect 4160 12248 4212 12300
rect 15844 12316 15896 12368
rect 3884 12223 3936 12232
rect 3884 12189 3893 12223
rect 3893 12189 3927 12223
rect 3927 12189 3936 12223
rect 3884 12180 3936 12189
rect 4804 12180 4856 12232
rect 6460 12180 6512 12232
rect 4528 12112 4580 12164
rect 9496 12180 9548 12232
rect 13084 12248 13136 12300
rect 10876 12180 10928 12232
rect 11336 12180 11388 12232
rect 13452 12248 13504 12300
rect 14556 12291 14608 12300
rect 14556 12257 14565 12291
rect 14565 12257 14599 12291
rect 14599 12257 14608 12291
rect 14556 12248 14608 12257
rect 14924 12248 14976 12300
rect 15936 12248 15988 12300
rect 1860 12087 1912 12096
rect 1860 12053 1869 12087
rect 1869 12053 1903 12087
rect 1903 12053 1912 12087
rect 1860 12044 1912 12053
rect 2044 12044 2096 12096
rect 2320 12087 2372 12096
rect 2320 12053 2329 12087
rect 2329 12053 2363 12087
rect 2363 12053 2372 12087
rect 2320 12044 2372 12053
rect 3240 12087 3292 12096
rect 3240 12053 3249 12087
rect 3249 12053 3283 12087
rect 3283 12053 3292 12087
rect 3240 12044 3292 12053
rect 3976 12044 4028 12096
rect 5724 12044 5776 12096
rect 9220 12112 9272 12164
rect 11796 12112 11848 12164
rect 12348 12155 12400 12164
rect 12348 12121 12366 12155
rect 12366 12121 12400 12155
rect 12348 12112 12400 12121
rect 14648 12180 14700 12232
rect 11244 12087 11296 12096
rect 11244 12053 11253 12087
rect 11253 12053 11287 12087
rect 11287 12053 11296 12087
rect 11244 12044 11296 12053
rect 11336 12044 11388 12096
rect 12808 12087 12860 12096
rect 12808 12053 12817 12087
rect 12817 12053 12851 12087
rect 12851 12053 12860 12087
rect 12808 12044 12860 12053
rect 13728 12087 13780 12096
rect 13728 12053 13737 12087
rect 13737 12053 13771 12087
rect 13771 12053 13780 12087
rect 13728 12044 13780 12053
rect 4698 11942 4750 11994
rect 4762 11942 4814 11994
rect 4826 11942 4878 11994
rect 4890 11942 4942 11994
rect 4954 11942 5006 11994
rect 8446 11942 8498 11994
rect 8510 11942 8562 11994
rect 8574 11942 8626 11994
rect 8638 11942 8690 11994
rect 8702 11942 8754 11994
rect 12194 11942 12246 11994
rect 12258 11942 12310 11994
rect 12322 11942 12374 11994
rect 12386 11942 12438 11994
rect 12450 11942 12502 11994
rect 1492 11883 1544 11892
rect 1492 11849 1501 11883
rect 1501 11849 1535 11883
rect 1535 11849 1544 11883
rect 1492 11840 1544 11849
rect 2596 11883 2648 11892
rect 2596 11849 2605 11883
rect 2605 11849 2639 11883
rect 2639 11849 2648 11883
rect 2596 11840 2648 11849
rect 4160 11840 4212 11892
rect 4344 11840 4396 11892
rect 9496 11883 9548 11892
rect 2412 11772 2464 11824
rect 2320 11704 2372 11756
rect 3148 11704 3200 11756
rect 3976 11772 4028 11824
rect 4528 11772 4580 11824
rect 9496 11849 9505 11883
rect 9505 11849 9539 11883
rect 9539 11849 9548 11883
rect 9496 11840 9548 11849
rect 9956 11840 10008 11892
rect 11336 11840 11388 11892
rect 11704 11840 11756 11892
rect 12992 11883 13044 11892
rect 12992 11849 13001 11883
rect 13001 11849 13035 11883
rect 13035 11849 13044 11883
rect 12992 11840 13044 11849
rect 13176 11883 13228 11892
rect 13176 11849 13185 11883
rect 13185 11849 13219 11883
rect 13219 11849 13228 11883
rect 13176 11840 13228 11849
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 14464 11840 14516 11892
rect 14740 11883 14792 11892
rect 14740 11849 14749 11883
rect 14749 11849 14783 11883
rect 14783 11849 14792 11883
rect 14740 11840 14792 11849
rect 15292 11840 15344 11892
rect 4068 11704 4120 11756
rect 10232 11704 10284 11756
rect 11244 11772 11296 11824
rect 3516 11679 3568 11688
rect 3516 11645 3525 11679
rect 3525 11645 3559 11679
rect 3559 11645 3568 11679
rect 3516 11636 3568 11645
rect 5448 11679 5500 11688
rect 5448 11645 5457 11679
rect 5457 11645 5491 11679
rect 5491 11645 5500 11679
rect 10876 11679 10928 11688
rect 5448 11636 5500 11645
rect 2136 11543 2188 11552
rect 2136 11509 2145 11543
rect 2145 11509 2179 11543
rect 2179 11509 2188 11543
rect 2136 11500 2188 11509
rect 2504 11500 2556 11552
rect 3240 11500 3292 11552
rect 10876 11645 10885 11679
rect 10885 11645 10919 11679
rect 10919 11645 10928 11679
rect 10876 11636 10928 11645
rect 12624 11704 12676 11756
rect 12716 11704 12768 11756
rect 12072 11636 12124 11688
rect 13544 11772 13596 11824
rect 15752 11772 15804 11824
rect 13820 11568 13872 11620
rect 14648 11636 14700 11688
rect 9220 11500 9272 11552
rect 11060 11500 11112 11552
rect 13360 11543 13412 11552
rect 13360 11509 13369 11543
rect 13369 11509 13403 11543
rect 13403 11509 13412 11543
rect 13360 11500 13412 11509
rect 13912 11500 13964 11552
rect 16028 11704 16080 11756
rect 15200 11500 15252 11552
rect 2824 11398 2876 11450
rect 2888 11398 2940 11450
rect 2952 11398 3004 11450
rect 3016 11398 3068 11450
rect 3080 11398 3132 11450
rect 6572 11398 6624 11450
rect 6636 11398 6688 11450
rect 6700 11398 6752 11450
rect 6764 11398 6816 11450
rect 6828 11398 6880 11450
rect 10320 11398 10372 11450
rect 10384 11398 10436 11450
rect 10448 11398 10500 11450
rect 10512 11398 10564 11450
rect 10576 11398 10628 11450
rect 14068 11398 14120 11450
rect 14132 11398 14184 11450
rect 14196 11398 14248 11450
rect 14260 11398 14312 11450
rect 14324 11398 14376 11450
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 5816 11339 5868 11348
rect 1768 11092 1820 11144
rect 2504 11203 2556 11212
rect 2504 11169 2513 11203
rect 2513 11169 2547 11203
rect 2547 11169 2556 11203
rect 2504 11160 2556 11169
rect 5816 11305 5825 11339
rect 5825 11305 5859 11339
rect 5859 11305 5868 11339
rect 5816 11296 5868 11305
rect 7288 11339 7340 11348
rect 7288 11305 7297 11339
rect 7297 11305 7331 11339
rect 7331 11305 7340 11339
rect 7288 11296 7340 11305
rect 9496 11296 9548 11348
rect 10140 11296 10192 11348
rect 2596 11092 2648 11144
rect 3516 11203 3568 11212
rect 3516 11169 3525 11203
rect 3525 11169 3559 11203
rect 3559 11169 3568 11203
rect 4068 11228 4120 11280
rect 3516 11160 3568 11169
rect 4344 11160 4396 11212
rect 3976 11092 4028 11144
rect 5448 11092 5500 11144
rect 6092 11024 6144 11076
rect 8852 11024 8904 11076
rect 9220 11092 9272 11144
rect 10876 11296 10928 11348
rect 12532 11296 12584 11348
rect 15292 11296 15344 11348
rect 16304 11296 16356 11348
rect 14648 11203 14700 11212
rect 14648 11169 14657 11203
rect 14657 11169 14691 11203
rect 14691 11169 14700 11203
rect 14648 11160 14700 11169
rect 15200 11160 15252 11212
rect 9588 11024 9640 11076
rect 16028 11092 16080 11144
rect 1492 10999 1544 11008
rect 1492 10965 1501 10999
rect 1501 10965 1535 10999
rect 1535 10965 1544 10999
rect 1492 10956 1544 10965
rect 3148 10956 3200 11008
rect 3332 10956 3384 11008
rect 8944 10999 8996 11008
rect 8944 10965 8953 10999
rect 8953 10965 8987 10999
rect 8987 10965 8996 10999
rect 8944 10956 8996 10965
rect 9312 10956 9364 11008
rect 9956 10956 10008 11008
rect 11888 10956 11940 11008
rect 14556 11067 14608 11076
rect 14556 11033 14565 11067
rect 14565 11033 14599 11067
rect 14599 11033 14608 11067
rect 14556 11024 14608 11033
rect 15200 11024 15252 11076
rect 15384 11024 15436 11076
rect 12072 10999 12124 11008
rect 12072 10965 12081 10999
rect 12081 10965 12115 10999
rect 12115 10965 12124 10999
rect 14096 10999 14148 11008
rect 12072 10956 12124 10965
rect 14096 10965 14105 10999
rect 14105 10965 14139 10999
rect 14139 10965 14148 10999
rect 14096 10956 14148 10965
rect 14648 10956 14700 11008
rect 15016 10956 15068 11008
rect 4698 10854 4750 10906
rect 4762 10854 4814 10906
rect 4826 10854 4878 10906
rect 4890 10854 4942 10906
rect 4954 10854 5006 10906
rect 8446 10854 8498 10906
rect 8510 10854 8562 10906
rect 8574 10854 8626 10906
rect 8638 10854 8690 10906
rect 8702 10854 8754 10906
rect 12194 10854 12246 10906
rect 12258 10854 12310 10906
rect 12322 10854 12374 10906
rect 12386 10854 12438 10906
rect 12450 10854 12502 10906
rect 1860 10795 1912 10804
rect 1860 10761 1869 10795
rect 1869 10761 1903 10795
rect 1903 10761 1912 10795
rect 1860 10752 1912 10761
rect 2136 10752 2188 10804
rect 4344 10795 4396 10804
rect 4344 10761 4353 10795
rect 4353 10761 4387 10795
rect 4387 10761 4396 10795
rect 4344 10752 4396 10761
rect 4528 10752 4580 10804
rect 6092 10752 6144 10804
rect 9956 10752 10008 10804
rect 10692 10752 10744 10804
rect 12532 10795 12584 10804
rect 12532 10761 12541 10795
rect 12541 10761 12575 10795
rect 12575 10761 12584 10795
rect 12532 10752 12584 10761
rect 13360 10752 13412 10804
rect 4068 10684 4120 10736
rect 5632 10684 5684 10736
rect 5816 10727 5868 10736
rect 5816 10693 5834 10727
rect 5834 10693 5868 10727
rect 5816 10684 5868 10693
rect 11060 10684 11112 10736
rect 12808 10684 12860 10736
rect 14096 10684 14148 10736
rect 2596 10548 2648 10600
rect 7104 10616 7156 10668
rect 7564 10659 7616 10668
rect 7564 10625 7582 10659
rect 7582 10625 7616 10659
rect 7564 10616 7616 10625
rect 9680 10616 9732 10668
rect 10048 10616 10100 10668
rect 3148 10548 3200 10600
rect 3516 10548 3568 10600
rect 4160 10591 4212 10600
rect 4160 10557 4169 10591
rect 4169 10557 4203 10591
rect 4203 10557 4212 10591
rect 4160 10548 4212 10557
rect 4344 10548 4396 10600
rect 4620 10548 4672 10600
rect 8944 10591 8996 10600
rect 4436 10480 4488 10532
rect 1676 10412 1728 10464
rect 5908 10412 5960 10464
rect 8944 10557 8953 10591
rect 8953 10557 8987 10591
rect 8987 10557 8996 10591
rect 8944 10548 8996 10557
rect 11888 10591 11940 10600
rect 11888 10557 11897 10591
rect 11897 10557 11931 10591
rect 11931 10557 11940 10591
rect 11888 10548 11940 10557
rect 8024 10455 8076 10464
rect 8024 10421 8033 10455
rect 8033 10421 8067 10455
rect 8067 10421 8076 10455
rect 8024 10412 8076 10421
rect 12624 10480 12676 10532
rect 12716 10480 12768 10532
rect 10784 10412 10836 10464
rect 15292 10412 15344 10464
rect 15936 10412 15988 10464
rect 2824 10310 2876 10362
rect 2888 10310 2940 10362
rect 2952 10310 3004 10362
rect 3016 10310 3068 10362
rect 3080 10310 3132 10362
rect 6572 10310 6624 10362
rect 6636 10310 6688 10362
rect 6700 10310 6752 10362
rect 6764 10310 6816 10362
rect 6828 10310 6880 10362
rect 10320 10310 10372 10362
rect 10384 10310 10436 10362
rect 10448 10310 10500 10362
rect 10512 10310 10564 10362
rect 10576 10310 10628 10362
rect 14068 10310 14120 10362
rect 14132 10310 14184 10362
rect 14196 10310 14248 10362
rect 14260 10310 14312 10362
rect 14324 10310 14376 10362
rect 1768 10251 1820 10260
rect 1768 10217 1777 10251
rect 1777 10217 1811 10251
rect 1811 10217 1820 10251
rect 1768 10208 1820 10217
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 2412 10140 2464 10192
rect 3516 10140 3568 10192
rect 4252 10072 4304 10124
rect 10784 10208 10836 10260
rect 3516 10004 3568 10056
rect 4160 10004 4212 10056
rect 1492 9911 1544 9920
rect 1492 9877 1501 9911
rect 1501 9877 1535 9911
rect 1535 9877 1544 9911
rect 1492 9868 1544 9877
rect 1952 9868 2004 9920
rect 2320 9868 2372 9920
rect 2504 9911 2556 9920
rect 2504 9877 2513 9911
rect 2513 9877 2547 9911
rect 2547 9877 2556 9911
rect 5908 10004 5960 10056
rect 7196 10004 7248 10056
rect 11152 10072 11204 10124
rect 15108 10115 15160 10124
rect 15108 10081 15117 10115
rect 15117 10081 15151 10115
rect 15151 10081 15160 10115
rect 15108 10072 15160 10081
rect 15016 10047 15068 10056
rect 8024 9936 8076 9988
rect 12072 9936 12124 9988
rect 2504 9868 2556 9877
rect 7288 9868 7340 9920
rect 11612 9868 11664 9920
rect 15016 10013 15025 10047
rect 15025 10013 15059 10047
rect 15059 10013 15068 10047
rect 15016 10004 15068 10013
rect 16212 10004 16264 10056
rect 14280 9936 14332 9988
rect 14464 9936 14516 9988
rect 14832 9936 14884 9988
rect 13084 9911 13136 9920
rect 13084 9877 13093 9911
rect 13093 9877 13127 9911
rect 13127 9877 13136 9911
rect 14556 9911 14608 9920
rect 13084 9868 13136 9877
rect 14556 9877 14565 9911
rect 14565 9877 14599 9911
rect 14599 9877 14608 9911
rect 14556 9868 14608 9877
rect 15568 9911 15620 9920
rect 15568 9877 15577 9911
rect 15577 9877 15611 9911
rect 15611 9877 15620 9911
rect 15568 9868 15620 9877
rect 4698 9766 4750 9818
rect 4762 9766 4814 9818
rect 4826 9766 4878 9818
rect 4890 9766 4942 9818
rect 4954 9766 5006 9818
rect 8446 9766 8498 9818
rect 8510 9766 8562 9818
rect 8574 9766 8626 9818
rect 8638 9766 8690 9818
rect 8702 9766 8754 9818
rect 12194 9766 12246 9818
rect 12258 9766 12310 9818
rect 12322 9766 12374 9818
rect 12386 9766 12438 9818
rect 12450 9766 12502 9818
rect 2504 9664 2556 9716
rect 7196 9664 7248 9716
rect 11152 9664 11204 9716
rect 13084 9664 13136 9716
rect 14280 9707 14332 9716
rect 14280 9673 14289 9707
rect 14289 9673 14323 9707
rect 14323 9673 14332 9707
rect 14280 9664 14332 9673
rect 14556 9664 14608 9716
rect 3884 9596 3936 9648
rect 1676 9571 1728 9580
rect 1676 9537 1685 9571
rect 1685 9537 1719 9571
rect 1719 9537 1728 9571
rect 1676 9528 1728 9537
rect 1952 9571 2004 9580
rect 1952 9537 1961 9571
rect 1961 9537 1995 9571
rect 1995 9537 2004 9571
rect 1952 9528 2004 9537
rect 2412 9528 2464 9580
rect 3332 9528 3384 9580
rect 3516 9528 3568 9580
rect 2504 9460 2556 9512
rect 1860 9392 1912 9444
rect 3792 9460 3844 9512
rect 4068 9528 4120 9580
rect 5908 9528 5960 9580
rect 7840 9596 7892 9648
rect 8116 9596 8168 9648
rect 10140 9596 10192 9648
rect 12532 9596 12584 9648
rect 12808 9528 12860 9580
rect 15016 9596 15068 9648
rect 15384 9596 15436 9648
rect 13820 9528 13872 9580
rect 14924 9528 14976 9580
rect 13636 9503 13688 9512
rect 13636 9469 13645 9503
rect 13645 9469 13679 9503
rect 13679 9469 13688 9503
rect 13636 9460 13688 9469
rect 15292 9503 15344 9512
rect 1492 9367 1544 9376
rect 1492 9333 1501 9367
rect 1501 9333 1535 9367
rect 1535 9333 1544 9367
rect 1492 9324 1544 9333
rect 1768 9367 1820 9376
rect 1768 9333 1777 9367
rect 1777 9333 1811 9367
rect 1811 9333 1820 9367
rect 1768 9324 1820 9333
rect 4252 9367 4304 9376
rect 4252 9333 4261 9367
rect 4261 9333 4295 9367
rect 4295 9333 4304 9367
rect 4252 9324 4304 9333
rect 5908 9324 5960 9376
rect 7564 9324 7616 9376
rect 8024 9367 8076 9376
rect 8024 9333 8033 9367
rect 8033 9333 8067 9367
rect 8067 9333 8076 9367
rect 8024 9324 8076 9333
rect 9588 9324 9640 9376
rect 15292 9469 15301 9503
rect 15301 9469 15335 9503
rect 15335 9469 15344 9503
rect 15292 9460 15344 9469
rect 2824 9222 2876 9274
rect 2888 9222 2940 9274
rect 2952 9222 3004 9274
rect 3016 9222 3068 9274
rect 3080 9222 3132 9274
rect 6572 9222 6624 9274
rect 6636 9222 6688 9274
rect 6700 9222 6752 9274
rect 6764 9222 6816 9274
rect 6828 9222 6880 9274
rect 10320 9222 10372 9274
rect 10384 9222 10436 9274
rect 10448 9222 10500 9274
rect 10512 9222 10564 9274
rect 10576 9222 10628 9274
rect 14068 9222 14120 9274
rect 14132 9222 14184 9274
rect 14196 9222 14248 9274
rect 14260 9222 14312 9274
rect 14324 9222 14376 9274
rect 2412 9163 2464 9172
rect 2412 9129 2421 9163
rect 2421 9129 2455 9163
rect 2455 9129 2464 9163
rect 2412 9120 2464 9129
rect 2596 9120 2648 9172
rect 9772 9120 9824 9172
rect 10048 9163 10100 9172
rect 10048 9129 10057 9163
rect 10057 9129 10091 9163
rect 10091 9129 10100 9163
rect 10048 9120 10100 9129
rect 13636 9120 13688 9172
rect 14924 9163 14976 9172
rect 14924 9129 14933 9163
rect 14933 9129 14967 9163
rect 14967 9129 14976 9163
rect 14924 9120 14976 9129
rect 3884 9052 3936 9104
rect 12808 9052 12860 9104
rect 13912 9052 13964 9104
rect 3516 9027 3568 9036
rect 3516 8993 3525 9027
rect 3525 8993 3559 9027
rect 3559 8993 3568 9027
rect 3516 8984 3568 8993
rect 2688 8916 2740 8968
rect 3700 8916 3752 8968
rect 5908 8959 5960 8968
rect 5908 8925 5917 8959
rect 5917 8925 5951 8959
rect 5951 8925 5960 8959
rect 5908 8916 5960 8925
rect 2872 8848 2924 8900
rect 3148 8848 3200 8900
rect 3332 8780 3384 8832
rect 4344 8848 4396 8900
rect 4528 8780 4580 8832
rect 5724 8780 5776 8832
rect 7932 8780 7984 8832
rect 8024 8780 8076 8832
rect 8852 8780 8904 8832
rect 11612 8916 11664 8968
rect 15108 8984 15160 9036
rect 14924 8916 14976 8968
rect 15292 8959 15344 8968
rect 15292 8925 15301 8959
rect 15301 8925 15335 8959
rect 15335 8925 15344 8959
rect 15292 8916 15344 8925
rect 15384 8959 15436 8968
rect 15384 8925 15393 8959
rect 15393 8925 15427 8959
rect 15427 8925 15436 8959
rect 15384 8916 15436 8925
rect 11888 8848 11940 8900
rect 12716 8848 12768 8900
rect 13176 8780 13228 8832
rect 13728 8823 13780 8832
rect 13728 8789 13737 8823
rect 13737 8789 13771 8823
rect 13771 8789 13780 8823
rect 13728 8780 13780 8789
rect 14464 8823 14516 8832
rect 14464 8789 14473 8823
rect 14473 8789 14507 8823
rect 14507 8789 14516 8823
rect 14464 8780 14516 8789
rect 14556 8823 14608 8832
rect 14556 8789 14565 8823
rect 14565 8789 14599 8823
rect 14599 8789 14608 8823
rect 14556 8780 14608 8789
rect 4698 8678 4750 8730
rect 4762 8678 4814 8730
rect 4826 8678 4878 8730
rect 4890 8678 4942 8730
rect 4954 8678 5006 8730
rect 8446 8678 8498 8730
rect 8510 8678 8562 8730
rect 8574 8678 8626 8730
rect 8638 8678 8690 8730
rect 8702 8678 8754 8730
rect 12194 8678 12246 8730
rect 12258 8678 12310 8730
rect 12322 8678 12374 8730
rect 12386 8678 12438 8730
rect 12450 8678 12502 8730
rect 2320 8576 2372 8628
rect 2504 8619 2556 8628
rect 2504 8585 2513 8619
rect 2513 8585 2547 8619
rect 2547 8585 2556 8619
rect 2872 8619 2924 8628
rect 2504 8576 2556 8585
rect 2872 8585 2881 8619
rect 2881 8585 2915 8619
rect 2915 8585 2924 8619
rect 2872 8576 2924 8585
rect 4068 8576 4120 8628
rect 4344 8576 4396 8628
rect 3148 8508 3200 8560
rect 3240 8508 3292 8560
rect 3516 8508 3568 8560
rect 5908 8576 5960 8628
rect 8024 8576 8076 8628
rect 13728 8576 13780 8628
rect 13820 8619 13872 8628
rect 13820 8585 13829 8619
rect 13829 8585 13863 8619
rect 13863 8585 13872 8619
rect 13820 8576 13872 8585
rect 14556 8576 14608 8628
rect 14648 8576 14700 8628
rect 15384 8619 15436 8628
rect 1860 8415 1912 8424
rect 1860 8381 1869 8415
rect 1869 8381 1903 8415
rect 1903 8381 1912 8415
rect 1860 8372 1912 8381
rect 3884 8440 3936 8492
rect 6276 8508 6328 8560
rect 4252 8440 4304 8492
rect 7380 8440 7432 8492
rect 13544 8440 13596 8492
rect 14648 8440 14700 8492
rect 8852 8415 8904 8424
rect 3240 8304 3292 8356
rect 4068 8304 4120 8356
rect 8852 8381 8861 8415
rect 8861 8381 8895 8415
rect 8895 8381 8904 8415
rect 8852 8372 8904 8381
rect 13912 8372 13964 8424
rect 14556 8372 14608 8424
rect 15384 8585 15393 8619
rect 15393 8585 15427 8619
rect 15427 8585 15436 8619
rect 15384 8576 15436 8585
rect 15476 8508 15528 8560
rect 14924 8415 14976 8424
rect 14924 8381 14933 8415
rect 14933 8381 14967 8415
rect 14967 8381 14976 8415
rect 14924 8372 14976 8381
rect 7472 8347 7524 8356
rect 7472 8313 7481 8347
rect 7481 8313 7515 8347
rect 7515 8313 7524 8347
rect 7472 8304 7524 8313
rect 11612 8304 11664 8356
rect 13176 8304 13228 8356
rect 13820 8304 13872 8356
rect 15200 8304 15252 8356
rect 5172 8236 5224 8288
rect 10784 8236 10836 8288
rect 12716 8279 12768 8288
rect 12716 8245 12725 8279
rect 12725 8245 12759 8279
rect 12759 8245 12768 8279
rect 12716 8236 12768 8245
rect 12992 8236 13044 8288
rect 14556 8236 14608 8288
rect 2824 8134 2876 8186
rect 2888 8134 2940 8186
rect 2952 8134 3004 8186
rect 3016 8134 3068 8186
rect 3080 8134 3132 8186
rect 6572 8134 6624 8186
rect 6636 8134 6688 8186
rect 6700 8134 6752 8186
rect 6764 8134 6816 8186
rect 6828 8134 6880 8186
rect 10320 8134 10372 8186
rect 10384 8134 10436 8186
rect 10448 8134 10500 8186
rect 10512 8134 10564 8186
rect 10576 8134 10628 8186
rect 14068 8134 14120 8186
rect 14132 8134 14184 8186
rect 14196 8134 14248 8186
rect 14260 8134 14312 8186
rect 14324 8134 14376 8186
rect 1492 8075 1544 8084
rect 1492 8041 1501 8075
rect 1501 8041 1535 8075
rect 1535 8041 1544 8075
rect 1492 8032 1544 8041
rect 3148 8032 3200 8084
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 11888 8032 11940 8084
rect 12900 8032 12952 8084
rect 13452 8032 13504 8084
rect 14464 8075 14516 8084
rect 3424 7896 3476 7948
rect 12624 7964 12676 8016
rect 4436 7828 4488 7880
rect 5172 7828 5224 7880
rect 8852 7828 8904 7880
rect 9404 7828 9456 7880
rect 3148 7760 3200 7812
rect 3976 7760 4028 7812
rect 4068 7760 4120 7812
rect 3608 7692 3660 7744
rect 5448 7692 5500 7744
rect 7932 7760 7984 7812
rect 9588 7803 9640 7812
rect 9588 7769 9622 7803
rect 9622 7769 9640 7803
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 14464 8041 14473 8075
rect 14473 8041 14507 8075
rect 14507 8041 14516 8075
rect 14464 8032 14516 8041
rect 14924 7896 14976 7948
rect 13636 7871 13688 7880
rect 9588 7760 9640 7769
rect 12624 7760 12676 7812
rect 13084 7760 13136 7812
rect 13636 7837 13645 7871
rect 13645 7837 13679 7871
rect 13679 7837 13688 7871
rect 13636 7828 13688 7837
rect 13912 7828 13964 7880
rect 14372 7760 14424 7812
rect 13452 7692 13504 7744
rect 13544 7692 13596 7744
rect 14464 7692 14516 7744
rect 14740 7692 14792 7744
rect 15016 7692 15068 7744
rect 15476 7735 15528 7744
rect 15476 7701 15485 7735
rect 15485 7701 15519 7735
rect 15519 7701 15528 7735
rect 15476 7692 15528 7701
rect 15660 7735 15712 7744
rect 15660 7701 15669 7735
rect 15669 7701 15703 7735
rect 15703 7701 15712 7735
rect 15660 7692 15712 7701
rect 4698 7590 4750 7642
rect 4762 7590 4814 7642
rect 4826 7590 4878 7642
rect 4890 7590 4942 7642
rect 4954 7590 5006 7642
rect 8446 7590 8498 7642
rect 8510 7590 8562 7642
rect 8574 7590 8626 7642
rect 8638 7590 8690 7642
rect 8702 7590 8754 7642
rect 12194 7590 12246 7642
rect 12258 7590 12310 7642
rect 12322 7590 12374 7642
rect 12386 7590 12438 7642
rect 12450 7590 12502 7642
rect 1676 7488 1728 7540
rect 2044 7488 2096 7540
rect 13452 7488 13504 7540
rect 15016 7488 15068 7540
rect 3148 7463 3200 7472
rect 3148 7429 3157 7463
rect 3157 7429 3191 7463
rect 3191 7429 3200 7463
rect 3148 7420 3200 7429
rect 2412 7352 2464 7404
rect 3976 7420 4028 7472
rect 5172 7420 5224 7472
rect 4160 7352 4212 7404
rect 5448 7395 5500 7404
rect 5448 7361 5466 7395
rect 5466 7361 5500 7395
rect 5448 7352 5500 7361
rect 5816 7352 5868 7404
rect 2228 7284 2280 7336
rect 3424 7327 3476 7336
rect 2320 7259 2372 7268
rect 2320 7225 2329 7259
rect 2329 7225 2363 7259
rect 2363 7225 2372 7259
rect 2320 7216 2372 7225
rect 3424 7293 3433 7327
rect 3433 7293 3467 7327
rect 3467 7293 3476 7327
rect 3424 7284 3476 7293
rect 3516 7216 3568 7268
rect 4620 7216 4672 7268
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 2504 7191 2556 7200
rect 2504 7157 2513 7191
rect 2513 7157 2547 7191
rect 2547 7157 2556 7191
rect 2504 7148 2556 7157
rect 3240 7148 3292 7200
rect 3608 7148 3660 7200
rect 4344 7191 4396 7200
rect 4344 7157 4353 7191
rect 4353 7157 4387 7191
rect 4387 7157 4396 7191
rect 4344 7148 4396 7157
rect 4436 7148 4488 7200
rect 5448 7148 5500 7200
rect 6460 7148 6512 7200
rect 8392 7352 8444 7404
rect 9312 7395 9364 7404
rect 9312 7361 9330 7395
rect 9330 7361 9364 7395
rect 9588 7395 9640 7404
rect 9312 7352 9364 7361
rect 9588 7361 9597 7395
rect 9597 7361 9631 7395
rect 9631 7361 9640 7395
rect 10784 7420 10836 7472
rect 9588 7352 9640 7361
rect 11152 7352 11204 7404
rect 11612 7420 11664 7472
rect 12716 7420 12768 7472
rect 12900 7420 12952 7472
rect 13360 7395 13412 7404
rect 13360 7361 13369 7395
rect 13369 7361 13403 7395
rect 13403 7361 13412 7395
rect 13360 7352 13412 7361
rect 11520 7327 11572 7336
rect 11520 7293 11529 7327
rect 11529 7293 11563 7327
rect 11563 7293 11572 7327
rect 11520 7284 11572 7293
rect 13452 7327 13504 7336
rect 13452 7293 13461 7327
rect 13461 7293 13495 7327
rect 13495 7293 13504 7327
rect 13452 7284 13504 7293
rect 14556 7420 14608 7472
rect 15384 7488 15436 7540
rect 15844 7488 15896 7540
rect 15108 7395 15160 7404
rect 15108 7361 15117 7395
rect 15117 7361 15151 7395
rect 15151 7361 15160 7395
rect 15108 7352 15160 7361
rect 14372 7327 14424 7336
rect 14372 7293 14381 7327
rect 14381 7293 14415 7327
rect 14415 7293 14424 7327
rect 14372 7284 14424 7293
rect 7012 7148 7064 7200
rect 8116 7191 8168 7200
rect 8116 7157 8125 7191
rect 8125 7157 8159 7191
rect 8159 7157 8168 7191
rect 8116 7148 8168 7157
rect 11336 7191 11388 7200
rect 11336 7157 11345 7191
rect 11345 7157 11379 7191
rect 11379 7157 11388 7191
rect 11336 7148 11388 7157
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 13176 7148 13228 7200
rect 15568 7216 15620 7268
rect 13820 7191 13872 7200
rect 13820 7157 13829 7191
rect 13829 7157 13863 7191
rect 13863 7157 13872 7191
rect 13820 7148 13872 7157
rect 14004 7148 14056 7200
rect 14556 7148 14608 7200
rect 14740 7191 14792 7200
rect 14740 7157 14749 7191
rect 14749 7157 14783 7191
rect 14783 7157 14792 7191
rect 14740 7148 14792 7157
rect 2824 7046 2876 7098
rect 2888 7046 2940 7098
rect 2952 7046 3004 7098
rect 3016 7046 3068 7098
rect 3080 7046 3132 7098
rect 6572 7046 6624 7098
rect 6636 7046 6688 7098
rect 6700 7046 6752 7098
rect 6764 7046 6816 7098
rect 6828 7046 6880 7098
rect 10320 7046 10372 7098
rect 10384 7046 10436 7098
rect 10448 7046 10500 7098
rect 10512 7046 10564 7098
rect 10576 7046 10628 7098
rect 14068 7046 14120 7098
rect 14132 7046 14184 7098
rect 14196 7046 14248 7098
rect 14260 7046 14312 7098
rect 14324 7046 14376 7098
rect 2044 6944 2096 6996
rect 8392 6944 8444 6996
rect 4160 6876 4212 6928
rect 1584 6851 1636 6860
rect 1584 6817 1593 6851
rect 1593 6817 1627 6851
rect 1627 6817 1636 6851
rect 1584 6808 1636 6817
rect 1952 6808 2004 6860
rect 2136 6808 2188 6860
rect 3332 6808 3384 6860
rect 9588 6944 9640 6996
rect 13084 6944 13136 6996
rect 1400 6740 1452 6792
rect 1860 6740 1912 6792
rect 2596 6783 2648 6792
rect 2596 6749 2605 6783
rect 2605 6749 2639 6783
rect 2639 6749 2648 6783
rect 2596 6740 2648 6749
rect 3884 6740 3936 6792
rect 6460 6740 6512 6792
rect 12072 6740 12124 6792
rect 13636 6808 13688 6860
rect 14556 6944 14608 6996
rect 13912 6740 13964 6792
rect 14740 6740 14792 6792
rect 2688 6672 2740 6724
rect 3332 6672 3384 6724
rect 2136 6647 2188 6656
rect 2136 6613 2145 6647
rect 2145 6613 2179 6647
rect 2179 6613 2188 6647
rect 2136 6604 2188 6613
rect 2504 6647 2556 6656
rect 2504 6613 2513 6647
rect 2513 6613 2547 6647
rect 2547 6613 2556 6647
rect 2504 6604 2556 6613
rect 2780 6647 2832 6656
rect 2780 6613 2789 6647
rect 2789 6613 2823 6647
rect 2823 6613 2832 6647
rect 3148 6647 3200 6656
rect 2780 6604 2832 6613
rect 3148 6613 3157 6647
rect 3157 6613 3191 6647
rect 3191 6613 3200 6647
rect 3148 6604 3200 6613
rect 3424 6604 3476 6656
rect 3792 6647 3844 6656
rect 3792 6613 3801 6647
rect 3801 6613 3835 6647
rect 3835 6613 3844 6647
rect 3792 6604 3844 6613
rect 5540 6647 5592 6656
rect 5540 6613 5549 6647
rect 5549 6613 5583 6647
rect 5583 6613 5592 6647
rect 5540 6604 5592 6613
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 11244 6672 11296 6724
rect 11336 6672 11388 6724
rect 12900 6672 12952 6724
rect 13268 6672 13320 6724
rect 13360 6672 13412 6724
rect 15016 6876 15068 6928
rect 14924 6740 14976 6792
rect 15292 6715 15344 6724
rect 7380 6604 7432 6613
rect 9680 6604 9732 6656
rect 11980 6647 12032 6656
rect 11980 6613 11989 6647
rect 11989 6613 12023 6647
rect 12023 6613 12032 6647
rect 11980 6604 12032 6613
rect 13636 6604 13688 6656
rect 15292 6681 15301 6715
rect 15301 6681 15335 6715
rect 15335 6681 15344 6715
rect 15292 6672 15344 6681
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 14740 6604 14792 6656
rect 4698 6502 4750 6554
rect 4762 6502 4814 6554
rect 4826 6502 4878 6554
rect 4890 6502 4942 6554
rect 4954 6502 5006 6554
rect 8446 6502 8498 6554
rect 8510 6502 8562 6554
rect 8574 6502 8626 6554
rect 8638 6502 8690 6554
rect 8702 6502 8754 6554
rect 12194 6502 12246 6554
rect 12258 6502 12310 6554
rect 12322 6502 12374 6554
rect 12386 6502 12438 6554
rect 12450 6502 12502 6554
rect 3792 6400 3844 6452
rect 6276 6400 6328 6452
rect 2780 6332 2832 6384
rect 3516 6332 3568 6384
rect 4344 6332 4396 6384
rect 2228 6307 2280 6316
rect 2228 6273 2237 6307
rect 2237 6273 2271 6307
rect 2271 6273 2280 6307
rect 2228 6264 2280 6273
rect 2596 6264 2648 6316
rect 6460 6332 6512 6384
rect 2780 6196 2832 6248
rect 3240 6196 3292 6248
rect 5540 6264 5592 6316
rect 6000 6264 6052 6316
rect 7932 6400 7984 6452
rect 9956 6400 10008 6452
rect 11428 6400 11480 6452
rect 11520 6400 11572 6452
rect 12072 6400 12124 6452
rect 12164 6400 12216 6452
rect 13820 6400 13872 6452
rect 14556 6443 14608 6452
rect 14556 6409 14565 6443
rect 14565 6409 14599 6443
rect 14599 6409 14608 6443
rect 14556 6400 14608 6409
rect 14832 6400 14884 6452
rect 15752 6400 15804 6452
rect 7656 6332 7708 6384
rect 7840 6332 7892 6384
rect 8760 6332 8812 6384
rect 10968 6332 11020 6384
rect 11704 6332 11756 6384
rect 14740 6332 14792 6384
rect 7932 6264 7984 6316
rect 8944 6307 8996 6316
rect 8944 6273 8978 6307
rect 8978 6273 8996 6307
rect 8944 6264 8996 6273
rect 9312 6264 9364 6316
rect 6460 6239 6512 6248
rect 1492 6171 1544 6180
rect 1492 6137 1501 6171
rect 1501 6137 1535 6171
rect 1535 6137 1544 6171
rect 1492 6128 1544 6137
rect 2596 6128 2648 6180
rect 1676 6060 1728 6112
rect 2044 6060 2096 6112
rect 3240 6060 3292 6112
rect 4712 6128 4764 6180
rect 6460 6205 6469 6239
rect 6469 6205 6503 6239
rect 6503 6205 6512 6239
rect 6460 6196 6512 6205
rect 7196 6239 7248 6248
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 8668 6239 8720 6248
rect 8668 6205 8677 6239
rect 8677 6205 8711 6239
rect 8711 6205 8720 6239
rect 8668 6196 8720 6205
rect 11888 6196 11940 6248
rect 12164 6196 12216 6248
rect 12348 6264 12400 6316
rect 14096 6307 14148 6316
rect 14096 6273 14105 6307
rect 14105 6273 14139 6307
rect 14139 6273 14148 6307
rect 14096 6264 14148 6273
rect 12624 6196 12676 6248
rect 13084 6239 13136 6248
rect 13084 6205 13093 6239
rect 13093 6205 13127 6239
rect 13127 6205 13136 6239
rect 13084 6196 13136 6205
rect 15016 6332 15068 6384
rect 15384 6307 15436 6316
rect 15384 6273 15393 6307
rect 15393 6273 15427 6307
rect 15427 6273 15436 6307
rect 15384 6264 15436 6273
rect 5172 6060 5224 6112
rect 6368 6060 6420 6112
rect 13452 6128 13504 6180
rect 13728 6128 13780 6180
rect 8116 6060 8168 6112
rect 8944 6060 8996 6112
rect 9772 6060 9824 6112
rect 11612 6060 11664 6112
rect 12164 6103 12216 6112
rect 12164 6069 12173 6103
rect 12173 6069 12207 6103
rect 12207 6069 12216 6103
rect 12164 6060 12216 6069
rect 12992 6060 13044 6112
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 2824 5958 2876 6010
rect 2888 5958 2940 6010
rect 2952 5958 3004 6010
rect 3016 5958 3068 6010
rect 3080 5958 3132 6010
rect 6572 5958 6624 6010
rect 6636 5958 6688 6010
rect 6700 5958 6752 6010
rect 6764 5958 6816 6010
rect 6828 5958 6880 6010
rect 10320 5958 10372 6010
rect 10384 5958 10436 6010
rect 10448 5958 10500 6010
rect 10512 5958 10564 6010
rect 10576 5958 10628 6010
rect 14068 5958 14120 6010
rect 14132 5958 14184 6010
rect 14196 5958 14248 6010
rect 14260 5958 14312 6010
rect 14324 5958 14376 6010
rect 3056 5856 3108 5908
rect 3424 5899 3476 5908
rect 3424 5865 3433 5899
rect 3433 5865 3467 5899
rect 3467 5865 3476 5899
rect 3424 5856 3476 5865
rect 5816 5899 5868 5908
rect 5816 5865 5825 5899
rect 5825 5865 5859 5899
rect 5859 5865 5868 5899
rect 5816 5856 5868 5865
rect 6276 5856 6328 5908
rect 7196 5856 7248 5908
rect 1400 5788 1452 5840
rect 1952 5788 2004 5840
rect 2872 5763 2924 5772
rect 1676 5695 1728 5704
rect 1676 5661 1685 5695
rect 1685 5661 1719 5695
rect 1719 5661 1728 5695
rect 1676 5652 1728 5661
rect 2872 5729 2881 5763
rect 2881 5729 2915 5763
rect 2915 5729 2924 5763
rect 2872 5720 2924 5729
rect 4068 5720 4120 5772
rect 8300 5856 8352 5908
rect 8668 5856 8720 5908
rect 9588 5899 9640 5908
rect 9588 5865 9597 5899
rect 9597 5865 9631 5899
rect 9631 5865 9640 5899
rect 9588 5856 9640 5865
rect 7564 5831 7616 5840
rect 7564 5797 7573 5831
rect 7573 5797 7607 5831
rect 7607 5797 7616 5831
rect 7564 5788 7616 5797
rect 7748 5831 7800 5840
rect 7748 5797 7757 5831
rect 7757 5797 7791 5831
rect 7791 5797 7800 5831
rect 7748 5788 7800 5797
rect 7840 5831 7892 5840
rect 7840 5797 7849 5831
rect 7849 5797 7883 5831
rect 7883 5797 7892 5831
rect 8116 5831 8168 5840
rect 7840 5788 7892 5797
rect 8116 5797 8125 5831
rect 8125 5797 8159 5831
rect 8159 5797 8168 5831
rect 10692 5856 10744 5908
rect 11244 5899 11296 5908
rect 11244 5865 11253 5899
rect 11253 5865 11287 5899
rect 11287 5865 11296 5899
rect 11244 5856 11296 5865
rect 12716 5856 12768 5908
rect 11152 5831 11204 5840
rect 8116 5788 8168 5797
rect 11152 5797 11161 5831
rect 11161 5797 11195 5831
rect 11195 5797 11204 5831
rect 11152 5788 11204 5797
rect 12624 5788 12676 5840
rect 8392 5720 8444 5772
rect 9312 5720 9364 5772
rect 9588 5720 9640 5772
rect 2780 5652 2832 5704
rect 3056 5695 3108 5704
rect 3056 5661 3065 5695
rect 3065 5661 3099 5695
rect 3099 5661 3108 5695
rect 3056 5652 3108 5661
rect 6460 5652 6512 5704
rect 7472 5652 7524 5704
rect 7932 5652 7984 5704
rect 9864 5652 9916 5704
rect 12072 5652 12124 5704
rect 12716 5652 12768 5704
rect 13728 5856 13780 5908
rect 15384 5899 15436 5908
rect 15384 5865 15393 5899
rect 15393 5865 15427 5899
rect 15427 5865 15436 5899
rect 15384 5856 15436 5865
rect 13360 5763 13412 5772
rect 13360 5729 13369 5763
rect 13369 5729 13403 5763
rect 13403 5729 13412 5763
rect 15108 5763 15160 5772
rect 13360 5720 13412 5729
rect 15108 5729 15117 5763
rect 15117 5729 15151 5763
rect 15151 5729 15160 5763
rect 15108 5720 15160 5729
rect 14188 5652 14240 5704
rect 15568 5695 15620 5704
rect 15568 5661 15577 5695
rect 15577 5661 15611 5695
rect 15611 5661 15620 5695
rect 15568 5652 15620 5661
rect 1584 5584 1636 5636
rect 1952 5584 2004 5636
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 1860 5516 1912 5568
rect 3424 5516 3476 5568
rect 3516 5516 3568 5568
rect 3792 5516 3844 5568
rect 3884 5516 3936 5568
rect 4160 5584 4212 5636
rect 4712 5584 4764 5636
rect 9312 5584 9364 5636
rect 9772 5584 9824 5636
rect 11796 5584 11848 5636
rect 12164 5584 12216 5636
rect 4436 5516 4488 5568
rect 7104 5516 7156 5568
rect 7196 5516 7248 5568
rect 8392 5516 8444 5568
rect 8760 5559 8812 5568
rect 8760 5525 8769 5559
rect 8769 5525 8803 5559
rect 8803 5525 8812 5559
rect 8760 5516 8812 5525
rect 9128 5516 9180 5568
rect 10324 5516 10376 5568
rect 10968 5516 11020 5568
rect 11152 5516 11204 5568
rect 11704 5516 11756 5568
rect 11980 5516 12032 5568
rect 13452 5584 13504 5636
rect 14280 5584 14332 5636
rect 14648 5627 14700 5636
rect 14648 5593 14657 5627
rect 14657 5593 14691 5627
rect 14691 5593 14700 5627
rect 14648 5584 14700 5593
rect 15936 5584 15988 5636
rect 12624 5516 12676 5568
rect 12716 5516 12768 5568
rect 13268 5559 13320 5568
rect 13268 5525 13277 5559
rect 13277 5525 13311 5559
rect 13311 5525 13320 5559
rect 13268 5516 13320 5525
rect 13820 5516 13872 5568
rect 14740 5559 14792 5568
rect 14740 5525 14749 5559
rect 14749 5525 14783 5559
rect 14783 5525 14792 5559
rect 14740 5516 14792 5525
rect 15384 5516 15436 5568
rect 4698 5414 4750 5466
rect 4762 5414 4814 5466
rect 4826 5414 4878 5466
rect 4890 5414 4942 5466
rect 4954 5414 5006 5466
rect 8446 5414 8498 5466
rect 8510 5414 8562 5466
rect 8574 5414 8626 5466
rect 8638 5414 8690 5466
rect 8702 5414 8754 5466
rect 12194 5414 12246 5466
rect 12258 5414 12310 5466
rect 12322 5414 12374 5466
rect 12386 5414 12438 5466
rect 12450 5414 12502 5466
rect 2228 5355 2280 5364
rect 2228 5321 2237 5355
rect 2237 5321 2271 5355
rect 2271 5321 2280 5355
rect 2228 5312 2280 5321
rect 2320 5355 2372 5364
rect 2320 5321 2329 5355
rect 2329 5321 2363 5355
rect 2363 5321 2372 5355
rect 2320 5312 2372 5321
rect 3148 5312 3200 5364
rect 3516 5355 3568 5364
rect 3516 5321 3525 5355
rect 3525 5321 3559 5355
rect 3559 5321 3568 5355
rect 3516 5312 3568 5321
rect 5080 5355 5132 5364
rect 5080 5321 5089 5355
rect 5089 5321 5123 5355
rect 5123 5321 5132 5355
rect 5080 5312 5132 5321
rect 5448 5355 5500 5364
rect 5448 5321 5457 5355
rect 5457 5321 5491 5355
rect 5491 5321 5500 5355
rect 5448 5312 5500 5321
rect 6460 5355 6512 5364
rect 6460 5321 6469 5355
rect 6469 5321 6503 5355
rect 6503 5321 6512 5355
rect 6460 5312 6512 5321
rect 6828 5312 6880 5364
rect 8300 5355 8352 5364
rect 8300 5321 8309 5355
rect 8309 5321 8343 5355
rect 8343 5321 8352 5355
rect 8300 5312 8352 5321
rect 10048 5312 10100 5364
rect 10232 5312 10284 5364
rect 10784 5312 10836 5364
rect 12072 5312 12124 5364
rect 13728 5312 13780 5364
rect 14188 5355 14240 5364
rect 14188 5321 14197 5355
rect 14197 5321 14231 5355
rect 14231 5321 14240 5355
rect 14188 5312 14240 5321
rect 15108 5312 15160 5364
rect 5172 5244 5224 5296
rect 5540 5244 5592 5296
rect 7196 5244 7248 5296
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 2504 5219 2556 5228
rect 2504 5185 2513 5219
rect 2513 5185 2547 5219
rect 2547 5185 2556 5219
rect 2504 5176 2556 5185
rect 3884 5219 3936 5228
rect 3884 5185 3893 5219
rect 3893 5185 3927 5219
rect 3927 5185 3936 5219
rect 3884 5176 3936 5185
rect 4436 5176 4488 5228
rect 5632 5176 5684 5228
rect 5816 5219 5868 5228
rect 5816 5185 5825 5219
rect 5825 5185 5859 5219
rect 5859 5185 5868 5219
rect 5816 5176 5868 5185
rect 6920 5219 6972 5228
rect 6920 5185 6929 5219
rect 6929 5185 6963 5219
rect 6963 5185 6972 5219
rect 6920 5176 6972 5185
rect 7380 5176 7432 5228
rect 7748 5219 7800 5228
rect 1768 5151 1820 5160
rect 1768 5117 1777 5151
rect 1777 5117 1811 5151
rect 1811 5117 1820 5151
rect 1768 5108 1820 5117
rect 2872 5151 2924 5160
rect 2872 5117 2881 5151
rect 2881 5117 2915 5151
rect 2915 5117 2924 5151
rect 2872 5108 2924 5117
rect 3332 5108 3384 5160
rect 4068 5151 4120 5160
rect 4068 5117 4077 5151
rect 4077 5117 4111 5151
rect 4111 5117 4120 5151
rect 4068 5108 4120 5117
rect 5080 5108 5132 5160
rect 5724 5108 5776 5160
rect 5908 5151 5960 5160
rect 5908 5117 5917 5151
rect 5917 5117 5951 5151
rect 5951 5117 5960 5151
rect 5908 5108 5960 5117
rect 7012 5108 7064 5160
rect 7472 5108 7524 5160
rect 6184 5040 6236 5092
rect 6276 5040 6328 5092
rect 2780 4972 2832 5024
rect 4068 4972 4120 5024
rect 4620 4972 4672 5024
rect 5540 4972 5592 5024
rect 6460 4972 6512 5024
rect 6828 5040 6880 5092
rect 7748 5185 7757 5219
rect 7757 5185 7791 5219
rect 7791 5185 7800 5219
rect 7748 5176 7800 5185
rect 8208 5176 8260 5228
rect 10140 5244 10192 5296
rect 12256 5244 12308 5296
rect 15016 5244 15068 5296
rect 7656 5108 7708 5160
rect 11520 5176 11572 5228
rect 13176 5176 13228 5228
rect 14096 5219 14148 5228
rect 14096 5185 14105 5219
rect 14105 5185 14139 5219
rect 14139 5185 14148 5219
rect 14096 5176 14148 5185
rect 14924 5176 14976 5228
rect 15476 5219 15528 5228
rect 15476 5185 15485 5219
rect 15485 5185 15519 5219
rect 15519 5185 15528 5219
rect 15476 5176 15528 5185
rect 7012 4972 7064 5024
rect 7104 4972 7156 5024
rect 7840 4972 7892 5024
rect 9404 5040 9456 5092
rect 9864 4972 9916 5024
rect 10232 5040 10284 5092
rect 11244 5108 11296 5160
rect 11428 5108 11480 5160
rect 12256 5108 12308 5160
rect 12532 5151 12584 5160
rect 12532 5117 12541 5151
rect 12541 5117 12575 5151
rect 12575 5117 12584 5151
rect 12532 5108 12584 5117
rect 13452 5151 13504 5160
rect 13452 5117 13461 5151
rect 13461 5117 13495 5151
rect 13495 5117 13504 5151
rect 13452 5108 13504 5117
rect 14280 5151 14332 5160
rect 14280 5117 14289 5151
rect 14289 5117 14323 5151
rect 14323 5117 14332 5151
rect 14280 5108 14332 5117
rect 14464 5108 14516 5160
rect 14648 5040 14700 5092
rect 10692 5015 10744 5024
rect 10692 4981 10701 5015
rect 10701 4981 10735 5015
rect 10735 4981 10744 5015
rect 10692 4972 10744 4981
rect 10876 5015 10928 5024
rect 10876 4981 10885 5015
rect 10885 4981 10919 5015
rect 10919 4981 10928 5015
rect 10876 4972 10928 4981
rect 12072 5015 12124 5024
rect 12072 4981 12081 5015
rect 12081 4981 12115 5015
rect 12115 4981 12124 5015
rect 12072 4972 12124 4981
rect 12164 4972 12216 5024
rect 13636 4972 13688 5024
rect 15108 5015 15160 5024
rect 15108 4981 15117 5015
rect 15117 4981 15151 5015
rect 15151 4981 15160 5015
rect 15108 4972 15160 4981
rect 15936 4972 15988 5024
rect 2824 4870 2876 4922
rect 2888 4870 2940 4922
rect 2952 4870 3004 4922
rect 3016 4870 3068 4922
rect 3080 4870 3132 4922
rect 6572 4870 6624 4922
rect 6636 4870 6688 4922
rect 6700 4870 6752 4922
rect 6764 4870 6816 4922
rect 6828 4870 6880 4922
rect 10320 4870 10372 4922
rect 10384 4870 10436 4922
rect 10448 4870 10500 4922
rect 10512 4870 10564 4922
rect 10576 4870 10628 4922
rect 14068 4870 14120 4922
rect 14132 4870 14184 4922
rect 14196 4870 14248 4922
rect 14260 4870 14312 4922
rect 14324 4870 14376 4922
rect 1768 4768 1820 4820
rect 4160 4768 4212 4820
rect 5632 4811 5684 4820
rect 2136 4700 2188 4752
rect 3884 4700 3936 4752
rect 5632 4777 5641 4811
rect 5641 4777 5675 4811
rect 5675 4777 5684 4811
rect 5632 4768 5684 4777
rect 5908 4768 5960 4820
rect 7656 4768 7708 4820
rect 9220 4768 9272 4820
rect 10232 4768 10284 4820
rect 10416 4768 10468 4820
rect 10784 4811 10836 4820
rect 10784 4777 10793 4811
rect 10793 4777 10827 4811
rect 10827 4777 10836 4811
rect 10784 4768 10836 4777
rect 10968 4811 11020 4820
rect 10968 4777 10977 4811
rect 10977 4777 11011 4811
rect 11011 4777 11020 4811
rect 10968 4768 11020 4777
rect 11520 4811 11572 4820
rect 11520 4777 11529 4811
rect 11529 4777 11563 4811
rect 11563 4777 11572 4811
rect 11520 4768 11572 4777
rect 14832 4768 14884 4820
rect 2596 4632 2648 4684
rect 2688 4632 2740 4684
rect 3240 4632 3292 4684
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 4160 4607 4212 4616
rect 4160 4573 4169 4607
rect 4169 4573 4203 4607
rect 4203 4573 4212 4607
rect 4160 4564 4212 4573
rect 5448 4564 5500 4616
rect 5908 4632 5960 4684
rect 6368 4632 6420 4684
rect 6460 4632 6512 4684
rect 7104 4675 7156 4684
rect 6092 4607 6144 4616
rect 6092 4573 6101 4607
rect 6101 4573 6135 4607
rect 6135 4573 6144 4607
rect 7104 4641 7113 4675
rect 7113 4641 7147 4675
rect 7147 4641 7156 4675
rect 7104 4632 7156 4641
rect 7196 4632 7248 4684
rect 7748 4632 7800 4684
rect 6092 4564 6144 4573
rect 7012 4564 7064 4616
rect 9404 4700 9456 4752
rect 9588 4700 9640 4752
rect 11336 4700 11388 4752
rect 8944 4632 8996 4684
rect 9680 4675 9732 4684
rect 9680 4641 9689 4675
rect 9689 4641 9723 4675
rect 9723 4641 9732 4675
rect 9680 4632 9732 4641
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 2320 4471 2372 4480
rect 2320 4437 2329 4471
rect 2329 4437 2363 4471
rect 2363 4437 2372 4471
rect 2320 4428 2372 4437
rect 2504 4428 2556 4480
rect 2688 4428 2740 4480
rect 2780 4471 2832 4480
rect 2780 4437 2789 4471
rect 2789 4437 2823 4471
rect 2823 4437 2832 4471
rect 2780 4428 2832 4437
rect 3056 4428 3108 4480
rect 3424 4428 3476 4480
rect 3792 4428 3844 4480
rect 6184 4496 6236 4548
rect 6644 4496 6696 4548
rect 7288 4496 7340 4548
rect 8852 4496 8904 4548
rect 10232 4564 10284 4616
rect 10968 4564 11020 4616
rect 12808 4632 12860 4684
rect 13452 4700 13504 4752
rect 13636 4675 13688 4684
rect 13636 4641 13645 4675
rect 13645 4641 13679 4675
rect 13679 4641 13688 4675
rect 13636 4632 13688 4641
rect 14648 4675 14700 4684
rect 12256 4564 12308 4616
rect 14648 4641 14657 4675
rect 14657 4641 14691 4675
rect 14691 4641 14700 4675
rect 14648 4632 14700 4641
rect 14464 4607 14516 4616
rect 4804 4471 4856 4480
rect 4804 4437 4813 4471
rect 4813 4437 4847 4471
rect 4847 4437 4856 4471
rect 4804 4428 4856 4437
rect 5080 4428 5132 4480
rect 5540 4428 5592 4480
rect 6368 4428 6420 4480
rect 6460 4428 6512 4480
rect 7748 4471 7800 4480
rect 7748 4437 7757 4471
rect 7757 4437 7791 4471
rect 7791 4437 7800 4471
rect 7748 4428 7800 4437
rect 8024 4428 8076 4480
rect 8300 4428 8352 4480
rect 10324 4496 10376 4548
rect 9956 4471 10008 4480
rect 9956 4437 9965 4471
rect 9965 4437 9999 4471
rect 9999 4437 10008 4471
rect 9956 4428 10008 4437
rect 11060 4428 11112 4480
rect 11520 4428 11572 4480
rect 12164 4428 12216 4480
rect 12440 4496 12492 4548
rect 12624 4496 12676 4548
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 15108 4607 15160 4616
rect 15108 4573 15117 4607
rect 15117 4573 15151 4607
rect 15151 4573 15160 4607
rect 15108 4564 15160 4573
rect 15384 4564 15436 4616
rect 12808 4471 12860 4480
rect 12808 4437 12817 4471
rect 12817 4437 12851 4471
rect 12851 4437 12860 4471
rect 12808 4428 12860 4437
rect 13176 4471 13228 4480
rect 13176 4437 13185 4471
rect 13185 4437 13219 4471
rect 13219 4437 13228 4471
rect 13176 4428 13228 4437
rect 14464 4428 14516 4480
rect 15384 4471 15436 4480
rect 15384 4437 15393 4471
rect 15393 4437 15427 4471
rect 15427 4437 15436 4471
rect 15384 4428 15436 4437
rect 16028 4428 16080 4480
rect 4698 4326 4750 4378
rect 4762 4326 4814 4378
rect 4826 4326 4878 4378
rect 4890 4326 4942 4378
rect 4954 4326 5006 4378
rect 8446 4326 8498 4378
rect 8510 4326 8562 4378
rect 8574 4326 8626 4378
rect 8638 4326 8690 4378
rect 8702 4326 8754 4378
rect 12194 4326 12246 4378
rect 12258 4326 12310 4378
rect 12322 4326 12374 4378
rect 12386 4326 12438 4378
rect 12450 4326 12502 4378
rect 1860 4224 1912 4276
rect 2044 4267 2096 4276
rect 2044 4233 2053 4267
rect 2053 4233 2087 4267
rect 2087 4233 2096 4267
rect 2044 4224 2096 4233
rect 3148 4224 3200 4276
rect 3332 4267 3384 4276
rect 3332 4233 3341 4267
rect 3341 4233 3375 4267
rect 3375 4233 3384 4267
rect 3332 4224 3384 4233
rect 3700 4224 3752 4276
rect 5172 4267 5224 4276
rect 5172 4233 5181 4267
rect 5181 4233 5215 4267
rect 5215 4233 5224 4267
rect 5172 4224 5224 4233
rect 5540 4267 5592 4276
rect 5540 4233 5549 4267
rect 5549 4233 5583 4267
rect 5583 4233 5592 4267
rect 5540 4224 5592 4233
rect 5724 4224 5776 4276
rect 6184 4224 6236 4276
rect 7012 4224 7064 4276
rect 7748 4224 7800 4276
rect 1584 4131 1636 4140
rect 1584 4097 1593 4131
rect 1593 4097 1627 4131
rect 1627 4097 1636 4131
rect 1584 4088 1636 4097
rect 2136 4131 2188 4140
rect 2136 4097 2145 4131
rect 2145 4097 2179 4131
rect 2179 4097 2188 4131
rect 2136 4088 2188 4097
rect 2780 4088 2832 4140
rect 2596 4020 2648 4072
rect 4068 4156 4120 4208
rect 4344 4088 4396 4140
rect 4528 4131 4580 4140
rect 4528 4097 4537 4131
rect 4537 4097 4571 4131
rect 4571 4097 4580 4131
rect 4528 4088 4580 4097
rect 7380 4156 7432 4208
rect 8300 4224 8352 4276
rect 9404 4267 9456 4276
rect 9404 4233 9413 4267
rect 9413 4233 9447 4267
rect 9447 4233 9456 4267
rect 9404 4224 9456 4233
rect 10324 4267 10376 4276
rect 10324 4233 10333 4267
rect 10333 4233 10367 4267
rect 10367 4233 10376 4267
rect 10324 4224 10376 4233
rect 11060 4224 11112 4276
rect 11520 4267 11572 4276
rect 9588 4156 9640 4208
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 6000 4088 6052 4140
rect 6184 4131 6236 4140
rect 6184 4097 6193 4131
rect 6193 4097 6227 4131
rect 6227 4097 6236 4131
rect 6184 4088 6236 4097
rect 6368 4088 6420 4140
rect 6644 4088 6696 4140
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 7748 4088 7800 4140
rect 8300 4088 8352 4140
rect 8760 4131 8812 4140
rect 8760 4097 8769 4131
rect 8769 4097 8803 4131
rect 8803 4097 8812 4131
rect 8760 4088 8812 4097
rect 9220 4088 9272 4140
rect 9496 4131 9548 4140
rect 9496 4097 9505 4131
rect 9505 4097 9539 4131
rect 9539 4097 9548 4131
rect 9496 4088 9548 4097
rect 9680 4088 9732 4140
rect 9864 4088 9916 4140
rect 10232 4156 10284 4208
rect 11520 4233 11529 4267
rect 11529 4233 11563 4267
rect 11563 4233 11572 4267
rect 11520 4224 11572 4233
rect 11980 4224 12032 4276
rect 12440 4224 12492 4276
rect 12900 4224 12952 4276
rect 13820 4224 13872 4276
rect 14464 4224 14516 4276
rect 6920 4020 6972 4072
rect 7288 4063 7340 4072
rect 7288 4029 7297 4063
rect 7297 4029 7331 4063
rect 7331 4029 7340 4063
rect 7288 4020 7340 4029
rect 7932 4020 7984 4072
rect 9772 4020 9824 4072
rect 7196 3952 7248 4004
rect 9864 3995 9916 4004
rect 9864 3961 9873 3995
rect 9873 3961 9907 3995
rect 9907 3961 9916 3995
rect 9864 3952 9916 3961
rect 1400 3927 1452 3936
rect 1400 3893 1409 3927
rect 1409 3893 1443 3927
rect 1443 3893 1452 3927
rect 1400 3884 1452 3893
rect 2228 3884 2280 3936
rect 2688 3884 2740 3936
rect 3424 3927 3476 3936
rect 3424 3893 3433 3927
rect 3433 3893 3467 3927
rect 3467 3893 3476 3927
rect 3424 3884 3476 3893
rect 3700 3884 3752 3936
rect 6092 3884 6144 3936
rect 6184 3884 6236 3936
rect 7380 3927 7432 3936
rect 7380 3893 7389 3927
rect 7389 3893 7423 3927
rect 7423 3893 7432 3927
rect 7380 3884 7432 3893
rect 8208 3884 8260 3936
rect 9036 3927 9088 3936
rect 9036 3893 9045 3927
rect 9045 3893 9079 3927
rect 9079 3893 9088 3927
rect 9036 3884 9088 3893
rect 9772 3884 9824 3936
rect 10784 4063 10836 4072
rect 10784 4029 10793 4063
rect 10793 4029 10827 4063
rect 10827 4029 10836 4063
rect 10784 4020 10836 4029
rect 10508 3952 10560 4004
rect 11244 4156 11296 4208
rect 11152 4088 11204 4140
rect 11796 4156 11848 4208
rect 11520 4088 11572 4140
rect 12164 4088 12216 4140
rect 13268 4088 13320 4140
rect 14832 4088 14884 4140
rect 15660 4131 15712 4140
rect 15660 4097 15669 4131
rect 15669 4097 15703 4131
rect 15703 4097 15712 4131
rect 15660 4088 15712 4097
rect 11704 4020 11756 4072
rect 12072 4063 12124 4072
rect 12072 4029 12081 4063
rect 12081 4029 12115 4063
rect 12115 4029 12124 4063
rect 12348 4063 12400 4072
rect 12072 4020 12124 4029
rect 12348 4029 12357 4063
rect 12357 4029 12391 4063
rect 12391 4029 12400 4063
rect 12348 4020 12400 4029
rect 13176 4063 13228 4072
rect 13176 4029 13185 4063
rect 13185 4029 13219 4063
rect 13219 4029 13228 4063
rect 13176 4020 13228 4029
rect 13360 4063 13412 4072
rect 13360 4029 13369 4063
rect 13369 4029 13403 4063
rect 13403 4029 13412 4063
rect 13360 4020 13412 4029
rect 11060 3952 11112 4004
rect 12072 3884 12124 3936
rect 12808 3884 12860 3936
rect 12900 3884 12952 3936
rect 13820 3884 13872 3936
rect 14648 4020 14700 4072
rect 15752 4020 15804 4072
rect 14648 3927 14700 3936
rect 14648 3893 14657 3927
rect 14657 3893 14691 3927
rect 14691 3893 14700 3927
rect 14648 3884 14700 3893
rect 2824 3782 2876 3834
rect 2888 3782 2940 3834
rect 2952 3782 3004 3834
rect 3016 3782 3068 3834
rect 3080 3782 3132 3834
rect 6572 3782 6624 3834
rect 6636 3782 6688 3834
rect 6700 3782 6752 3834
rect 6764 3782 6816 3834
rect 6828 3782 6880 3834
rect 10320 3782 10372 3834
rect 10384 3782 10436 3834
rect 10448 3782 10500 3834
rect 10512 3782 10564 3834
rect 10576 3782 10628 3834
rect 14068 3782 14120 3834
rect 14132 3782 14184 3834
rect 14196 3782 14248 3834
rect 14260 3782 14312 3834
rect 14324 3782 14376 3834
rect 2320 3680 2372 3732
rect 2780 3680 2832 3732
rect 5172 3680 5224 3732
rect 5540 3680 5592 3732
rect 1860 3655 1912 3664
rect 1860 3621 1869 3655
rect 1869 3621 1903 3655
rect 1903 3621 1912 3655
rect 1860 3612 1912 3621
rect 3700 3612 3752 3664
rect 3240 3587 3292 3596
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 3240 3553 3249 3587
rect 3249 3553 3283 3587
rect 3283 3553 3292 3587
rect 3240 3544 3292 3553
rect 4528 3544 4580 3596
rect 1492 3408 1544 3460
rect 3424 3476 3476 3528
rect 4068 3519 4120 3528
rect 4068 3485 4077 3519
rect 4077 3485 4111 3519
rect 4111 3485 4120 3519
rect 4068 3476 4120 3485
rect 4252 3476 4304 3528
rect 4436 3408 4488 3460
rect 5816 3680 5868 3732
rect 6460 3680 6512 3732
rect 9496 3680 9548 3732
rect 9956 3680 10008 3732
rect 10784 3680 10836 3732
rect 12532 3680 12584 3732
rect 13084 3680 13136 3732
rect 6368 3612 6420 3664
rect 6644 3587 6696 3596
rect 6644 3553 6653 3587
rect 6653 3553 6687 3587
rect 6687 3553 6696 3587
rect 6644 3544 6696 3553
rect 7472 3587 7524 3596
rect 7472 3553 7481 3587
rect 7481 3553 7515 3587
rect 7515 3553 7524 3587
rect 7472 3544 7524 3553
rect 5080 3476 5132 3528
rect 5540 3519 5592 3528
rect 5540 3485 5549 3519
rect 5549 3485 5583 3519
rect 5583 3485 5592 3519
rect 5540 3476 5592 3485
rect 7104 3476 7156 3528
rect 7288 3476 7340 3528
rect 7748 3519 7800 3528
rect 7748 3485 7757 3519
rect 7757 3485 7791 3519
rect 7791 3485 7800 3519
rect 7748 3476 7800 3485
rect 9036 3612 9088 3664
rect 8944 3544 8996 3596
rect 9680 3544 9732 3596
rect 10600 3544 10652 3596
rect 9312 3476 9364 3528
rect 8760 3451 8812 3460
rect 8760 3417 8769 3451
rect 8769 3417 8803 3451
rect 8803 3417 8812 3451
rect 8760 3408 8812 3417
rect 9588 3408 9640 3460
rect 10140 3476 10192 3528
rect 10968 3476 11020 3528
rect 11244 3544 11296 3596
rect 11980 3587 12032 3596
rect 11980 3553 11989 3587
rect 11989 3553 12023 3587
rect 12023 3553 12032 3587
rect 11980 3544 12032 3553
rect 12624 3544 12676 3596
rect 13176 3544 13228 3596
rect 13360 3680 13412 3732
rect 15108 3680 15160 3732
rect 13728 3612 13780 3664
rect 14924 3612 14976 3664
rect 14832 3587 14884 3596
rect 14832 3553 14841 3587
rect 14841 3553 14875 3587
rect 14875 3553 14884 3587
rect 14832 3544 14884 3553
rect 15568 3544 15620 3596
rect 1584 3383 1636 3392
rect 1584 3349 1593 3383
rect 1593 3349 1627 3383
rect 1627 3349 1636 3383
rect 1584 3340 1636 3349
rect 1860 3340 1912 3392
rect 2228 3383 2280 3392
rect 2228 3349 2237 3383
rect 2237 3349 2271 3383
rect 2271 3349 2280 3383
rect 2228 3340 2280 3349
rect 3148 3383 3200 3392
rect 3148 3349 3157 3383
rect 3157 3349 3191 3383
rect 3191 3349 3200 3383
rect 3148 3340 3200 3349
rect 3884 3383 3936 3392
rect 3884 3349 3893 3383
rect 3893 3349 3927 3383
rect 3927 3349 3936 3383
rect 3884 3340 3936 3349
rect 5172 3340 5224 3392
rect 5540 3340 5592 3392
rect 6276 3340 6328 3392
rect 7012 3340 7064 3392
rect 7564 3340 7616 3392
rect 7932 3340 7984 3392
rect 8944 3340 8996 3392
rect 9312 3383 9364 3392
rect 9312 3349 9321 3383
rect 9321 3349 9355 3383
rect 9355 3349 9364 3383
rect 9312 3340 9364 3349
rect 9404 3383 9456 3392
rect 9404 3349 9413 3383
rect 9413 3349 9447 3383
rect 9447 3349 9456 3383
rect 10048 3383 10100 3392
rect 9404 3340 9456 3349
rect 10048 3349 10057 3383
rect 10057 3349 10091 3383
rect 10091 3349 10100 3383
rect 10048 3340 10100 3349
rect 12900 3476 12952 3528
rect 13728 3476 13780 3528
rect 14740 3476 14792 3528
rect 15016 3476 15068 3528
rect 11152 3408 11204 3460
rect 11244 3408 11296 3460
rect 12440 3408 12492 3460
rect 13912 3408 13964 3460
rect 10968 3383 11020 3392
rect 10968 3349 10977 3383
rect 10977 3349 11011 3383
rect 11011 3349 11020 3383
rect 10968 3340 11020 3349
rect 12624 3383 12676 3392
rect 12624 3349 12633 3383
rect 12633 3349 12667 3383
rect 12667 3349 12676 3383
rect 12624 3340 12676 3349
rect 13176 3340 13228 3392
rect 13636 3340 13688 3392
rect 14464 3340 14516 3392
rect 15016 3340 15068 3392
rect 4698 3238 4750 3290
rect 4762 3238 4814 3290
rect 4826 3238 4878 3290
rect 4890 3238 4942 3290
rect 4954 3238 5006 3290
rect 8446 3238 8498 3290
rect 8510 3238 8562 3290
rect 8574 3238 8626 3290
rect 8638 3238 8690 3290
rect 8702 3238 8754 3290
rect 12194 3238 12246 3290
rect 12258 3238 12310 3290
rect 12322 3238 12374 3290
rect 12386 3238 12438 3290
rect 12450 3238 12502 3290
rect 2688 3068 2740 3120
rect 3148 3136 3200 3188
rect 4528 3136 4580 3188
rect 2044 3000 2096 3052
rect 2412 3000 2464 3052
rect 2780 3043 2832 3052
rect 2780 3009 2789 3043
rect 2789 3009 2823 3043
rect 2823 3009 2832 3043
rect 2780 3000 2832 3009
rect 3976 3068 4028 3120
rect 5172 3136 5224 3188
rect 5448 3136 5500 3188
rect 6092 3136 6144 3188
rect 6276 3136 6328 3188
rect 3884 3000 3936 3052
rect 4620 3000 4672 3052
rect 5264 3000 5316 3052
rect 4344 2975 4396 2984
rect 4344 2941 4353 2975
rect 4353 2941 4387 2975
rect 4387 2941 4396 2975
rect 4344 2932 4396 2941
rect 5172 2932 5224 2984
rect 5632 3000 5684 3052
rect 5908 2932 5960 2984
rect 2688 2864 2740 2916
rect 3148 2864 3200 2916
rect 6828 3136 6880 3188
rect 7104 3136 7156 3188
rect 7656 3136 7708 3188
rect 8944 3179 8996 3188
rect 8944 3145 8953 3179
rect 8953 3145 8987 3179
rect 8987 3145 8996 3179
rect 8944 3136 8996 3145
rect 9312 3136 9364 3188
rect 7840 3068 7892 3120
rect 10048 3136 10100 3188
rect 7196 3043 7248 3052
rect 7196 3009 7205 3043
rect 7205 3009 7239 3043
rect 7239 3009 7248 3043
rect 7196 3000 7248 3009
rect 7748 3000 7800 3052
rect 8116 3043 8168 3052
rect 8116 3009 8125 3043
rect 8125 3009 8159 3043
rect 8159 3009 8168 3043
rect 8116 3000 8168 3009
rect 8208 3000 8260 3052
rect 7472 2932 7524 2984
rect 7840 2975 7892 2984
rect 7840 2941 7849 2975
rect 7849 2941 7883 2975
rect 7883 2941 7892 2975
rect 7840 2932 7892 2941
rect 10232 3068 10284 3120
rect 9312 3000 9364 3052
rect 9588 3000 9640 3052
rect 9864 3043 9916 3052
rect 9864 3009 9873 3043
rect 9873 3009 9907 3043
rect 9907 3009 9916 3043
rect 9864 3000 9916 3009
rect 9680 2932 9732 2984
rect 9956 2975 10008 2984
rect 9956 2941 9965 2975
rect 9965 2941 9999 2975
rect 9999 2941 10008 2975
rect 9956 2932 10008 2941
rect 6920 2864 6972 2916
rect 7196 2864 7248 2916
rect 8392 2864 8444 2916
rect 9404 2864 9456 2916
rect 1216 2796 1268 2848
rect 2044 2839 2096 2848
rect 2044 2805 2053 2839
rect 2053 2805 2087 2839
rect 2087 2805 2096 2839
rect 2044 2796 2096 2805
rect 2596 2839 2648 2848
rect 2596 2805 2605 2839
rect 2605 2805 2639 2839
rect 2639 2805 2648 2839
rect 3240 2839 3292 2848
rect 2596 2796 2648 2805
rect 3240 2805 3249 2839
rect 3249 2805 3283 2839
rect 3283 2805 3292 2839
rect 3240 2796 3292 2805
rect 4712 2796 4764 2848
rect 5172 2839 5224 2848
rect 5172 2805 5181 2839
rect 5181 2805 5215 2839
rect 5215 2805 5224 2839
rect 5172 2796 5224 2805
rect 5724 2796 5776 2848
rect 7012 2796 7064 2848
rect 7104 2796 7156 2848
rect 8484 2839 8536 2848
rect 8484 2805 8493 2839
rect 8493 2805 8527 2839
rect 8527 2805 8536 2839
rect 8484 2796 8536 2805
rect 10600 2864 10652 2916
rect 11336 3136 11388 3188
rect 12072 3136 12124 3188
rect 12624 3136 12676 3188
rect 12808 3179 12860 3188
rect 12808 3145 12817 3179
rect 12817 3145 12851 3179
rect 12851 3145 12860 3179
rect 12808 3136 12860 3145
rect 10876 3068 10928 3120
rect 11428 3068 11480 3120
rect 12716 3111 12768 3120
rect 12716 3077 12725 3111
rect 12725 3077 12759 3111
rect 12759 3077 12768 3111
rect 12716 3068 12768 3077
rect 11980 2932 12032 2984
rect 13820 3000 13872 3052
rect 14096 3043 14148 3052
rect 14096 3009 14105 3043
rect 14105 3009 14139 3043
rect 14139 3009 14148 3043
rect 14096 3000 14148 3009
rect 14556 3043 14608 3052
rect 13268 2932 13320 2984
rect 13636 2932 13688 2984
rect 14556 3009 14565 3043
rect 14565 3009 14599 3043
rect 14599 3009 14608 3043
rect 14556 3000 14608 3009
rect 15844 3000 15896 3052
rect 14372 2932 14424 2984
rect 13820 2864 13872 2916
rect 11612 2796 11664 2848
rect 11796 2796 11848 2848
rect 12072 2796 12124 2848
rect 13176 2796 13228 2848
rect 13452 2796 13504 2848
rect 15384 2796 15436 2848
rect 2824 2694 2876 2746
rect 2888 2694 2940 2746
rect 2952 2694 3004 2746
rect 3016 2694 3068 2746
rect 3080 2694 3132 2746
rect 6572 2694 6624 2746
rect 6636 2694 6688 2746
rect 6700 2694 6752 2746
rect 6764 2694 6816 2746
rect 6828 2694 6880 2746
rect 10320 2694 10372 2746
rect 10384 2694 10436 2746
rect 10448 2694 10500 2746
rect 10512 2694 10564 2746
rect 10576 2694 10628 2746
rect 14068 2694 14120 2746
rect 14132 2694 14184 2746
rect 14196 2694 14248 2746
rect 14260 2694 14312 2746
rect 14324 2694 14376 2746
rect 8208 2592 8260 2644
rect 9036 2635 9088 2644
rect 9036 2601 9045 2635
rect 9045 2601 9079 2635
rect 9079 2601 9088 2635
rect 9036 2592 9088 2601
rect 9772 2592 9824 2644
rect 10968 2592 11020 2644
rect 15016 2592 15068 2644
rect 2044 2456 2096 2508
rect 1860 2431 1912 2440
rect 1860 2397 1869 2431
rect 1869 2397 1903 2431
rect 1903 2397 1912 2431
rect 2228 2431 2280 2440
rect 1860 2388 1912 2397
rect 2228 2397 2237 2431
rect 2237 2397 2271 2431
rect 2271 2397 2280 2431
rect 2228 2388 2280 2397
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 2780 2388 2832 2440
rect 3148 2388 3200 2440
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 7840 2524 7892 2576
rect 8024 2567 8076 2576
rect 8024 2533 8033 2567
rect 8033 2533 8067 2567
rect 8067 2533 8076 2567
rect 8024 2524 8076 2533
rect 9496 2524 9548 2576
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 6000 2456 6052 2508
rect 6092 2456 6144 2508
rect 5172 2431 5224 2440
rect 5172 2397 5181 2431
rect 5181 2397 5215 2431
rect 5215 2397 5224 2431
rect 5816 2431 5868 2440
rect 5172 2388 5224 2397
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 6184 2431 6236 2440
rect 6184 2397 6193 2431
rect 6193 2397 6227 2431
rect 6227 2397 6236 2431
rect 6184 2388 6236 2397
rect 8300 2456 8352 2508
rect 8484 2499 8536 2508
rect 8484 2465 8493 2499
rect 8493 2465 8527 2499
rect 8527 2465 8536 2499
rect 8484 2456 8536 2465
rect 9588 2456 9640 2508
rect 9864 2499 9916 2508
rect 9864 2465 9873 2499
rect 9873 2465 9907 2499
rect 9907 2465 9916 2499
rect 9864 2456 9916 2465
rect 10324 2456 10376 2508
rect 7380 2388 7432 2440
rect 7932 2431 7984 2440
rect 7932 2397 7941 2431
rect 7941 2397 7975 2431
rect 7975 2397 7984 2431
rect 7932 2388 7984 2397
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 3608 2320 3660 2372
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 1952 2252 2004 2304
rect 2320 2252 2372 2304
rect 2688 2252 2740 2304
rect 3424 2252 3476 2304
rect 3792 2252 3844 2304
rect 4160 2252 4212 2304
rect 4528 2295 4580 2304
rect 4528 2261 4537 2295
rect 4537 2261 4571 2295
rect 4571 2261 4580 2295
rect 4528 2252 4580 2261
rect 5080 2252 5132 2304
rect 5264 2252 5316 2304
rect 5908 2252 5960 2304
rect 6276 2252 6328 2304
rect 6460 2295 6512 2304
rect 6460 2261 6469 2295
rect 6469 2261 6503 2295
rect 6503 2261 6512 2295
rect 6460 2252 6512 2261
rect 6736 2295 6788 2304
rect 6736 2261 6745 2295
rect 6745 2261 6779 2295
rect 6779 2261 6788 2295
rect 6736 2252 6788 2261
rect 7472 2252 7524 2304
rect 8944 2252 8996 2304
rect 9680 2320 9732 2372
rect 10232 2252 10284 2304
rect 10416 2320 10468 2372
rect 10692 2388 10744 2440
rect 10600 2320 10652 2372
rect 11428 2388 11480 2440
rect 11704 2431 11756 2440
rect 11704 2397 11713 2431
rect 11713 2397 11747 2431
rect 11747 2397 11756 2431
rect 11704 2388 11756 2397
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 12624 2388 12676 2440
rect 12900 2431 12952 2440
rect 12900 2397 12909 2431
rect 12909 2397 12943 2431
rect 12943 2397 12952 2431
rect 12900 2388 12952 2397
rect 11244 2320 11296 2372
rect 13544 2388 13596 2440
rect 14372 2431 14424 2440
rect 14372 2397 14381 2431
rect 14381 2397 14415 2431
rect 14415 2397 14424 2431
rect 14372 2388 14424 2397
rect 15200 2456 15252 2508
rect 15476 2456 15528 2508
rect 13084 2320 13136 2372
rect 4698 2150 4750 2202
rect 4762 2150 4814 2202
rect 4826 2150 4878 2202
rect 4890 2150 4942 2202
rect 4954 2150 5006 2202
rect 8446 2150 8498 2202
rect 8510 2150 8562 2202
rect 8574 2150 8626 2202
rect 8638 2150 8690 2202
rect 8702 2150 8754 2202
rect 12194 2150 12246 2202
rect 12258 2150 12310 2202
rect 12322 2150 12374 2202
rect 12386 2150 12438 2202
rect 12450 2150 12502 2202
rect 6460 2048 6512 2100
rect 5816 1980 5868 2032
rect 7932 2048 7984 2100
rect 15384 2048 15436 2100
rect 9680 1980 9732 2032
rect 9864 1980 9916 2032
rect 11612 1980 11664 2032
rect 11060 1912 11112 1964
rect 10048 1504 10100 1556
rect 11704 1504 11756 1556
<< metal2 >>
rect 1030 19200 1086 20000
rect 1398 19200 1454 20000
rect 1766 19200 1822 20000
rect 2134 19200 2190 20000
rect 2502 19200 2558 20000
rect 2870 19200 2926 20000
rect 3238 19200 3294 20000
rect 3606 19200 3662 20000
rect 3974 19200 4030 20000
rect 4342 19200 4398 20000
rect 4710 19200 4766 20000
rect 5078 19200 5134 20000
rect 5446 19200 5502 20000
rect 5814 19200 5870 20000
rect 6182 19200 6238 20000
rect 6550 19200 6606 20000
rect 6918 19200 6974 20000
rect 7286 19200 7342 20000
rect 7654 19200 7710 20000
rect 8022 19200 8078 20000
rect 8390 19200 8446 20000
rect 8758 19200 8814 20000
rect 9126 19200 9182 20000
rect 9494 19200 9550 20000
rect 9862 19200 9918 20000
rect 10230 19200 10286 20000
rect 10598 19200 10654 20000
rect 10966 19200 11022 20000
rect 11334 19200 11390 20000
rect 11702 19200 11758 20000
rect 12070 19200 12126 20000
rect 12438 19200 12494 20000
rect 12806 19200 12862 20000
rect 13174 19200 13230 20000
rect 13542 19200 13598 20000
rect 13910 19200 13966 20000
rect 14278 19200 14334 20000
rect 14384 19230 14596 19258
rect 1044 17066 1072 19200
rect 1306 18592 1362 18601
rect 1306 18527 1362 18536
rect 1032 17060 1084 17066
rect 1032 17002 1084 17008
rect 1044 14074 1072 17002
rect 1320 15858 1348 18527
rect 1412 16454 1440 19200
rect 1780 17338 1808 19200
rect 2148 17338 2176 19200
rect 2318 17640 2374 17649
rect 2318 17575 2374 17584
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 2136 17332 2188 17338
rect 2136 17274 2188 17280
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1780 16794 1808 17138
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 2332 16726 2360 17575
rect 2516 17338 2544 19200
rect 2778 19136 2834 19145
rect 2778 19071 2834 19080
rect 2504 17332 2556 17338
rect 2504 17274 2556 17280
rect 2412 17196 2464 17202
rect 2412 17138 2464 17144
rect 1952 16720 2004 16726
rect 1950 16688 1952 16697
rect 2320 16720 2372 16726
rect 2004 16688 2006 16697
rect 2320 16662 2372 16668
rect 1950 16623 2006 16632
rect 2136 16584 2188 16590
rect 2136 16526 2188 16532
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 1400 16448 1452 16454
rect 1400 16390 1452 16396
rect 2148 16250 2176 16526
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 1492 15904 1544 15910
rect 1320 15830 1440 15858
rect 1492 15846 1544 15852
rect 1412 15706 1440 15830
rect 1504 15745 1532 15846
rect 1490 15736 1546 15745
rect 1400 15700 1452 15706
rect 2240 15706 2268 16526
rect 2318 16144 2374 16153
rect 2318 16079 2320 16088
rect 2372 16079 2374 16088
rect 2320 16050 2372 16056
rect 2424 15706 2452 17138
rect 2792 17082 2820 19071
rect 2884 17338 2912 19200
rect 3252 17338 3280 19200
rect 3620 17338 3648 19200
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 3240 17332 3292 17338
rect 3240 17274 3292 17280
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 2700 17054 2820 17082
rect 3148 17128 3200 17134
rect 3148 17070 3200 17076
rect 2700 16674 2728 17054
rect 2824 16892 3132 16901
rect 2824 16890 2830 16892
rect 2886 16890 2910 16892
rect 2966 16890 2990 16892
rect 3046 16890 3070 16892
rect 3126 16890 3132 16892
rect 2886 16838 2888 16890
rect 3068 16838 3070 16890
rect 2824 16836 2830 16838
rect 2886 16836 2910 16838
rect 2966 16836 2990 16838
rect 3046 16836 3070 16838
rect 3126 16836 3132 16838
rect 2824 16827 3132 16836
rect 3160 16794 3188 17070
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 3252 16726 3280 17138
rect 3344 16794 3372 17138
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 3240 16720 3292 16726
rect 2504 16652 2556 16658
rect 2700 16646 2820 16674
rect 3240 16662 3292 16668
rect 2504 16594 2556 16600
rect 1490 15671 1546 15680
rect 2228 15700 2280 15706
rect 1400 15642 1452 15648
rect 2228 15642 2280 15648
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2136 15632 2188 15638
rect 2136 15574 2188 15580
rect 2042 15464 2098 15473
rect 2042 15399 2098 15408
rect 2056 15366 2084 15399
rect 2148 15366 2176 15574
rect 2044 15360 2096 15366
rect 2136 15360 2188 15366
rect 2044 15302 2096 15308
rect 2134 15328 2136 15337
rect 2412 15360 2464 15366
rect 2188 15328 2190 15337
rect 2134 15263 2190 15272
rect 2410 15328 2412 15337
rect 2464 15328 2466 15337
rect 2410 15263 2466 15272
rect 1950 15056 2006 15065
rect 1584 15020 1636 15026
rect 1950 14991 1952 15000
rect 1584 14962 1636 14968
rect 2004 14991 2006 15000
rect 1952 14962 2004 14968
rect 1492 14816 1544 14822
rect 1490 14784 1492 14793
rect 1544 14784 1546 14793
rect 1490 14719 1546 14728
rect 1596 14618 1624 14962
rect 2412 14884 2464 14890
rect 2412 14826 2464 14832
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1032 14068 1084 14074
rect 1032 14010 1084 14016
rect 1688 13938 1716 14758
rect 1950 13968 2006 13977
rect 1676 13932 1728 13938
rect 1950 13903 2006 13912
rect 1676 13874 1728 13880
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1490 13832 1546 13841
rect 1412 6798 1440 13806
rect 1490 13767 1492 13776
rect 1544 13767 1546 13776
rect 1492 13738 1544 13744
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 1504 12889 1532 13126
rect 1490 12880 1546 12889
rect 1490 12815 1546 12824
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1490 11928 1546 11937
rect 1490 11863 1492 11872
rect 1544 11863 1546 11872
rect 1492 11834 1544 11840
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1492 11008 1544 11014
rect 1490 10976 1492 10985
rect 1544 10976 1546 10985
rect 1490 10911 1546 10920
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 10062 1716 10406
rect 1780 10266 1808 11086
rect 1872 10810 1900 12038
rect 1860 10804 1912 10810
rect 1860 10746 1912 10752
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1676 10056 1728 10062
rect 1490 10024 1546 10033
rect 1676 9998 1728 10004
rect 1964 10010 1992 13903
rect 2228 13864 2280 13870
rect 2228 13806 2280 13812
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 2056 11354 2084 12038
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2148 10810 2176 11494
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 1964 9982 2084 10010
rect 1490 9959 1546 9968
rect 1504 9926 1532 9959
rect 1492 9920 1544 9926
rect 1492 9862 1544 9868
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 1582 9616 1638 9625
rect 1964 9586 1992 9862
rect 1582 9551 1638 9560
rect 1676 9580 1728 9586
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1504 9081 1532 9318
rect 1490 9072 1546 9081
rect 1490 9007 1546 9016
rect 1490 8120 1546 8129
rect 1490 8055 1492 8064
rect 1544 8055 1546 8064
rect 1492 8026 1544 8032
rect 1492 7200 1544 7206
rect 1490 7168 1492 7177
rect 1544 7168 1546 7177
rect 1490 7103 1546 7112
rect 1596 6866 1624 9551
rect 1676 9522 1728 9528
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 1688 7546 1716 9522
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1490 6216 1546 6225
rect 1490 6151 1492 6160
rect 1544 6151 1546 6160
rect 1492 6122 1544 6128
rect 1400 5840 1452 5846
rect 1400 5782 1452 5788
rect 1412 4026 1440 5782
rect 1596 5642 1624 6802
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1688 5710 1716 6054
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1584 5636 1636 5642
rect 1584 5578 1636 5584
rect 1492 5568 1544 5574
rect 1780 5522 1808 9318
rect 1872 8430 1900 9386
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 2056 7546 2084 9982
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2056 7002 2084 7482
rect 2240 7426 2268 13806
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2332 13326 2360 13670
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2332 12986 2360 13126
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2332 11762 2360 12038
rect 2424 11830 2452 14826
rect 2516 14822 2544 16594
rect 2688 16516 2740 16522
rect 2688 16458 2740 16464
rect 2700 16425 2728 16458
rect 2686 16416 2742 16425
rect 2686 16351 2742 16360
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 2688 16108 2740 16114
rect 2688 16050 2740 16056
rect 2608 15638 2636 16050
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 2700 15586 2728 16050
rect 2792 15978 2820 16646
rect 3240 16584 3292 16590
rect 3240 16526 3292 16532
rect 3608 16584 3660 16590
rect 3608 16526 3660 16532
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3146 16416 3202 16425
rect 3146 16351 3202 16360
rect 2780 15972 2832 15978
rect 2780 15914 2832 15920
rect 2824 15804 3132 15813
rect 2824 15802 2830 15804
rect 2886 15802 2910 15804
rect 2966 15802 2990 15804
rect 3046 15802 3070 15804
rect 3126 15802 3132 15804
rect 2886 15750 2888 15802
rect 3068 15750 3070 15802
rect 2824 15748 2830 15750
rect 2886 15748 2910 15750
rect 2966 15748 2990 15750
rect 3046 15748 3070 15750
rect 3126 15748 3132 15750
rect 2824 15739 3132 15748
rect 2700 15570 2820 15586
rect 2700 15564 2832 15570
rect 2700 15558 2780 15564
rect 2780 15506 2832 15512
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 2792 15178 2820 15302
rect 2700 15150 2820 15178
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2516 12850 2544 14758
rect 2700 14600 2728 15150
rect 3068 14929 3096 15302
rect 3160 15094 3188 16351
rect 3148 15088 3200 15094
rect 3148 15030 3200 15036
rect 3054 14920 3110 14929
rect 3252 14890 3280 16526
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 3436 15706 3464 15982
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 3422 15600 3478 15609
rect 3332 15564 3384 15570
rect 3422 15535 3478 15544
rect 3332 15506 3384 15512
rect 3054 14855 3110 14864
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 2824 14716 3132 14725
rect 2824 14714 2830 14716
rect 2886 14714 2910 14716
rect 2966 14714 2990 14716
rect 3046 14714 3070 14716
rect 3126 14714 3132 14716
rect 2886 14662 2888 14714
rect 3068 14662 3070 14714
rect 2824 14660 2830 14662
rect 2886 14660 2910 14662
rect 2966 14660 2990 14662
rect 3046 14660 3070 14662
rect 3126 14660 3132 14662
rect 2824 14651 3132 14660
rect 2700 14572 2820 14600
rect 2596 14544 2648 14550
rect 2596 14486 2648 14492
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2608 11898 2636 14486
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2700 13297 2728 14350
rect 2792 14006 2820 14572
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 2780 14000 2832 14006
rect 2780 13942 2832 13948
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 2884 13870 2912 13942
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 3068 13716 3096 14418
rect 3160 14414 3188 14758
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 3068 13688 3188 13716
rect 2824 13628 3132 13637
rect 2824 13626 2830 13628
rect 2886 13626 2910 13628
rect 2966 13626 2990 13628
rect 3046 13626 3070 13628
rect 3126 13626 3132 13628
rect 2886 13574 2888 13626
rect 3068 13574 3070 13626
rect 2824 13572 2830 13574
rect 2886 13572 2910 13574
rect 2966 13572 2990 13574
rect 3046 13572 3070 13574
rect 3126 13572 3132 13574
rect 2824 13563 3132 13572
rect 3160 13530 3188 13688
rect 3148 13524 3200 13530
rect 3148 13466 3200 13472
rect 3160 13394 3188 13466
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 2686 13288 2742 13297
rect 2686 13223 2742 13232
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 2824 12540 3132 12549
rect 2824 12538 2830 12540
rect 2886 12538 2910 12540
rect 2966 12538 2990 12540
rect 3046 12538 3070 12540
rect 3126 12538 3132 12540
rect 2886 12486 2888 12538
rect 3068 12486 3070 12538
rect 2824 12484 2830 12486
rect 2886 12484 2910 12486
rect 2966 12484 2990 12486
rect 3046 12484 3070 12486
rect 3126 12484 3132 12486
rect 2824 12475 3132 12484
rect 3160 12442 3188 12786
rect 3238 12608 3294 12617
rect 3238 12543 3294 12552
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3252 12102 3280 12543
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2412 11824 2464 11830
rect 2412 11766 2464 11772
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2424 10198 2452 11766
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2516 11218 2544 11494
rect 2608 11234 2636 11834
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 2824 11452 3132 11461
rect 2824 11450 2830 11452
rect 2886 11450 2910 11452
rect 2966 11450 2990 11452
rect 3046 11450 3070 11452
rect 3126 11450 3132 11452
rect 2886 11398 2888 11450
rect 3068 11398 3070 11450
rect 2824 11396 2830 11398
rect 2886 11396 2910 11398
rect 2966 11396 2990 11398
rect 3046 11396 3070 11398
rect 3126 11396 3132 11398
rect 2824 11387 3132 11396
rect 3160 11234 3188 11698
rect 3252 11558 3280 12038
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 3252 11393 3280 11494
rect 3238 11384 3294 11393
rect 3238 11319 3294 11328
rect 2504 11212 2556 11218
rect 2608 11206 2728 11234
rect 3160 11206 3280 11234
rect 2504 11154 2556 11160
rect 2596 11144 2648 11150
rect 2596 11086 2648 11092
rect 2608 10606 2636 11086
rect 2596 10600 2648 10606
rect 2596 10542 2648 10548
rect 2412 10192 2464 10198
rect 2412 10134 2464 10140
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 2332 8634 2360 9862
rect 2516 9722 2544 9862
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2424 9178 2452 9522
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2516 8634 2544 9454
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2608 8514 2636 9114
rect 2700 8974 2728 11206
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10606 3188 10950
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 2824 10364 3132 10373
rect 2824 10362 2830 10364
rect 2886 10362 2910 10364
rect 2966 10362 2990 10364
rect 3046 10362 3070 10364
rect 3126 10362 3132 10364
rect 2886 10310 2888 10362
rect 3068 10310 3070 10362
rect 2824 10308 2830 10310
rect 2886 10308 2910 10310
rect 2966 10308 2990 10310
rect 3046 10308 3070 10310
rect 3126 10308 3132 10310
rect 2824 10299 3132 10308
rect 2824 9276 3132 9285
rect 2824 9274 2830 9276
rect 2886 9274 2910 9276
rect 2966 9274 2990 9276
rect 3046 9274 3070 9276
rect 3126 9274 3132 9276
rect 2886 9222 2888 9274
rect 3068 9222 3070 9274
rect 2824 9220 2830 9222
rect 2886 9220 2910 9222
rect 2966 9220 2990 9222
rect 3046 9220 3070 9222
rect 3126 9220 3132 9222
rect 2824 9211 3132 9220
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 3160 8906 3188 10542
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 2884 8634 2912 8842
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3252 8566 3280 11206
rect 3344 11014 3372 15506
rect 3436 15366 3464 15535
rect 3424 15360 3476 15366
rect 3424 15302 3476 15308
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 3436 14958 3464 15098
rect 3424 14952 3476 14958
rect 3528 14929 3556 16050
rect 3620 15337 3648 16526
rect 3700 16448 3752 16454
rect 3700 16390 3752 16396
rect 3606 15328 3662 15337
rect 3606 15263 3662 15272
rect 3712 15026 3740 16390
rect 3896 15570 3924 16526
rect 3988 16454 4016 19200
rect 4068 17808 4120 17814
rect 4068 17750 4120 17756
rect 4080 17338 4108 17750
rect 4356 17338 4384 19200
rect 4724 17524 4752 19200
rect 4632 17496 4752 17524
rect 4632 17338 4660 17496
rect 4698 17436 5006 17445
rect 4698 17434 4704 17436
rect 4760 17434 4784 17436
rect 4840 17434 4864 17436
rect 4920 17434 4944 17436
rect 5000 17434 5006 17436
rect 4760 17382 4762 17434
rect 4942 17382 4944 17434
rect 4698 17380 4704 17382
rect 4760 17380 4784 17382
rect 4840 17380 4864 17382
rect 4920 17380 4944 17382
rect 5000 17380 5006 17382
rect 4698 17371 5006 17380
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4436 17264 4488 17270
rect 4436 17206 4488 17212
rect 4710 17232 4766 17241
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 3976 16448 4028 16454
rect 3976 16390 4028 16396
rect 4080 16250 4108 16526
rect 4160 16516 4212 16522
rect 4160 16458 4212 16464
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 3976 16176 4028 16182
rect 3976 16118 4028 16124
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3882 15328 3938 15337
rect 3804 15162 3832 15302
rect 3882 15263 3938 15272
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 3700 15020 3752 15026
rect 3700 14962 3752 14968
rect 3608 14952 3660 14958
rect 3424 14894 3476 14900
rect 3514 14920 3570 14929
rect 3608 14894 3660 14900
rect 3514 14855 3570 14864
rect 3620 14822 3648 14894
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3422 14104 3478 14113
rect 3422 14039 3478 14048
rect 3436 14006 3464 14039
rect 3424 14000 3476 14006
rect 3424 13942 3476 13948
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 3436 12986 3464 13330
rect 3528 13326 3556 14214
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3332 11008 3384 11014
rect 3332 10950 3384 10956
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3344 8838 3372 9522
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 2148 7398 2268 7426
rect 2516 8486 2636 8514
rect 3148 8560 3200 8566
rect 3148 8502 3200 8508
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 2412 7404 2464 7410
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 1872 5574 1900 6734
rect 1964 5846 1992 6802
rect 2056 6202 2084 6938
rect 2148 6866 2176 7398
rect 2412 7346 2464 7352
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 2318 7304 2374 7313
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2136 6656 2188 6662
rect 2134 6624 2136 6633
rect 2188 6624 2190 6633
rect 2134 6559 2190 6568
rect 2240 6474 2268 7278
rect 2318 7239 2320 7248
rect 2372 7239 2374 7248
rect 2320 7210 2372 7216
rect 2240 6446 2360 6474
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2056 6174 2176 6202
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 1952 5840 2004 5846
rect 1952 5782 2004 5788
rect 1952 5636 2004 5642
rect 1952 5578 2004 5584
rect 1492 5510 1544 5516
rect 1504 5273 1532 5510
rect 1688 5494 1808 5522
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1490 5264 1546 5273
rect 1490 5199 1546 5208
rect 1688 4622 1716 5494
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 1780 4826 1808 5102
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1492 4480 1544 4486
rect 1492 4422 1544 4428
rect 1504 4321 1532 4422
rect 1490 4312 1546 4321
rect 1872 4282 1900 5170
rect 1490 4247 1546 4256
rect 1860 4276 1912 4282
rect 1860 4218 1912 4224
rect 1584 4140 1636 4146
rect 1584 4082 1636 4088
rect 1596 4049 1624 4082
rect 1582 4040 1638 4049
rect 1412 3998 1532 4026
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 1412 3534 1440 3878
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 1504 3466 1532 3998
rect 1582 3975 1638 3984
rect 1860 3664 1912 3670
rect 1858 3632 1860 3641
rect 1912 3632 1914 3641
rect 1858 3567 1914 3576
rect 1492 3460 1544 3466
rect 1492 3402 1544 3408
rect 1584 3392 1636 3398
rect 1582 3360 1584 3369
rect 1860 3392 1912 3398
rect 1636 3360 1638 3369
rect 1860 3334 1912 3340
rect 1582 3295 1638 3304
rect 1216 2848 1268 2854
rect 1216 2790 1268 2796
rect 1228 800 1256 2790
rect 1872 2446 1900 3334
rect 1964 3040 1992 5578
rect 2056 4282 2084 6054
rect 2148 4842 2176 6174
rect 2240 5370 2268 6258
rect 2332 5370 2360 6446
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2148 4814 2268 4842
rect 2136 4752 2188 4758
rect 2136 4694 2188 4700
rect 2044 4276 2096 4282
rect 2044 4218 2096 4224
rect 2148 4146 2176 4694
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2240 3942 2268 4814
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2332 3738 2360 4422
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2228 3392 2280 3398
rect 2228 3334 2280 3340
rect 2044 3052 2096 3058
rect 1964 3012 2044 3040
rect 2044 2994 2096 3000
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 2056 2514 2084 2790
rect 2044 2508 2096 2514
rect 2044 2450 2096 2456
rect 2240 2446 2268 3334
rect 2424 3058 2452 7346
rect 2516 7206 2544 8486
rect 2824 8188 3132 8197
rect 2824 8186 2830 8188
rect 2886 8186 2910 8188
rect 2966 8186 2990 8188
rect 3046 8186 3070 8188
rect 3126 8186 3132 8188
rect 2886 8134 2888 8186
rect 3068 8134 3070 8186
rect 2824 8132 2830 8134
rect 2886 8132 2910 8134
rect 2966 8132 2990 8134
rect 3046 8132 3070 8134
rect 3126 8132 3132 8134
rect 2824 8123 3132 8132
rect 3160 8090 3188 8502
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3148 7812 3200 7818
rect 3148 7754 3200 7760
rect 3160 7478 3188 7754
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3252 7206 3280 8298
rect 3436 8072 3464 12650
rect 3712 12374 3740 14962
rect 3792 14952 3844 14958
rect 3792 14894 3844 14900
rect 3804 14482 3832 14894
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3804 13870 3832 14418
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 3804 13258 3832 13806
rect 3792 13252 3844 13258
rect 3792 13194 3844 13200
rect 3804 12918 3832 13194
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 3896 12434 3924 15263
rect 3988 14958 4016 16118
rect 4068 16040 4120 16046
rect 4066 16008 4068 16017
rect 4120 16008 4122 16017
rect 4172 15978 4200 16458
rect 4264 16250 4292 17138
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4344 16108 4396 16114
rect 4344 16050 4396 16056
rect 4066 15943 4122 15952
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 3976 14952 4028 14958
rect 3976 14894 4028 14900
rect 4172 14278 4200 15914
rect 4356 15910 4384 16050
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4448 15706 4476 17206
rect 4710 17167 4712 17176
rect 4764 17167 4766 17176
rect 4712 17138 4764 17144
rect 4528 16584 4580 16590
rect 4526 16552 4528 16561
rect 4580 16552 4582 16561
rect 4582 16510 4660 16538
rect 4526 16487 4582 16496
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4342 15600 4398 15609
rect 4252 15564 4304 15570
rect 4342 15535 4398 15544
rect 4252 15506 4304 15512
rect 4264 15026 4292 15506
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 4356 14822 4384 15535
rect 4540 15502 4568 15846
rect 4632 15745 4660 16510
rect 5092 16402 5120 19200
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 5368 17202 5396 17682
rect 5460 17338 5488 19200
rect 5828 17898 5856 19200
rect 5736 17870 5856 17898
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5356 17196 5408 17202
rect 5356 17138 5408 17144
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 5172 17128 5224 17134
rect 5460 17105 5488 17138
rect 5172 17070 5224 17076
rect 5446 17096 5502 17105
rect 5184 16794 5212 17070
rect 5446 17031 5502 17040
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 5172 16448 5224 16454
rect 5092 16396 5172 16402
rect 5092 16390 5224 16396
rect 5092 16374 5212 16390
rect 4698 16348 5006 16357
rect 4698 16346 4704 16348
rect 4760 16346 4784 16348
rect 4840 16346 4864 16348
rect 4920 16346 4944 16348
rect 5000 16346 5006 16348
rect 4760 16294 4762 16346
rect 4942 16294 4944 16346
rect 4698 16292 4704 16294
rect 4760 16292 4784 16294
rect 4840 16292 4864 16294
rect 4920 16292 4944 16294
rect 5000 16292 5006 16294
rect 4698 16283 5006 16292
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5172 16040 5224 16046
rect 5172 15982 5224 15988
rect 4618 15736 4674 15745
rect 4618 15671 4674 15680
rect 4528 15496 4580 15502
rect 4528 15438 4580 15444
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4632 15162 4660 15302
rect 4698 15260 5006 15269
rect 4698 15258 4704 15260
rect 4760 15258 4784 15260
rect 4840 15258 4864 15260
rect 4920 15258 4944 15260
rect 5000 15258 5006 15260
rect 4760 15206 4762 15258
rect 4942 15206 4944 15258
rect 4698 15204 4704 15206
rect 4760 15204 4784 15206
rect 4840 15204 4864 15206
rect 4920 15204 4944 15206
rect 5000 15204 5006 15206
rect 4698 15195 5006 15204
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 4436 15020 4488 15026
rect 4436 14962 4488 14968
rect 5080 15020 5132 15026
rect 5080 14962 5132 14968
rect 4344 14816 4396 14822
rect 4344 14758 4396 14764
rect 4250 14512 4306 14521
rect 4250 14447 4306 14456
rect 4264 14278 4292 14447
rect 4448 14414 4476 14962
rect 5092 14618 5120 14962
rect 5184 14958 5212 15982
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4172 13870 4200 14214
rect 4264 14006 4292 14214
rect 4252 14000 4304 14006
rect 4250 13968 4252 13977
rect 4304 13968 4306 13977
rect 4250 13903 4306 13912
rect 4160 13864 4212 13870
rect 4158 13832 4160 13841
rect 4212 13832 4214 13841
rect 4158 13767 4214 13776
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4080 12918 4108 13466
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 3804 12406 3924 12434
rect 3700 12368 3752 12374
rect 3700 12310 3752 12316
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3528 11218 3556 11630
rect 3516 11212 3568 11218
rect 3516 11154 3568 11160
rect 3528 10606 3556 11154
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3528 10198 3556 10542
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3528 9586 3556 9998
rect 3804 9602 3832 12406
rect 4172 12306 4200 12786
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 3884 12232 3936 12238
rect 3882 12200 3884 12209
rect 3936 12200 3938 12209
rect 3882 12135 3938 12144
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3988 11830 4016 12038
rect 4172 11898 4200 12242
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 3988 11150 4016 11766
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 4080 11286 4108 11698
rect 4068 11280 4120 11286
rect 4068 11222 4120 11228
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 4080 10826 4108 11222
rect 4356 11218 4384 11834
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 3988 10798 4108 10826
rect 4356 10810 4384 11154
rect 4344 10804 4396 10810
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3620 9574 3832 9602
rect 3884 9648 3936 9654
rect 3884 9590 3936 9596
rect 3528 9042 3556 9522
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3516 8560 3568 8566
rect 3516 8502 3568 8508
rect 3344 8044 3464 8072
rect 2504 7200 2556 7206
rect 2504 7142 2556 7148
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 2516 6662 2544 7142
rect 2824 7100 3132 7109
rect 2824 7098 2830 7100
rect 2886 7098 2910 7100
rect 2966 7098 2990 7100
rect 3046 7098 3070 7100
rect 3126 7098 3132 7100
rect 2886 7046 2888 7098
rect 3068 7046 3070 7098
rect 2824 7044 2830 7046
rect 2886 7044 2910 7046
rect 2966 7044 2990 7046
rect 3046 7044 3070 7046
rect 3126 7044 3132 7046
rect 2824 7035 3132 7044
rect 3344 6866 3372 8044
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3436 7342 3464 7890
rect 3528 7732 3556 8502
rect 3620 7857 3648 9574
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3606 7848 3662 7857
rect 3606 7783 3662 7792
rect 3608 7744 3660 7750
rect 3528 7704 3608 7732
rect 3608 7686 3660 7692
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2516 5681 2544 6598
rect 2608 6322 2636 6734
rect 2688 6724 2740 6730
rect 3332 6724 3384 6730
rect 2688 6666 2740 6672
rect 3252 6684 3332 6712
rect 2596 6316 2648 6322
rect 2596 6258 2648 6264
rect 2596 6180 2648 6186
rect 2596 6122 2648 6128
rect 2502 5672 2558 5681
rect 2502 5607 2558 5616
rect 2502 5264 2558 5273
rect 2502 5199 2504 5208
rect 2556 5199 2558 5208
rect 2504 5170 2556 5176
rect 2608 4690 2636 6122
rect 2700 4690 2728 6666
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 2792 6390 2820 6598
rect 2780 6384 2832 6390
rect 2780 6326 2832 6332
rect 2780 6248 2832 6254
rect 2778 6216 2780 6225
rect 2832 6216 2834 6225
rect 2778 6151 2834 6160
rect 2824 6012 3132 6021
rect 2824 6010 2830 6012
rect 2886 6010 2910 6012
rect 2966 6010 2990 6012
rect 3046 6010 3070 6012
rect 3126 6010 3132 6012
rect 2886 5958 2888 6010
rect 3068 5958 3070 6010
rect 2824 5956 2830 5958
rect 2886 5956 2910 5958
rect 2966 5956 2990 5958
rect 3046 5956 3070 5958
rect 3126 5956 3132 5958
rect 2824 5947 3132 5956
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2792 5030 2820 5646
rect 2884 5166 2912 5714
rect 3068 5710 3096 5850
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 3160 5370 3188 6598
rect 3252 6254 3280 6684
rect 3332 6666 3384 6672
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3240 6248 3292 6254
rect 3240 6190 3292 6196
rect 3252 6118 3280 6190
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 3146 5128 3202 5137
rect 3146 5063 3202 5072
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2824 4924 3132 4933
rect 2824 4922 2830 4924
rect 2886 4922 2910 4924
rect 2966 4922 2990 4924
rect 3046 4922 3070 4924
rect 3126 4922 3132 4924
rect 2886 4870 2888 4922
rect 3068 4870 3070 4922
rect 2824 4868 2830 4870
rect 2886 4868 2910 4870
rect 2966 4868 2990 4870
rect 3046 4868 3070 4870
rect 3126 4868 3132 4870
rect 2824 4859 3132 4868
rect 3054 4720 3110 4729
rect 2596 4684 2648 4690
rect 2596 4626 2648 4632
rect 2688 4684 2740 4690
rect 3054 4655 3110 4664
rect 2688 4626 2740 4632
rect 2504 4480 2556 4486
rect 2504 4422 2556 4428
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 1952 2304 2004 2310
rect 1952 2246 2004 2252
rect 2320 2304 2372 2310
rect 2320 2246 2372 2252
rect 1596 800 1624 2246
rect 1964 800 1992 2246
rect 2332 800 2360 2246
rect 2516 1465 2544 4422
rect 2608 4078 2636 4626
rect 2700 4486 2728 4626
rect 2778 4584 2834 4593
rect 2778 4519 2834 4528
rect 2792 4486 2820 4519
rect 3068 4486 3096 4655
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 3068 4162 3096 4422
rect 3160 4282 3188 5063
rect 3252 4690 3280 6054
rect 3436 5914 3464 6598
rect 3528 6390 3556 7210
rect 3620 7206 3648 7686
rect 3608 7200 3660 7206
rect 3608 7142 3660 7148
rect 3516 6384 3568 6390
rect 3516 6326 3568 6332
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3528 5574 3556 6326
rect 3620 6225 3648 7142
rect 3606 6216 3662 6225
rect 3606 6151 3662 6160
rect 3424 5568 3476 5574
rect 3330 5536 3386 5545
rect 3424 5510 3476 5516
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 3330 5471 3386 5480
rect 3344 5250 3372 5471
rect 3436 5352 3464 5510
rect 3516 5364 3568 5370
rect 3436 5324 3516 5352
rect 3516 5306 3568 5312
rect 3344 5222 3464 5250
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 2700 4146 2820 4162
rect 2700 4140 2832 4146
rect 2700 4134 2780 4140
rect 2596 4072 2648 4078
rect 2596 4014 2648 4020
rect 2700 3942 2728 4134
rect 3068 4134 3188 4162
rect 2780 4082 2832 4088
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2700 3126 2728 3878
rect 2824 3836 3132 3845
rect 2824 3834 2830 3836
rect 2886 3834 2910 3836
rect 2966 3834 2990 3836
rect 3046 3834 3070 3836
rect 3126 3834 3132 3836
rect 2886 3782 2888 3834
rect 3068 3782 3070 3834
rect 2824 3780 2830 3782
rect 2886 3780 2910 3782
rect 2966 3780 2990 3782
rect 3046 3780 3070 3782
rect 3126 3780 3132 3782
rect 2824 3771 3132 3780
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2688 3120 2740 3126
rect 2688 3062 2740 3068
rect 2792 3058 2820 3674
rect 3160 3482 3188 4134
rect 3252 3602 3280 4626
rect 3344 4282 3372 5102
rect 3436 4486 3464 5222
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3712 4282 3740 8910
rect 3804 6882 3832 9454
rect 3896 9110 3924 9590
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3896 8498 3924 9046
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3896 8090 3924 8434
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 3988 7818 4016 10798
rect 4344 10746 4396 10752
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 4080 9586 4108 10678
rect 4356 10606 4384 10746
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4172 10062 4200 10542
rect 4448 10538 4476 14350
rect 4698 14172 5006 14181
rect 4698 14170 4704 14172
rect 4760 14170 4784 14172
rect 4840 14170 4864 14172
rect 4920 14170 4944 14172
rect 5000 14170 5006 14172
rect 4760 14118 4762 14170
rect 4942 14118 4944 14170
rect 4698 14116 4704 14118
rect 4760 14116 4784 14118
rect 4840 14116 4864 14118
rect 4920 14116 4944 14118
rect 5000 14116 5006 14118
rect 4698 14107 5006 14116
rect 5184 14006 5212 14894
rect 5276 14249 5304 16050
rect 5460 15706 5488 16934
rect 5632 16516 5684 16522
rect 5632 16458 5684 16464
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5356 15632 5408 15638
rect 5356 15574 5408 15580
rect 5368 15162 5396 15574
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5368 14414 5396 15098
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5262 14240 5318 14249
rect 5262 14175 5318 14184
rect 5460 14074 5488 15506
rect 5552 14890 5580 15846
rect 5644 15434 5672 16458
rect 5736 16454 5764 17870
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5736 15570 5764 16050
rect 5828 15706 5856 17138
rect 6196 17066 6224 19200
rect 6564 17270 6592 19200
rect 6932 17338 6960 19200
rect 7012 17604 7064 17610
rect 7012 17546 7064 17552
rect 6920 17332 6972 17338
rect 6920 17274 6972 17280
rect 6552 17264 6604 17270
rect 6552 17206 6604 17212
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6184 17060 6236 17066
rect 6184 17002 6236 17008
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5908 16040 5960 16046
rect 5908 15982 5960 15988
rect 5816 15700 5868 15706
rect 5816 15642 5868 15648
rect 5724 15564 5776 15570
rect 5724 15506 5776 15512
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5632 15428 5684 15434
rect 5632 15370 5684 15376
rect 5630 15056 5686 15065
rect 5630 14991 5686 15000
rect 5644 14890 5672 14991
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5540 14884 5592 14890
rect 5540 14826 5592 14832
rect 5632 14884 5684 14890
rect 5632 14826 5684 14832
rect 5736 14618 5764 14894
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5828 14498 5856 15438
rect 5920 14958 5948 15982
rect 6012 15162 6040 16186
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6104 16017 6132 16050
rect 6090 16008 6146 16017
rect 6090 15943 6146 15952
rect 6288 15570 6316 16730
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 6380 15706 6408 16390
rect 6368 15700 6420 15706
rect 6368 15642 6420 15648
rect 6276 15564 6328 15570
rect 6276 15506 6328 15512
rect 6092 15428 6144 15434
rect 6092 15370 6144 15376
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 5908 14952 5960 14958
rect 5908 14894 5960 14900
rect 5736 14470 5856 14498
rect 5920 14482 5948 14894
rect 5908 14476 5960 14482
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4540 13326 4568 13670
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4698 13084 5006 13093
rect 4698 13082 4704 13084
rect 4760 13082 4784 13084
rect 4840 13082 4864 13084
rect 4920 13082 4944 13084
rect 5000 13082 5006 13084
rect 4760 13030 4762 13082
rect 4942 13030 4944 13082
rect 4698 13028 4704 13030
rect 4760 13028 4784 13030
rect 4840 13028 4864 13030
rect 4920 13028 4944 13030
rect 5000 13028 5006 13030
rect 4698 13019 5006 13028
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4816 12238 4844 12718
rect 5264 12368 5316 12374
rect 5264 12310 5316 12316
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4540 11830 4568 12106
rect 4698 11996 5006 12005
rect 4698 11994 4704 11996
rect 4760 11994 4784 11996
rect 4840 11994 4864 11996
rect 4920 11994 4944 11996
rect 5000 11994 5006 11996
rect 4760 11942 4762 11994
rect 4942 11942 4944 11994
rect 4698 11940 4704 11942
rect 4760 11940 4784 11942
rect 4840 11940 4864 11942
rect 4920 11940 4944 11942
rect 5000 11940 5006 11942
rect 4698 11931 5006 11940
rect 4528 11824 4580 11830
rect 4528 11766 4580 11772
rect 4540 10810 4568 11766
rect 4698 10908 5006 10917
rect 4698 10906 4704 10908
rect 4760 10906 4784 10908
rect 4840 10906 4864 10908
rect 4920 10906 4944 10908
rect 5000 10906 5006 10908
rect 4760 10854 4762 10906
rect 4942 10854 4944 10906
rect 4698 10852 4704 10854
rect 4760 10852 4784 10854
rect 4840 10852 4864 10854
rect 4920 10852 4944 10854
rect 5000 10852 5006 10854
rect 4698 10843 5006 10852
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4436 10532 4488 10538
rect 4436 10474 4488 10480
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 4080 8634 4108 9522
rect 4264 9466 4292 10066
rect 4264 9438 4384 9466
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4264 8498 4292 9318
rect 4356 8906 4384 9438
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4356 8634 4384 8842
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4080 8242 4108 8298
rect 4448 8242 4476 10474
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4080 8214 4476 8242
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 3988 7478 4016 7754
rect 3976 7472 4028 7478
rect 3976 7414 4028 7420
rect 3804 6854 4016 6882
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6458 3832 6598
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3896 5574 3924 6734
rect 3988 5681 4016 6854
rect 4080 5778 4108 7754
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4172 6934 4200 7346
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4068 5772 4120 5778
rect 4068 5714 4120 5720
rect 3974 5672 4030 5681
rect 3974 5607 4030 5616
rect 4160 5636 4212 5642
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3804 5001 3832 5510
rect 3896 5234 3924 5510
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3790 4992 3846 5001
rect 3790 4927 3846 4936
rect 3896 4758 3924 5170
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3712 3942 3740 4218
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 3436 3534 3464 3878
rect 3712 3670 3740 3878
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 3424 3528 3476 3534
rect 3160 3454 3280 3482
rect 3424 3470 3476 3476
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 3160 3194 3188 3334
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 3252 2961 3280 3454
rect 3238 2952 3294 2961
rect 2688 2916 2740 2922
rect 2688 2858 2740 2864
rect 3148 2916 3200 2922
rect 3238 2887 3294 2896
rect 3148 2858 3200 2864
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 2608 2446 2636 2790
rect 2700 2530 2728 2858
rect 2824 2748 3132 2757
rect 2824 2746 2830 2748
rect 2886 2746 2910 2748
rect 2966 2746 2990 2748
rect 3046 2746 3070 2748
rect 3126 2746 3132 2748
rect 2886 2694 2888 2746
rect 3068 2694 3070 2746
rect 2824 2692 2830 2694
rect 2886 2692 2910 2694
rect 2966 2692 2990 2694
rect 3046 2692 3070 2694
rect 3126 2692 3132 2694
rect 2824 2683 3132 2692
rect 2700 2502 2820 2530
rect 2792 2446 2820 2502
rect 3160 2446 3188 2858
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 2688 2304 2740 2310
rect 2688 2246 2740 2252
rect 2502 1456 2558 1465
rect 2502 1391 2558 1400
rect 2700 800 2728 2246
rect 3252 1442 3280 2790
rect 3804 2446 3832 4422
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3896 3058 3924 3334
rect 3988 3126 4016 5607
rect 4160 5578 4212 5584
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 4080 5030 4108 5102
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4214 4108 4966
rect 4172 4826 4200 5578
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 4172 3641 4200 4558
rect 4158 3632 4214 3641
rect 4158 3567 4214 3576
rect 4264 3534 4292 8214
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4448 7206 4476 7822
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4356 6390 4384 7142
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 4356 4146 4384 6326
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4448 5234 4476 5510
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4540 4146 4568 8774
rect 4632 7274 4660 10542
rect 4698 9820 5006 9829
rect 4698 9818 4704 9820
rect 4760 9818 4784 9820
rect 4840 9818 4864 9820
rect 4920 9818 4944 9820
rect 5000 9818 5006 9820
rect 4760 9766 4762 9818
rect 4942 9766 4944 9818
rect 4698 9764 4704 9766
rect 4760 9764 4784 9766
rect 4840 9764 4864 9766
rect 4920 9764 4944 9766
rect 5000 9764 5006 9766
rect 4698 9755 5006 9764
rect 4698 8732 5006 8741
rect 4698 8730 4704 8732
rect 4760 8730 4784 8732
rect 4840 8730 4864 8732
rect 4920 8730 4944 8732
rect 5000 8730 5006 8732
rect 4760 8678 4762 8730
rect 4942 8678 4944 8730
rect 4698 8676 4704 8678
rect 4760 8676 4784 8678
rect 4840 8676 4864 8678
rect 4920 8676 4944 8678
rect 5000 8676 5006 8678
rect 4698 8667 5006 8676
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 7886 5212 8230
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 4698 7644 5006 7653
rect 4698 7642 4704 7644
rect 4760 7642 4784 7644
rect 4840 7642 4864 7644
rect 4920 7642 4944 7644
rect 5000 7642 5006 7644
rect 4760 7590 4762 7642
rect 4942 7590 4944 7642
rect 4698 7588 4704 7590
rect 4760 7588 4784 7590
rect 4840 7588 4864 7590
rect 4920 7588 4944 7590
rect 5000 7588 5006 7590
rect 4698 7579 5006 7588
rect 5184 7478 5212 7822
rect 5172 7472 5224 7478
rect 5172 7414 5224 7420
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4698 6556 5006 6565
rect 4698 6554 4704 6556
rect 4760 6554 4784 6556
rect 4840 6554 4864 6556
rect 4920 6554 4944 6556
rect 5000 6554 5006 6556
rect 4760 6502 4762 6554
rect 4942 6502 4944 6554
rect 4698 6500 4704 6502
rect 4760 6500 4784 6502
rect 4840 6500 4864 6502
rect 4920 6500 4944 6502
rect 5000 6500 5006 6502
rect 4698 6491 5006 6500
rect 5276 6202 5304 12310
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5460 11150 5488 11630
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5644 10742 5672 14350
rect 5736 14346 5764 14470
rect 5908 14418 5960 14424
rect 5724 14340 5776 14346
rect 5724 14282 5776 14288
rect 5736 12102 5764 14282
rect 5816 13932 5868 13938
rect 5920 13920 5948 14418
rect 6012 14346 6040 15098
rect 6000 14340 6052 14346
rect 6000 14282 6052 14288
rect 5868 13892 5948 13920
rect 5816 13874 5868 13880
rect 5920 13530 5948 13892
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 6012 13326 6040 13874
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5828 10742 5856 11290
rect 6104 11082 6132 15370
rect 6182 15192 6238 15201
rect 6182 15127 6238 15136
rect 6196 15094 6224 15127
rect 6472 15094 6500 17138
rect 6572 16892 6880 16901
rect 6572 16890 6578 16892
rect 6634 16890 6658 16892
rect 6714 16890 6738 16892
rect 6794 16890 6818 16892
rect 6874 16890 6880 16892
rect 6634 16838 6636 16890
rect 6816 16838 6818 16890
rect 6572 16836 6578 16838
rect 6634 16836 6658 16838
rect 6714 16836 6738 16838
rect 6794 16836 6818 16838
rect 6874 16836 6880 16838
rect 6572 16827 6880 16836
rect 7024 16640 7052 17546
rect 7300 17134 7328 19200
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7392 17338 7420 17478
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 6932 16612 7052 16640
rect 7102 16688 7158 16697
rect 7102 16623 7158 16632
rect 7196 16652 7248 16658
rect 6932 16538 6960 16612
rect 7116 16590 7144 16623
rect 7196 16594 7248 16600
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 6840 16510 6960 16538
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 6840 16250 6868 16510
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6920 16176 6972 16182
rect 6920 16118 6972 16124
rect 6572 15804 6880 15813
rect 6572 15802 6578 15804
rect 6634 15802 6658 15804
rect 6714 15802 6738 15804
rect 6794 15802 6818 15804
rect 6874 15802 6880 15804
rect 6634 15750 6636 15802
rect 6816 15750 6818 15802
rect 6572 15748 6578 15750
rect 6634 15748 6658 15750
rect 6714 15748 6738 15750
rect 6794 15748 6818 15750
rect 6874 15748 6880 15750
rect 6572 15739 6880 15748
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 6840 15162 6868 15302
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6184 15088 6236 15094
rect 6184 15030 6236 15036
rect 6460 15088 6512 15094
rect 6932 15065 6960 16118
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 6460 15030 6512 15036
rect 6918 15056 6974 15065
rect 6828 15020 6880 15026
rect 6918 14991 6974 15000
rect 6828 14962 6880 14968
rect 6840 14906 6868 14962
rect 6840 14878 6960 14906
rect 6460 14816 6512 14822
rect 6288 14776 6460 14804
rect 6288 14414 6316 14776
rect 6460 14758 6512 14764
rect 6572 14716 6880 14725
rect 6572 14714 6578 14716
rect 6634 14714 6658 14716
rect 6714 14714 6738 14716
rect 6794 14714 6818 14716
rect 6874 14714 6880 14716
rect 6634 14662 6636 14714
rect 6816 14662 6818 14714
rect 6572 14660 6578 14662
rect 6634 14660 6658 14662
rect 6714 14660 6738 14662
rect 6794 14660 6818 14662
rect 6874 14660 6880 14662
rect 6572 14651 6880 14660
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 6184 14340 6236 14346
rect 6184 14282 6236 14288
rect 6196 13512 6224 14282
rect 6276 13524 6328 13530
rect 6196 13484 6276 13512
rect 6276 13466 6328 13472
rect 6380 13190 6408 14418
rect 6932 14346 6960 14878
rect 7024 14618 7052 16050
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 7116 14958 7144 15438
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 6460 14272 6512 14278
rect 6460 14214 6512 14220
rect 6472 13938 6500 14214
rect 6840 14006 6868 14282
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 6572 13628 6880 13637
rect 6572 13626 6578 13628
rect 6634 13626 6658 13628
rect 6714 13626 6738 13628
rect 6794 13626 6818 13628
rect 6874 13626 6880 13628
rect 6634 13574 6636 13626
rect 6816 13574 6818 13626
rect 6572 13572 6578 13574
rect 6634 13572 6658 13574
rect 6714 13572 6738 13574
rect 6794 13572 6818 13574
rect 6874 13572 6880 13574
rect 6572 13563 6880 13572
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6380 12442 6408 13126
rect 6656 12986 6684 13194
rect 6644 12980 6696 12986
rect 6472 12940 6644 12968
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6472 12238 6500 12940
rect 6644 12922 6696 12928
rect 6572 12540 6880 12549
rect 6572 12538 6578 12540
rect 6634 12538 6658 12540
rect 6714 12538 6738 12540
rect 6794 12538 6818 12540
rect 6874 12538 6880 12540
rect 6634 12486 6636 12538
rect 6816 12486 6818 12538
rect 6572 12484 6578 12486
rect 6634 12484 6658 12486
rect 6714 12484 6738 12486
rect 6794 12484 6818 12486
rect 6874 12484 6880 12486
rect 6572 12475 6880 12484
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6572 11452 6880 11461
rect 6572 11450 6578 11452
rect 6634 11450 6658 11452
rect 6714 11450 6738 11452
rect 6794 11450 6818 11452
rect 6874 11450 6880 11452
rect 6634 11398 6636 11450
rect 6816 11398 6818 11450
rect 6572 11396 6578 11398
rect 6634 11396 6658 11398
rect 6714 11396 6738 11398
rect 6794 11396 6818 11398
rect 6874 11396 6880 11398
rect 6572 11387 6880 11396
rect 6092 11076 6144 11082
rect 6092 11018 6144 11024
rect 6104 10810 6132 11018
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 5632 10736 5684 10742
rect 5632 10678 5684 10684
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 7116 10674 7144 14894
rect 7208 14498 7236 16594
rect 7300 15570 7328 16594
rect 7380 16584 7432 16590
rect 7484 16572 7512 17614
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7576 16697 7604 17274
rect 7668 17066 7696 19200
rect 8036 17542 8064 19200
rect 8208 17604 8260 17610
rect 8208 17546 8260 17552
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 7932 17196 7984 17202
rect 7932 17138 7984 17144
rect 7656 17060 7708 17066
rect 7656 17002 7708 17008
rect 7944 16794 7972 17138
rect 8036 16998 8064 17274
rect 8220 17218 8248 17546
rect 8404 17524 8432 19200
rect 8312 17496 8432 17524
rect 8772 17524 8800 19200
rect 8772 17496 8892 17524
rect 8312 17338 8340 17496
rect 8446 17436 8754 17445
rect 8446 17434 8452 17436
rect 8508 17434 8532 17436
rect 8588 17434 8612 17436
rect 8668 17434 8692 17436
rect 8748 17434 8754 17436
rect 8508 17382 8510 17434
rect 8690 17382 8692 17434
rect 8446 17380 8452 17382
rect 8508 17380 8532 17382
rect 8588 17380 8612 17382
rect 8668 17380 8692 17382
rect 8748 17380 8754 17382
rect 8446 17371 8754 17380
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8220 17190 8432 17218
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 8024 16992 8076 16998
rect 8024 16934 8076 16940
rect 8036 16794 8064 16934
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 7748 16720 7800 16726
rect 7562 16688 7618 16697
rect 7562 16623 7618 16632
rect 7668 16680 7748 16708
rect 7432 16544 7512 16572
rect 7380 16526 7432 16532
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7392 15434 7420 16526
rect 7668 16522 7696 16680
rect 7748 16662 7800 16668
rect 8220 16658 8248 17070
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 7746 16552 7802 16561
rect 7656 16516 7708 16522
rect 7746 16487 7802 16496
rect 7932 16516 7984 16522
rect 7656 16458 7708 16464
rect 7760 16250 7788 16487
rect 7932 16458 7984 16464
rect 7748 16244 7800 16250
rect 7748 16186 7800 16192
rect 7656 16040 7708 16046
rect 7656 15982 7708 15988
rect 7760 15994 7788 16186
rect 7944 16182 7972 16458
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 8128 16250 8156 16390
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 7932 16176 7984 16182
rect 7932 16118 7984 16124
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 7564 15904 7616 15910
rect 7668 15881 7696 15982
rect 7760 15966 7972 15994
rect 7564 15846 7616 15852
rect 7654 15872 7710 15881
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7380 15428 7432 15434
rect 7380 15370 7432 15376
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7300 14618 7328 14962
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7208 14470 7328 14498
rect 7194 14376 7250 14385
rect 7194 14311 7250 14320
rect 7208 13977 7236 14311
rect 7194 13968 7250 13977
rect 7194 13903 7250 13912
rect 7300 11354 7328 14470
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5920 10062 5948 10406
rect 6572 10364 6880 10373
rect 6572 10362 6578 10364
rect 6634 10362 6658 10364
rect 6714 10362 6738 10364
rect 6794 10362 6818 10364
rect 6874 10362 6880 10364
rect 6634 10310 6636 10362
rect 6816 10310 6818 10362
rect 6572 10308 6578 10310
rect 6634 10308 6658 10310
rect 6714 10308 6738 10310
rect 6794 10308 6818 10310
rect 6874 10308 6880 10310
rect 6572 10299 6880 10308
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 5920 9586 5948 9998
rect 7208 9722 7236 9998
rect 7300 9926 7328 11290
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7196 9716 7248 9722
rect 7392 9674 7420 15370
rect 7484 15366 7512 15642
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7484 14278 7512 15302
rect 7576 15162 7604 15846
rect 7654 15807 7710 15816
rect 7840 15564 7892 15570
rect 7840 15506 7892 15512
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7484 13818 7512 14214
rect 7576 14006 7604 14894
rect 7668 14618 7696 15030
rect 7760 15026 7788 15098
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7748 14884 7800 14890
rect 7748 14826 7800 14832
rect 7852 14872 7880 15506
rect 7944 15042 7972 15966
rect 8128 15094 8156 16050
rect 8220 15502 8248 16594
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 8220 15201 8248 15302
rect 8206 15192 8262 15201
rect 8206 15127 8262 15136
rect 8116 15088 8168 15094
rect 7944 15014 8064 15042
rect 8116 15030 8168 15036
rect 7932 14884 7984 14890
rect 7852 14844 7932 14872
rect 7760 14657 7788 14826
rect 7746 14648 7802 14657
rect 7656 14612 7708 14618
rect 7746 14583 7802 14592
rect 7656 14554 7708 14560
rect 7852 14482 7880 14844
rect 7932 14826 7984 14832
rect 7840 14476 7892 14482
rect 7840 14418 7892 14424
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7564 14000 7616 14006
rect 7564 13942 7616 13948
rect 7484 13790 7604 13818
rect 7576 12434 7604 13790
rect 7668 13326 7696 14010
rect 7656 13320 7708 13326
rect 7656 13262 7708 13268
rect 7852 12442 7880 14418
rect 8036 14074 8064 15014
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8116 14952 8168 14958
rect 8116 14894 8168 14900
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8128 14006 8156 14894
rect 8220 14074 8248 14962
rect 8312 14618 8340 17002
rect 8404 16454 8432 17190
rect 8864 16590 8892 17496
rect 8942 17232 8998 17241
rect 8942 17167 8998 17176
rect 8956 16726 8984 17167
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 8944 16720 8996 16726
rect 8944 16662 8996 16668
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 9048 16538 9076 16934
rect 9140 16674 9168 19200
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9310 16824 9366 16833
rect 9310 16759 9366 16768
rect 9324 16726 9352 16759
rect 9312 16720 9364 16726
rect 9140 16646 9260 16674
rect 9312 16662 9364 16668
rect 9232 16590 9260 16646
rect 9128 16584 9180 16590
rect 9126 16552 9128 16561
rect 9220 16584 9272 16590
rect 9180 16552 9182 16561
rect 9048 16510 9126 16538
rect 9220 16526 9272 16532
rect 9126 16487 9182 16496
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8852 16448 8904 16454
rect 8852 16390 8904 16396
rect 8446 16348 8754 16357
rect 8446 16346 8452 16348
rect 8508 16346 8532 16348
rect 8588 16346 8612 16348
rect 8668 16346 8692 16348
rect 8748 16346 8754 16348
rect 8508 16294 8510 16346
rect 8690 16294 8692 16346
rect 8446 16292 8452 16294
rect 8508 16292 8532 16294
rect 8588 16292 8612 16294
rect 8668 16292 8692 16294
rect 8748 16292 8754 16294
rect 8446 16283 8754 16292
rect 8864 16266 8892 16390
rect 8864 16238 9076 16266
rect 8944 16108 8996 16114
rect 8944 16050 8996 16056
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 8496 15910 8524 15982
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 8404 15638 8432 15846
rect 8392 15632 8444 15638
rect 8392 15574 8444 15580
rect 8392 15360 8444 15366
rect 8373 15308 8392 15348
rect 8373 15302 8444 15308
rect 8373 15144 8401 15302
rect 8446 15260 8754 15269
rect 8446 15258 8452 15260
rect 8508 15258 8532 15260
rect 8588 15258 8612 15260
rect 8668 15258 8692 15260
rect 8748 15258 8754 15260
rect 8508 15206 8510 15258
rect 8690 15206 8692 15258
rect 8446 15204 8452 15206
rect 8508 15204 8532 15206
rect 8588 15204 8612 15206
rect 8668 15204 8692 15206
rect 8748 15204 8754 15206
rect 8446 15195 8754 15204
rect 8864 15162 8892 15982
rect 8956 15706 8984 16050
rect 8944 15700 8996 15706
rect 8944 15642 8996 15648
rect 9048 15502 9076 16238
rect 9128 16176 9180 16182
rect 9128 16118 9180 16124
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8852 15156 8904 15162
rect 8373 15116 8432 15144
rect 8404 14822 8432 15116
rect 8852 15098 8904 15104
rect 8760 15088 8812 15094
rect 8760 15030 8812 15036
rect 8850 15056 8906 15065
rect 8668 14884 8720 14890
rect 8668 14826 8720 14832
rect 8392 14816 8444 14822
rect 8576 14816 8628 14822
rect 8392 14758 8444 14764
rect 8574 14784 8576 14793
rect 8628 14784 8630 14793
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8404 14498 8432 14758
rect 8574 14719 8630 14728
rect 8574 14648 8630 14657
rect 8680 14634 8708 14826
rect 8630 14606 8708 14634
rect 8772 14618 8800 15030
rect 8850 14991 8906 15000
rect 8760 14612 8812 14618
rect 8574 14583 8630 14592
rect 8760 14554 8812 14560
rect 8312 14470 8432 14498
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 7840 12436 7892 12442
rect 7576 12406 7696 12434
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7196 9658 7248 9664
rect 7300 9646 7420 9674
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5920 9382 5948 9522
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5920 8974 5948 9318
rect 6572 9276 6880 9285
rect 6572 9274 6578 9276
rect 6634 9274 6658 9276
rect 6714 9274 6738 9276
rect 6794 9274 6818 9276
rect 6874 9274 6880 9276
rect 6634 9222 6636 9274
rect 6816 9222 6818 9274
rect 6572 9220 6578 9222
rect 6634 9220 6658 9222
rect 6714 9220 6738 9222
rect 6794 9220 6818 9222
rect 6874 9220 6880 9222
rect 6572 9211 6880 9220
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5460 7410 5488 7686
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 5092 6174 5304 6202
rect 4724 5642 4752 6122
rect 5092 5817 5120 6174
rect 5172 6112 5224 6118
rect 5224 6072 5304 6100
rect 5172 6054 5224 6060
rect 5078 5808 5134 5817
rect 5078 5743 5134 5752
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4698 5468 5006 5477
rect 4698 5466 4704 5468
rect 4760 5466 4784 5468
rect 4840 5466 4864 5468
rect 4920 5466 4944 5468
rect 5000 5466 5006 5468
rect 4760 5414 4762 5466
rect 4942 5414 4944 5466
rect 4698 5412 4704 5414
rect 4760 5412 4784 5414
rect 4840 5412 4864 5414
rect 4920 5412 4944 5414
rect 5000 5412 5006 5414
rect 4698 5403 5006 5412
rect 5092 5370 5120 5743
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5092 5166 5120 5306
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4068 3528 4120 3534
rect 4066 3496 4068 3505
rect 4252 3528 4304 3534
rect 4120 3496 4122 3505
rect 4252 3470 4304 3476
rect 4066 3431 4122 3440
rect 3976 3120 4028 3126
rect 3976 3062 4028 3068
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 4356 2990 4384 4082
rect 4434 3632 4490 3641
rect 4434 3567 4490 3576
rect 4528 3596 4580 3602
rect 4448 3466 4476 3567
rect 4528 3538 4580 3544
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 4540 3194 4568 3538
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4632 3058 4660 4966
rect 4802 4584 4858 4593
rect 4802 4519 4858 4528
rect 4816 4486 4844 4519
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4698 4380 5006 4389
rect 4698 4378 4704 4380
rect 4760 4378 4784 4380
rect 4840 4378 4864 4380
rect 4920 4378 4944 4380
rect 5000 4378 5006 4380
rect 4760 4326 4762 4378
rect 4942 4326 4944 4378
rect 4698 4324 4704 4326
rect 4760 4324 4784 4326
rect 4840 4324 4864 4326
rect 4920 4324 4944 4326
rect 5000 4324 5006 4326
rect 4698 4315 5006 4324
rect 5092 3534 5120 4422
rect 5184 4282 5212 5238
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5184 3398 5212 3674
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 4698 3292 5006 3301
rect 4698 3290 4704 3292
rect 4760 3290 4784 3292
rect 4840 3290 4864 3292
rect 4920 3290 4944 3292
rect 5000 3290 5006 3292
rect 4760 3238 4762 3290
rect 4942 3238 4944 3290
rect 4698 3236 4704 3238
rect 4760 3236 4784 3238
rect 4840 3236 4864 3238
rect 4920 3236 4944 3238
rect 5000 3236 5006 3238
rect 4698 3227 5006 3236
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 5184 2990 5212 3130
rect 5276 3058 5304 6072
rect 5460 5370 5488 7142
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5552 6322 5580 6598
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5552 5030 5580 5238
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5644 4826 5672 5170
rect 5736 5166 5764 8774
rect 5920 8634 5948 8910
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 5828 5914 5856 7346
rect 6288 6458 6316 8502
rect 6572 8188 6880 8197
rect 6572 8186 6578 8188
rect 6634 8186 6658 8188
rect 6714 8186 6738 8188
rect 6794 8186 6818 8188
rect 6874 8186 6880 8188
rect 6634 8134 6636 8186
rect 6816 8134 6818 8186
rect 6572 8132 6578 8134
rect 6634 8132 6658 8134
rect 6714 8132 6738 8134
rect 6794 8132 6818 8134
rect 6874 8132 6880 8134
rect 6572 8123 6880 8132
rect 7300 7313 7328 9646
rect 7576 9382 7604 10610
rect 7564 9376 7616 9382
rect 7564 9318 7616 9324
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7286 7304 7342 7313
rect 7286 7239 7342 7248
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6472 6798 6500 7142
rect 6572 7100 6880 7109
rect 6572 7098 6578 7100
rect 6634 7098 6658 7100
rect 6714 7098 6738 7100
rect 6794 7098 6818 7100
rect 6874 7098 6880 7100
rect 6634 7046 6636 7098
rect 6816 7046 6818 7098
rect 6572 7044 6578 7046
rect 6634 7044 6658 7046
rect 6714 7044 6738 7046
rect 6794 7044 6818 7046
rect 6874 7044 6880 7046
rect 6572 7035 6880 7044
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5630 4720 5686 4729
rect 5630 4655 5686 4664
rect 5448 4616 5500 4622
rect 5644 4570 5672 4655
rect 5500 4564 5672 4570
rect 5448 4558 5672 4564
rect 5460 4542 5672 4558
rect 5540 4480 5592 4486
rect 5446 4448 5502 4457
rect 5540 4422 5592 4428
rect 5446 4383 5502 4392
rect 5460 4049 5488 4383
rect 5552 4282 5580 4422
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5644 4146 5672 4542
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5446 4040 5502 4049
rect 5446 3975 5502 3984
rect 5540 3732 5592 3738
rect 5460 3692 5540 3720
rect 5460 3194 5488 3692
rect 5540 3674 5592 3680
rect 5538 3632 5594 3641
rect 5538 3567 5594 3576
rect 5552 3534 5580 3567
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5540 3392 5592 3398
rect 5538 3360 5540 3369
rect 5592 3360 5594 3369
rect 5538 3295 5594 3304
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 5644 3058 5672 4082
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 5172 2984 5224 2990
rect 5172 2926 5224 2932
rect 5736 2938 5764 4218
rect 5828 3738 5856 5170
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5920 4826 5948 5102
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5816 3732 5868 3738
rect 5816 3674 5868 3680
rect 5920 2990 5948 4626
rect 6012 4146 6040 6258
rect 6288 6066 6316 6394
rect 6472 6390 6500 6734
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6472 6254 6500 6326
rect 6460 6248 6512 6254
rect 6366 6216 6422 6225
rect 6460 6190 6512 6196
rect 6366 6151 6422 6160
rect 6380 6118 6408 6151
rect 6196 6038 6316 6066
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6196 5098 6224 6038
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6288 5098 6316 5850
rect 6184 5092 6236 5098
rect 6184 5034 6236 5040
rect 6276 5092 6328 5098
rect 6276 5034 6328 5040
rect 6090 4992 6146 5001
rect 6090 4927 6146 4936
rect 6104 4622 6132 4927
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6184 4548 6236 4554
rect 6184 4490 6236 4496
rect 6196 4282 6224 4490
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6196 4146 6224 4218
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6104 3369 6132 3878
rect 6090 3360 6146 3369
rect 6090 3295 6146 3304
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 5908 2984 5960 2990
rect 5736 2910 5856 2938
rect 5908 2926 5960 2932
rect 4712 2848 4764 2854
rect 4712 2790 4764 2796
rect 5172 2848 5224 2854
rect 5724 2848 5776 2854
rect 5172 2790 5224 2796
rect 5644 2808 5724 2836
rect 4724 2446 4752 2790
rect 5184 2446 5212 2790
rect 3792 2440 3844 2446
rect 3606 2408 3662 2417
rect 3792 2382 3844 2388
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 3606 2343 3608 2352
rect 3660 2343 3662 2352
rect 3608 2314 3660 2320
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 3068 1414 3280 1442
rect 3068 800 3096 1414
rect 3436 800 3464 2246
rect 3804 800 3832 2246
rect 4172 800 4200 2246
rect 4540 800 4568 2246
rect 4698 2204 5006 2213
rect 4698 2202 4704 2204
rect 4760 2202 4784 2204
rect 4840 2202 4864 2204
rect 4920 2202 4944 2204
rect 5000 2202 5006 2204
rect 4760 2150 4762 2202
rect 4942 2150 4944 2202
rect 4698 2148 4704 2150
rect 4760 2148 4784 2150
rect 4840 2148 4864 2150
rect 4920 2148 4944 2150
rect 5000 2148 5006 2150
rect 4698 2139 5006 2148
rect 5092 1170 5120 2246
rect 4908 1142 5120 1170
rect 4908 800 4936 1142
rect 5276 800 5304 2246
rect 5644 800 5672 2808
rect 5724 2790 5776 2796
rect 5828 2774 5856 2910
rect 5828 2746 6040 2774
rect 6012 2514 6040 2746
rect 6104 2514 6132 3130
rect 6000 2508 6052 2514
rect 6000 2450 6052 2456
rect 6092 2508 6144 2514
rect 6092 2450 6144 2456
rect 6196 2446 6224 3878
rect 6288 3516 6316 5034
rect 6380 4690 6408 6054
rect 6472 5710 6500 6190
rect 6572 6012 6880 6021
rect 6572 6010 6578 6012
rect 6634 6010 6658 6012
rect 6714 6010 6738 6012
rect 6794 6010 6818 6012
rect 6874 6010 6880 6012
rect 6634 5958 6636 6010
rect 6816 5958 6818 6010
rect 6572 5956 6578 5958
rect 6634 5956 6658 5958
rect 6714 5956 6738 5958
rect 6794 5956 6818 5958
rect 6874 5956 6880 5958
rect 6572 5947 6880 5956
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6472 5370 6500 5646
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6840 5098 6868 5306
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6472 4690 6500 4966
rect 6572 4924 6880 4933
rect 6572 4922 6578 4924
rect 6634 4922 6658 4924
rect 6714 4922 6738 4924
rect 6794 4922 6818 4924
rect 6874 4922 6880 4924
rect 6634 4870 6636 4922
rect 6816 4870 6818 4922
rect 6572 4868 6578 4870
rect 6634 4868 6658 4870
rect 6714 4868 6738 4870
rect 6794 4868 6818 4870
rect 6874 4868 6880 4870
rect 6572 4859 6880 4868
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6826 4584 6882 4593
rect 6644 4548 6696 4554
rect 6826 4519 6882 4528
rect 6644 4490 6696 4496
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 6380 4146 6408 4422
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6380 3670 6408 4082
rect 6472 3738 6500 4422
rect 6656 4146 6684 4490
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6840 3924 6868 4519
rect 6932 4078 6960 5170
rect 7024 5166 7052 7142
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7208 5914 7236 6190
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 7116 5030 7144 5510
rect 7208 5302 7236 5510
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 7024 4622 7052 4966
rect 7116 4690 7144 4966
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6840 3896 6960 3924
rect 6572 3836 6880 3845
rect 6572 3834 6578 3836
rect 6634 3834 6658 3836
rect 6714 3834 6738 3836
rect 6794 3834 6818 3836
rect 6874 3834 6880 3836
rect 6634 3782 6636 3834
rect 6816 3782 6818 3834
rect 6572 3780 6578 3782
rect 6634 3780 6658 3782
rect 6714 3780 6738 3782
rect 6794 3780 6818 3782
rect 6874 3780 6880 3782
rect 6572 3771 6880 3780
rect 6460 3732 6512 3738
rect 6932 3720 6960 3896
rect 6460 3674 6512 3680
rect 6840 3692 6960 3720
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 6644 3596 6696 3602
rect 6472 3556 6644 3584
rect 6472 3516 6500 3556
rect 6644 3538 6696 3544
rect 6288 3488 6500 3516
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 6288 3194 6316 3334
rect 6840 3194 6868 3692
rect 7024 3618 7052 4218
rect 7208 4128 7236 4626
rect 7300 4554 7328 7239
rect 7392 6662 7420 8434
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7392 5234 7420 6598
rect 7484 5710 7512 8298
rect 7668 6390 7696 12406
rect 7840 12378 7892 12384
rect 7852 9654 7880 12378
rect 8024 10464 8076 10470
rect 8024 10406 8076 10412
rect 8036 9994 8064 10406
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 7840 9648 7892 9654
rect 7840 9590 7892 9596
rect 7746 9480 7802 9489
rect 7746 9415 7802 9424
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7562 5944 7618 5953
rect 7562 5879 7618 5888
rect 7576 5846 7604 5879
rect 7760 5846 7788 9415
rect 8036 9382 8064 9930
rect 8312 9674 8340 14470
rect 8864 14414 8892 14991
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8446 14172 8754 14181
rect 8446 14170 8452 14172
rect 8508 14170 8532 14172
rect 8588 14170 8612 14172
rect 8668 14170 8692 14172
rect 8748 14170 8754 14172
rect 8508 14118 8510 14170
rect 8690 14118 8692 14170
rect 8446 14116 8452 14118
rect 8508 14116 8532 14118
rect 8588 14116 8612 14118
rect 8668 14116 8692 14118
rect 8748 14116 8754 14118
rect 8446 14107 8754 14116
rect 8446 13084 8754 13093
rect 8446 13082 8452 13084
rect 8508 13082 8532 13084
rect 8588 13082 8612 13084
rect 8668 13082 8692 13084
rect 8748 13082 8754 13084
rect 8508 13030 8510 13082
rect 8690 13030 8692 13082
rect 8446 13028 8452 13030
rect 8508 13028 8532 13030
rect 8588 13028 8612 13030
rect 8668 13028 8692 13030
rect 8748 13028 8754 13030
rect 8446 13019 8754 13028
rect 8864 12714 8892 14350
rect 8956 14278 8984 15302
rect 9048 14482 9076 15438
rect 9140 14482 9168 16118
rect 9232 14618 9260 16526
rect 9312 16516 9364 16522
rect 9312 16458 9364 16464
rect 9324 15042 9352 16458
rect 9416 16096 9444 17070
rect 9508 16454 9536 19200
rect 9680 17196 9732 17202
rect 9876 17184 9904 19200
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10046 17232 10102 17241
rect 9732 17156 9904 17184
rect 9956 17196 10008 17202
rect 9680 17138 9732 17144
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9600 16810 9628 16934
rect 9600 16782 9720 16810
rect 9588 16720 9640 16726
rect 9588 16662 9640 16668
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9496 16108 9548 16114
rect 9416 16068 9496 16096
rect 9496 16050 9548 16056
rect 9508 15910 9536 16050
rect 9600 16046 9628 16662
rect 9692 16590 9720 16782
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9416 15162 9444 15506
rect 9404 15156 9456 15162
rect 9404 15098 9456 15104
rect 9324 15014 9444 15042
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 9220 14612 9272 14618
rect 9220 14554 9272 14560
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8956 13938 8984 14214
rect 9048 14074 9076 14418
rect 9036 14068 9088 14074
rect 9036 14010 9088 14016
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 9140 13530 9168 14418
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9036 13456 9088 13462
rect 9036 13398 9088 13404
rect 9048 12866 9076 13398
rect 9140 12986 9168 13466
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9048 12838 9168 12866
rect 9324 12850 9352 14894
rect 9416 14482 9444 15014
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9416 13841 9444 14418
rect 9402 13832 9458 13841
rect 9402 13767 9458 13776
rect 8852 12708 8904 12714
rect 8852 12650 8904 12656
rect 9036 12640 9088 12646
rect 9036 12582 9088 12588
rect 9048 12434 9076 12582
rect 8864 12406 9076 12434
rect 8446 11996 8754 12005
rect 8446 11994 8452 11996
rect 8508 11994 8532 11996
rect 8588 11994 8612 11996
rect 8668 11994 8692 11996
rect 8748 11994 8754 11996
rect 8508 11942 8510 11994
rect 8690 11942 8692 11994
rect 8446 11940 8452 11942
rect 8508 11940 8532 11942
rect 8588 11940 8612 11942
rect 8668 11940 8692 11942
rect 8748 11940 8754 11942
rect 8446 11931 8754 11940
rect 8864 11082 8892 12406
rect 8852 11076 8904 11082
rect 8852 11018 8904 11024
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8446 10908 8754 10917
rect 8446 10906 8452 10908
rect 8508 10906 8532 10908
rect 8588 10906 8612 10908
rect 8668 10906 8692 10908
rect 8748 10906 8754 10908
rect 8508 10854 8510 10906
rect 8690 10854 8692 10906
rect 8446 10852 8452 10854
rect 8508 10852 8532 10854
rect 8588 10852 8612 10854
rect 8668 10852 8692 10854
rect 8748 10852 8754 10854
rect 8446 10843 8754 10852
rect 8956 10606 8984 10950
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8446 9820 8754 9829
rect 8446 9818 8452 9820
rect 8508 9818 8532 9820
rect 8588 9818 8612 9820
rect 8668 9818 8692 9820
rect 8748 9818 8754 9820
rect 8508 9766 8510 9818
rect 8690 9766 8692 9818
rect 8446 9764 8452 9766
rect 8508 9764 8532 9766
rect 8588 9764 8612 9766
rect 8668 9764 8692 9766
rect 8748 9764 8754 9766
rect 8446 9755 8754 9764
rect 8116 9648 8168 9654
rect 8116 9590 8168 9596
rect 8220 9646 8340 9674
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 8036 8838 8064 9318
rect 7932 8832 7984 8838
rect 7932 8774 7984 8780
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 7944 7818 7972 8774
rect 8036 8634 8064 8774
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7932 7812 7984 7818
rect 7932 7754 7984 7760
rect 7944 6458 7972 7754
rect 8128 7206 8156 9590
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7852 5846 7880 6326
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 7564 5840 7616 5846
rect 7564 5782 7616 5788
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 7840 5840 7892 5846
rect 7840 5782 7892 5788
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7484 5166 7512 5646
rect 7760 5556 7788 5782
rect 7576 5528 7788 5556
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7378 4856 7434 4865
rect 7378 4791 7434 4800
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 7300 4321 7328 4490
rect 7286 4312 7342 4321
rect 7286 4247 7342 4256
rect 7392 4214 7420 4791
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7116 4100 7236 4128
rect 7116 3641 7144 4100
rect 7288 4072 7340 4078
rect 7288 4014 7340 4020
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 6932 3590 7052 3618
rect 7102 3632 7158 3641
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6932 2922 6960 3590
rect 7102 3567 7158 3576
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 6920 2916 6972 2922
rect 6920 2858 6972 2864
rect 7024 2854 7052 3334
rect 7116 3194 7144 3470
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 7208 3058 7236 3946
rect 7300 3534 7328 4014
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 7104 2848 7156 2854
rect 7208 2825 7236 2858
rect 7104 2790 7156 2796
rect 7194 2816 7250 2825
rect 6572 2748 6880 2757
rect 6572 2746 6578 2748
rect 6634 2746 6658 2748
rect 6714 2746 6738 2748
rect 6794 2746 6818 2748
rect 6874 2746 6880 2748
rect 6634 2694 6636 2746
rect 6816 2694 6818 2746
rect 6572 2692 6578 2694
rect 6634 2692 6658 2694
rect 6714 2692 6738 2694
rect 6794 2692 6818 2694
rect 6874 2692 6880 2694
rect 6572 2683 6880 2692
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 5828 2038 5856 2382
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 6736 2304 6788 2310
rect 6736 2246 6788 2252
rect 5816 2032 5868 2038
rect 5816 1974 5868 1980
rect 5920 1170 5948 2246
rect 6288 1170 6316 2246
rect 6472 2106 6500 2246
rect 6460 2100 6512 2106
rect 6460 2042 6512 2048
rect 5920 1142 6040 1170
rect 6288 1142 6408 1170
rect 6012 800 6040 1142
rect 6380 800 6408 1142
rect 6748 800 6776 2246
rect 7116 800 7144 2790
rect 7194 2751 7250 2760
rect 7392 2446 7420 3878
rect 7484 3602 7512 5102
rect 7576 4146 7604 5528
rect 7746 5400 7802 5409
rect 7746 5335 7802 5344
rect 7760 5234 7788 5335
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7656 5160 7708 5166
rect 7852 5114 7880 5782
rect 7944 5710 7972 6258
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 8128 5846 8156 6054
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 7656 5102 7708 5108
rect 7668 4826 7696 5102
rect 7760 5086 7880 5114
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7484 2990 7512 3538
rect 7576 3398 7604 4082
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7668 3194 7696 4762
rect 7760 4690 7788 5086
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 7760 4282 7788 4422
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7760 3534 7788 4082
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7760 3058 7788 3470
rect 7852 3126 7880 4966
rect 7944 4078 7972 5646
rect 8022 5400 8078 5409
rect 8220 5386 8248 9646
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8446 8732 8754 8741
rect 8446 8730 8452 8732
rect 8508 8730 8532 8732
rect 8588 8730 8612 8732
rect 8668 8730 8692 8732
rect 8748 8730 8754 8732
rect 8508 8678 8510 8730
rect 8690 8678 8692 8730
rect 8446 8676 8452 8678
rect 8508 8676 8532 8678
rect 8588 8676 8612 8678
rect 8668 8676 8692 8678
rect 8748 8676 8754 8678
rect 8446 8667 8754 8676
rect 8864 8430 8892 8774
rect 8852 8424 8904 8430
rect 8852 8366 8904 8372
rect 8864 7886 8892 8366
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8446 7644 8754 7653
rect 8446 7642 8452 7644
rect 8508 7642 8532 7644
rect 8588 7642 8612 7644
rect 8668 7642 8692 7644
rect 8748 7642 8754 7644
rect 8508 7590 8510 7642
rect 8690 7590 8692 7642
rect 8446 7588 8452 7590
rect 8508 7588 8532 7590
rect 8588 7588 8612 7590
rect 8668 7588 8692 7590
rect 8748 7588 8754 7590
rect 8446 7579 8754 7588
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8404 7002 8432 7346
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8446 6556 8754 6565
rect 8446 6554 8452 6556
rect 8508 6554 8532 6556
rect 8588 6554 8612 6556
rect 8668 6554 8692 6556
rect 8748 6554 8754 6556
rect 8508 6502 8510 6554
rect 8690 6502 8692 6554
rect 8446 6500 8452 6502
rect 8508 6500 8532 6502
rect 8588 6500 8612 6502
rect 8668 6500 8692 6502
rect 8748 6500 8754 6502
rect 8446 6491 8754 6500
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8680 5914 8708 6190
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 8022 5335 8078 5344
rect 8128 5358 8248 5386
rect 8312 5370 8340 5850
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 8404 5574 8432 5714
rect 8772 5574 8800 6326
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8956 6118 8984 6258
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8446 5468 8754 5477
rect 8446 5466 8452 5468
rect 8508 5466 8532 5468
rect 8588 5466 8612 5468
rect 8668 5466 8692 5468
rect 8748 5466 8754 5468
rect 8508 5414 8510 5466
rect 8690 5414 8692 5466
rect 8446 5412 8452 5414
rect 8508 5412 8532 5414
rect 8588 5412 8612 5414
rect 8668 5412 8692 5414
rect 8748 5412 8754 5414
rect 8446 5403 8754 5412
rect 8300 5364 8352 5370
rect 8036 4570 8064 5335
rect 8128 4865 8156 5358
rect 8300 5306 8352 5312
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8114 4856 8170 4865
rect 8114 4791 8170 4800
rect 8036 4542 8156 4570
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7932 3392 7984 3398
rect 7930 3360 7932 3369
rect 7984 3360 7986 3369
rect 7930 3295 7986 3304
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7472 2984 7524 2990
rect 7760 2961 7788 2994
rect 7852 2990 7880 3062
rect 7840 2984 7892 2990
rect 7472 2926 7524 2932
rect 7746 2952 7802 2961
rect 7840 2926 7892 2932
rect 7746 2887 7802 2896
rect 8036 2582 8064 4422
rect 8128 3058 8156 4542
rect 8220 3942 8248 5170
rect 8956 4690 8984 6054
rect 9140 5953 9168 12838
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 9220 12164 9272 12170
rect 9220 12106 9272 12112
rect 9232 11558 9260 12106
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9232 11150 9260 11494
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9324 11014 9352 12650
rect 9508 12646 9536 15846
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9508 11898 9536 12174
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9496 11348 9548 11354
rect 9600 11336 9628 15982
rect 9692 15162 9720 16390
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 14657 9720 14758
rect 9678 14648 9734 14657
rect 9678 14583 9734 14592
rect 9784 14362 9812 17156
rect 10152 17202 10180 17614
rect 10046 17167 10102 17176
rect 10140 17196 10192 17202
rect 9956 17138 10008 17144
rect 9864 16176 9916 16182
rect 9968 16164 9996 17138
rect 10060 17134 10088 17167
rect 10140 17138 10192 17144
rect 10244 17134 10272 19200
rect 10612 17184 10640 19200
rect 10692 17196 10744 17202
rect 10612 17156 10692 17184
rect 10692 17138 10744 17144
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10152 16658 10180 16934
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 10060 16250 10088 16390
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 9916 16136 9996 16164
rect 10244 16130 10272 17070
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10320 16892 10628 16901
rect 10320 16890 10326 16892
rect 10382 16890 10406 16892
rect 10462 16890 10486 16892
rect 10542 16890 10566 16892
rect 10622 16890 10628 16892
rect 10382 16838 10384 16890
rect 10564 16838 10566 16890
rect 10320 16836 10326 16838
rect 10382 16836 10406 16838
rect 10462 16836 10486 16838
rect 10542 16836 10566 16838
rect 10622 16836 10628 16838
rect 10320 16827 10628 16836
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 9864 16118 9916 16124
rect 10060 16102 10272 16130
rect 9956 16040 10008 16046
rect 9954 16008 9956 16017
rect 10008 16008 10010 16017
rect 9954 15943 10010 15952
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9862 15736 9918 15745
rect 9862 15671 9918 15680
rect 9876 15502 9904 15671
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9968 15162 9996 15846
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9956 14884 10008 14890
rect 9956 14826 10008 14832
rect 9968 14482 9996 14826
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9692 14334 9812 14362
rect 9862 14376 9918 14385
rect 9692 13462 9720 14334
rect 9862 14311 9918 14320
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9784 13530 9812 14214
rect 9876 13920 9904 14311
rect 9956 14272 10008 14278
rect 9954 14240 9956 14249
rect 10008 14240 10010 14249
rect 9954 14175 10010 14184
rect 9956 13932 10008 13938
rect 9876 13892 9956 13920
rect 9956 13874 10008 13880
rect 9956 13796 10008 13802
rect 9956 13738 10008 13744
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9772 13524 9824 13530
rect 9772 13466 9824 13472
rect 9680 13456 9732 13462
rect 9680 13398 9732 13404
rect 9784 12918 9812 13466
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 9876 12730 9904 13670
rect 9548 11308 9628 11336
rect 9496 11290 9548 11296
rect 9600 11082 9628 11308
rect 9692 12702 9904 12730
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9692 10674 9720 12702
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9416 7698 9444 7822
rect 9600 7818 9628 9318
rect 9784 9178 9812 12582
rect 9968 11898 9996 13738
rect 10060 13190 10088 16102
rect 10336 15960 10364 16594
rect 10600 16584 10652 16590
rect 10600 16526 10652 16532
rect 10612 16182 10640 16526
rect 10704 16425 10732 16934
rect 10784 16720 10836 16726
rect 10784 16662 10836 16668
rect 10690 16416 10746 16425
rect 10690 16351 10746 16360
rect 10508 16176 10560 16182
rect 10508 16118 10560 16124
rect 10600 16176 10652 16182
rect 10600 16118 10652 16124
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10152 15932 10364 15960
rect 10152 15162 10180 15932
rect 10428 15892 10456 15982
rect 10520 15978 10548 16118
rect 10704 16017 10732 16351
rect 10690 16008 10746 16017
rect 10508 15972 10560 15978
rect 10690 15943 10746 15952
rect 10508 15914 10560 15920
rect 10244 15864 10456 15892
rect 10692 15904 10744 15910
rect 10244 15706 10272 15864
rect 10692 15846 10744 15852
rect 10320 15804 10628 15813
rect 10320 15802 10326 15804
rect 10382 15802 10406 15804
rect 10462 15802 10486 15804
rect 10542 15802 10566 15804
rect 10622 15802 10628 15804
rect 10382 15750 10384 15802
rect 10564 15750 10566 15802
rect 10320 15748 10326 15750
rect 10382 15748 10406 15750
rect 10462 15748 10486 15750
rect 10542 15748 10566 15750
rect 10622 15748 10628 15750
rect 10320 15739 10628 15748
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10508 15428 10560 15434
rect 10508 15370 10560 15376
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10140 15156 10192 15162
rect 10140 15098 10192 15104
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10152 13326 10180 14894
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 9968 11014 9996 11834
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9968 10810 9996 10950
rect 9956 10804 10008 10810
rect 10060 10792 10088 12922
rect 10152 11354 10180 13262
rect 10244 11762 10272 15302
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10428 14822 10456 15098
rect 10520 14822 10548 15370
rect 10416 14816 10468 14822
rect 10416 14758 10468 14764
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10320 14716 10628 14725
rect 10320 14714 10326 14716
rect 10382 14714 10406 14716
rect 10462 14714 10486 14716
rect 10542 14714 10566 14716
rect 10622 14714 10628 14716
rect 10382 14662 10384 14714
rect 10564 14662 10566 14714
rect 10320 14660 10326 14662
rect 10382 14660 10406 14662
rect 10462 14660 10486 14662
rect 10542 14660 10566 14662
rect 10622 14660 10628 14662
rect 10320 14651 10628 14660
rect 10704 14346 10732 15846
rect 10796 15434 10824 16662
rect 10784 15428 10836 15434
rect 10784 15370 10836 15376
rect 10782 15192 10838 15201
rect 10782 15127 10838 15136
rect 10796 14958 10824 15127
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10782 14784 10838 14793
rect 10782 14719 10838 14728
rect 10692 14340 10744 14346
rect 10692 14282 10744 14288
rect 10796 14278 10824 14719
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10320 13628 10628 13637
rect 10320 13626 10326 13628
rect 10382 13626 10406 13628
rect 10462 13626 10486 13628
rect 10542 13626 10566 13628
rect 10622 13626 10628 13628
rect 10382 13574 10384 13626
rect 10564 13574 10566 13626
rect 10320 13572 10326 13574
rect 10382 13572 10406 13574
rect 10462 13572 10486 13574
rect 10542 13572 10566 13574
rect 10622 13572 10628 13574
rect 10320 13563 10628 13572
rect 10598 13016 10654 13025
rect 10598 12951 10600 12960
rect 10652 12951 10654 12960
rect 10600 12922 10652 12928
rect 10320 12540 10628 12549
rect 10320 12538 10326 12540
rect 10382 12538 10406 12540
rect 10462 12538 10486 12540
rect 10542 12538 10566 12540
rect 10622 12538 10628 12540
rect 10382 12486 10384 12538
rect 10564 12486 10566 12538
rect 10320 12484 10326 12486
rect 10382 12484 10406 12486
rect 10462 12484 10486 12486
rect 10542 12484 10566 12486
rect 10622 12484 10628 12486
rect 10320 12475 10628 12484
rect 10232 11756 10284 11762
rect 10232 11698 10284 11704
rect 10320 11452 10628 11461
rect 10320 11450 10326 11452
rect 10382 11450 10406 11452
rect 10462 11450 10486 11452
rect 10542 11450 10566 11452
rect 10622 11450 10628 11452
rect 10382 11398 10384 11450
rect 10564 11398 10566 11450
rect 10320 11396 10326 11398
rect 10382 11396 10406 11398
rect 10462 11396 10486 11398
rect 10542 11396 10566 11398
rect 10622 11396 10628 11398
rect 10320 11387 10628 11396
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10704 10810 10732 14010
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10796 12986 10824 13126
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10796 12714 10824 12922
rect 10784 12708 10836 12714
rect 10784 12650 10836 12656
rect 10782 12608 10838 12617
rect 10782 12543 10838 12552
rect 10692 10804 10744 10810
rect 10060 10764 10272 10792
rect 9956 10746 10008 10752
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 10060 9178 10088 10610
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9416 7670 9628 7698
rect 9600 7410 9628 7670
rect 9312 7404 9364 7410
rect 9588 7404 9640 7410
rect 9364 7364 9444 7392
rect 9312 7346 9364 7352
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9126 5944 9182 5953
rect 9126 5879 9182 5888
rect 9140 5574 9168 5879
rect 9218 5808 9274 5817
rect 9324 5778 9352 6258
rect 9218 5743 9274 5752
rect 9312 5772 9364 5778
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9232 4826 9260 5743
rect 9312 5714 9364 5720
rect 9312 5636 9364 5642
rect 9312 5578 9364 5584
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8312 4282 8340 4422
rect 8446 4380 8754 4389
rect 8446 4378 8452 4380
rect 8508 4378 8532 4380
rect 8588 4378 8612 4380
rect 8668 4378 8692 4380
rect 8748 4378 8754 4380
rect 8508 4326 8510 4378
rect 8690 4326 8692 4378
rect 8446 4324 8452 4326
rect 8508 4324 8532 4326
rect 8588 4324 8612 4326
rect 8668 4324 8692 4326
rect 8748 4324 8754 4326
rect 8446 4315 8754 4324
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8220 3058 8248 3878
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 7840 2576 7892 2582
rect 7840 2518 7892 2524
rect 8024 2576 8076 2582
rect 8024 2518 8076 2524
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 7484 800 7512 2246
rect 7852 800 7880 2518
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 7944 2106 7972 2382
rect 7932 2100 7984 2106
rect 7932 2042 7984 2048
rect 8220 800 8248 2586
rect 8312 2514 8340 4082
rect 8772 3466 8800 4082
rect 8760 3460 8812 3466
rect 8760 3402 8812 3408
rect 8446 3292 8754 3301
rect 8446 3290 8452 3292
rect 8508 3290 8532 3292
rect 8588 3290 8612 3292
rect 8668 3290 8692 3292
rect 8748 3290 8754 3292
rect 8508 3238 8510 3290
rect 8690 3238 8692 3290
rect 8446 3236 8452 3238
rect 8508 3236 8532 3238
rect 8588 3236 8612 3238
rect 8668 3236 8692 3238
rect 8748 3236 8754 3238
rect 8446 3227 8754 3236
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 8404 2446 8432 2858
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8496 2514 8524 2790
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8446 2204 8754 2213
rect 8446 2202 8452 2204
rect 8508 2202 8532 2204
rect 8588 2202 8612 2204
rect 8668 2202 8692 2204
rect 8748 2202 8754 2204
rect 8508 2150 8510 2202
rect 8690 2150 8692 2202
rect 8446 2148 8452 2150
rect 8508 2148 8532 2150
rect 8588 2148 8612 2150
rect 8668 2148 8692 2150
rect 8748 2148 8754 2150
rect 8446 2139 8754 2148
rect 8588 870 8708 898
rect 8588 800 8616 870
rect 1214 0 1270 800
rect 1582 0 1638 800
rect 1950 0 2006 800
rect 2318 0 2374 800
rect 2686 0 2742 800
rect 3054 0 3110 800
rect 3422 0 3478 800
rect 3790 0 3846 800
rect 4158 0 4214 800
rect 4526 0 4582 800
rect 4894 0 4950 800
rect 5262 0 5318 800
rect 5630 0 5686 800
rect 5998 0 6054 800
rect 6366 0 6422 800
rect 6734 0 6790 800
rect 7102 0 7158 800
rect 7470 0 7526 800
rect 7838 0 7894 800
rect 8206 0 8262 800
rect 8574 0 8630 800
rect 8680 762 8708 870
rect 8864 762 8892 4490
rect 8956 3602 8984 4626
rect 9232 4146 9260 4762
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9048 3670 9076 3878
rect 9036 3664 9088 3670
rect 9036 3606 9088 3612
rect 8944 3596 8996 3602
rect 9232 3584 9260 4082
rect 8944 3538 8996 3544
rect 9201 3556 9260 3584
rect 9201 3516 9229 3556
rect 9324 3534 9352 5578
rect 9416 5098 9444 7364
rect 9588 7346 9640 7352
rect 9600 7002 9628 7346
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 9600 5914 9628 6938
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9600 5778 9628 5850
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 9404 4752 9456 4758
rect 9404 4694 9456 4700
rect 9588 4752 9640 4758
rect 9588 4694 9640 4700
rect 9416 4282 9444 4694
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9600 4214 9628 4694
rect 9692 4690 9720 6598
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9784 5642 9812 6054
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 9772 5636 9824 5642
rect 9772 5578 9824 5584
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9402 3768 9458 3777
rect 9508 3738 9536 4082
rect 9402 3703 9458 3712
rect 9496 3732 9548 3738
rect 9048 3488 9229 3516
rect 9312 3528 9364 3534
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8956 3194 8984 3334
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9048 2650 9076 3488
rect 9312 3470 9364 3476
rect 9416 3482 9444 3703
rect 9496 3674 9548 3680
rect 9692 3602 9720 4082
rect 9784 4078 9812 5578
rect 9876 5030 9904 5646
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9876 4865 9904 4966
rect 9862 4856 9918 4865
rect 9862 4791 9918 4800
rect 9968 4604 9996 6394
rect 10152 5409 10180 9590
rect 10138 5400 10194 5409
rect 10048 5364 10100 5370
rect 10244 5370 10272 10764
rect 10692 10746 10744 10752
rect 10796 10554 10824 12543
rect 10888 12442 10916 17138
rect 10980 16590 11008 19200
rect 11150 17096 11206 17105
rect 11060 17060 11112 17066
rect 11150 17031 11206 17040
rect 11060 17002 11112 17008
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10980 15502 11008 16390
rect 11072 15706 11100 17002
rect 11164 16697 11192 17031
rect 11150 16688 11206 16697
rect 11150 16623 11206 16632
rect 11244 16516 11296 16522
rect 11348 16504 11376 19200
rect 11716 17202 11744 19200
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11296 16476 11376 16504
rect 11244 16458 11296 16464
rect 11150 16144 11206 16153
rect 11150 16079 11206 16088
rect 11336 16108 11388 16114
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 11060 15496 11112 15502
rect 11060 15438 11112 15444
rect 10968 15088 11020 15094
rect 10966 15056 10968 15065
rect 11020 15056 11022 15065
rect 10966 14991 11022 15000
rect 10966 14104 11022 14113
rect 10966 14039 11022 14048
rect 10980 14006 11008 14039
rect 10968 14000 11020 14006
rect 10968 13942 11020 13948
rect 10980 13190 11008 13942
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10968 12912 11020 12918
rect 10968 12854 11020 12860
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10980 12322 11008 12854
rect 11072 12374 11100 15438
rect 11164 15366 11192 16079
rect 11336 16050 11388 16056
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11150 15192 11206 15201
rect 11150 15127 11206 15136
rect 11164 13462 11192 15127
rect 11256 15026 11284 15846
rect 11348 15162 11376 16050
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11440 14618 11468 15302
rect 11428 14612 11480 14618
rect 11428 14554 11480 14560
rect 11532 14550 11560 16526
rect 11624 16250 11652 16730
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 11520 14544 11572 14550
rect 11520 14486 11572 14492
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11152 13456 11204 13462
rect 11152 13398 11204 13404
rect 11164 12986 11192 13398
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 10888 12294 11008 12322
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 10888 12238 10916 12294
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10888 11694 10916 12174
rect 11256 12102 11284 14418
rect 11428 13796 11480 13802
rect 11428 13738 11480 13744
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11348 12238 11376 13670
rect 11440 12782 11468 13738
rect 11624 13530 11652 14894
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11624 13326 11652 13466
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11624 12850 11652 13262
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11428 12776 11480 12782
rect 11426 12744 11428 12753
rect 11480 12744 11482 12753
rect 11426 12679 11482 12688
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11256 11830 11284 12038
rect 11348 11898 11376 12038
rect 11716 11898 11744 17138
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11808 16697 11836 17070
rect 11794 16688 11850 16697
rect 11794 16623 11850 16632
rect 12084 16590 12112 19200
rect 12452 17524 12480 19200
rect 12452 17496 12572 17524
rect 12194 17436 12502 17445
rect 12194 17434 12200 17436
rect 12256 17434 12280 17436
rect 12336 17434 12360 17436
rect 12416 17434 12440 17436
rect 12496 17434 12502 17436
rect 12256 17382 12258 17434
rect 12438 17382 12440 17434
rect 12194 17380 12200 17382
rect 12256 17380 12280 17382
rect 12336 17380 12360 17382
rect 12416 17380 12440 17382
rect 12496 17380 12502 17382
rect 12194 17371 12502 17380
rect 12544 17202 12572 17496
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12728 16969 12756 17070
rect 12714 16960 12770 16969
rect 12714 16895 12770 16904
rect 12714 16688 12770 16697
rect 12714 16623 12716 16632
rect 12768 16623 12770 16632
rect 12716 16594 12768 16600
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 12194 16348 12502 16357
rect 12194 16346 12200 16348
rect 12256 16346 12280 16348
rect 12336 16346 12360 16348
rect 12416 16346 12440 16348
rect 12496 16346 12502 16348
rect 12256 16294 12258 16346
rect 12438 16294 12440 16346
rect 12194 16292 12200 16294
rect 12256 16292 12280 16294
rect 12336 16292 12360 16294
rect 12416 16292 12440 16294
rect 12496 16292 12502 16294
rect 12194 16283 12502 16292
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 12084 15570 12112 16186
rect 12820 16182 12848 19200
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 12808 16176 12860 16182
rect 12808 16118 12860 16124
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12532 15972 12584 15978
rect 12532 15914 12584 15920
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 12360 15638 12388 15846
rect 12348 15632 12400 15638
rect 12348 15574 12400 15580
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 11808 15201 11836 15506
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11794 15192 11850 15201
rect 11794 15127 11850 15136
rect 11796 15088 11848 15094
rect 11796 15030 11848 15036
rect 11808 14958 11836 15030
rect 11796 14952 11848 14958
rect 11794 14920 11796 14929
rect 11848 14920 11850 14929
rect 11794 14855 11850 14864
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11808 13734 11836 14214
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11808 12170 11836 13670
rect 11900 13512 11928 15438
rect 11980 15428 12032 15434
rect 11980 15370 12032 15376
rect 11992 14890 12020 15370
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 12084 15162 12112 15302
rect 12194 15260 12502 15269
rect 12194 15258 12200 15260
rect 12256 15258 12280 15260
rect 12336 15258 12360 15260
rect 12416 15258 12440 15260
rect 12496 15258 12502 15260
rect 12256 15206 12258 15258
rect 12438 15206 12440 15258
rect 12194 15204 12200 15206
rect 12256 15204 12280 15206
rect 12336 15204 12360 15206
rect 12416 15204 12440 15206
rect 12496 15204 12502 15206
rect 12194 15195 12502 15204
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11992 14278 12020 14486
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11980 13524 12032 13530
rect 11900 13484 11980 13512
rect 11980 13466 12032 13472
rect 12084 13190 12112 14894
rect 12452 14822 12480 14962
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12452 14618 12480 14758
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12544 14414 12572 15914
rect 12636 15706 12664 15982
rect 13004 15722 13032 16050
rect 12624 15700 12676 15706
rect 12624 15642 12676 15648
rect 12820 15694 13032 15722
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12194 14172 12502 14181
rect 12194 14170 12200 14172
rect 12256 14170 12280 14172
rect 12336 14170 12360 14172
rect 12416 14170 12440 14172
rect 12496 14170 12502 14172
rect 12256 14118 12258 14170
rect 12438 14118 12440 14170
rect 12194 14116 12200 14118
rect 12256 14116 12280 14118
rect 12336 14116 12360 14118
rect 12416 14116 12440 14118
rect 12496 14116 12502 14118
rect 12194 14107 12502 14116
rect 12636 13258 12664 14894
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 12194 13084 12502 13093
rect 12194 13082 12200 13084
rect 12256 13082 12280 13084
rect 12336 13082 12360 13084
rect 12416 13082 12440 13084
rect 12496 13082 12502 13084
rect 12256 13030 12258 13082
rect 12438 13030 12440 13082
rect 12194 13028 12200 13030
rect 12256 13028 12280 13030
rect 12336 13028 12360 13030
rect 12416 13028 12440 13030
rect 12496 13028 12502 13030
rect 12194 13019 12502 13028
rect 12728 12986 12756 15438
rect 12820 15366 12848 15694
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12808 15360 12860 15366
rect 12806 15328 12808 15337
rect 12860 15328 12862 15337
rect 12806 15263 12862 15272
rect 12912 15178 12940 15506
rect 12820 15150 12940 15178
rect 12820 13938 12848 15150
rect 12992 14952 13044 14958
rect 12912 14900 12992 14906
rect 12912 14894 13044 14900
rect 12912 14878 13032 14894
rect 12912 14346 12940 14878
rect 13096 14770 13124 17138
rect 13188 17134 13216 19200
rect 13556 17898 13584 19200
rect 13556 17870 13676 17898
rect 13544 17740 13596 17746
rect 13544 17682 13596 17688
rect 13452 17604 13504 17610
rect 13452 17546 13504 17552
rect 13464 17338 13492 17546
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13450 17096 13506 17105
rect 13450 17031 13506 17040
rect 13358 16824 13414 16833
rect 13358 16759 13414 16768
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 13176 15972 13228 15978
rect 13176 15914 13228 15920
rect 13004 14742 13124 14770
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12912 13734 12940 14282
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12820 13258 12848 13466
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12360 12170 12388 12922
rect 12728 12889 12756 12922
rect 12714 12880 12770 12889
rect 12714 12815 12770 12824
rect 12912 12782 12940 13670
rect 12900 12776 12952 12782
rect 12900 12718 12952 12724
rect 12900 12368 12952 12374
rect 12900 12310 12952 12316
rect 11796 12164 11848 12170
rect 11796 12106 11848 12112
rect 12348 12164 12400 12170
rect 12348 12106 12400 12112
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12194 11996 12502 12005
rect 12194 11994 12200 11996
rect 12256 11994 12280 11996
rect 12336 11994 12360 11996
rect 12416 11994 12440 11996
rect 12496 11994 12502 11996
rect 12256 11942 12258 11994
rect 12438 11942 12440 11994
rect 12194 11940 12200 11942
rect 12256 11940 12280 11942
rect 12336 11940 12360 11942
rect 12416 11940 12440 11942
rect 12496 11940 12502 11942
rect 12194 11931 12502 11940
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11244 11824 11296 11830
rect 11244 11766 11296 11772
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 12072 11688 12124 11694
rect 12072 11630 12124 11636
rect 10888 11354 10916 11630
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 11072 10742 11100 11494
rect 12084 11014 12112 11630
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 11060 10736 11112 10742
rect 11060 10678 11112 10684
rect 11900 10606 11928 10950
rect 10704 10526 10824 10554
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 10320 10364 10628 10373
rect 10320 10362 10326 10364
rect 10382 10362 10406 10364
rect 10462 10362 10486 10364
rect 10542 10362 10566 10364
rect 10622 10362 10628 10364
rect 10382 10310 10384 10362
rect 10564 10310 10566 10362
rect 10320 10308 10326 10310
rect 10382 10308 10406 10310
rect 10462 10308 10486 10310
rect 10542 10308 10566 10310
rect 10622 10308 10628 10310
rect 10320 10299 10628 10308
rect 10320 9276 10628 9285
rect 10320 9274 10326 9276
rect 10382 9274 10406 9276
rect 10462 9274 10486 9276
rect 10542 9274 10566 9276
rect 10622 9274 10628 9276
rect 10382 9222 10384 9274
rect 10564 9222 10566 9274
rect 10320 9220 10326 9222
rect 10382 9220 10406 9222
rect 10462 9220 10486 9222
rect 10542 9220 10566 9222
rect 10622 9220 10628 9222
rect 10320 9211 10628 9220
rect 10320 8188 10628 8197
rect 10320 8186 10326 8188
rect 10382 8186 10406 8188
rect 10462 8186 10486 8188
rect 10542 8186 10566 8188
rect 10622 8186 10628 8188
rect 10382 8134 10384 8186
rect 10564 8134 10566 8186
rect 10320 8132 10326 8134
rect 10382 8132 10406 8134
rect 10462 8132 10486 8134
rect 10542 8132 10566 8134
rect 10622 8132 10628 8134
rect 10320 8123 10628 8132
rect 10320 7100 10628 7109
rect 10320 7098 10326 7100
rect 10382 7098 10406 7100
rect 10462 7098 10486 7100
rect 10542 7098 10566 7100
rect 10622 7098 10628 7100
rect 10382 7046 10384 7098
rect 10564 7046 10566 7098
rect 10320 7044 10326 7046
rect 10382 7044 10406 7046
rect 10462 7044 10486 7046
rect 10542 7044 10566 7046
rect 10622 7044 10628 7046
rect 10320 7035 10628 7044
rect 10320 6012 10628 6021
rect 10320 6010 10326 6012
rect 10382 6010 10406 6012
rect 10462 6010 10486 6012
rect 10542 6010 10566 6012
rect 10622 6010 10628 6012
rect 10382 5958 10384 6010
rect 10564 5958 10566 6010
rect 10320 5956 10326 5958
rect 10382 5956 10406 5958
rect 10462 5956 10486 5958
rect 10542 5956 10566 5958
rect 10622 5956 10628 5958
rect 10320 5947 10628 5956
rect 10704 5914 10732 10526
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10796 10266 10824 10406
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11164 9722 11192 10066
rect 12084 9994 12112 10950
rect 12194 10908 12502 10917
rect 12194 10906 12200 10908
rect 12256 10906 12280 10908
rect 12336 10906 12360 10908
rect 12416 10906 12440 10908
rect 12496 10906 12502 10908
rect 12256 10854 12258 10906
rect 12438 10854 12440 10906
rect 12194 10852 12200 10854
rect 12256 10852 12280 10854
rect 12336 10852 12360 10854
rect 12416 10852 12440 10854
rect 12496 10852 12502 10854
rect 12194 10843 12502 10852
rect 12544 10810 12572 11290
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11624 8974 11652 9862
rect 12194 9820 12502 9829
rect 12194 9818 12200 9820
rect 12256 9818 12280 9820
rect 12336 9818 12360 9820
rect 12416 9818 12440 9820
rect 12496 9818 12502 9820
rect 12256 9766 12258 9818
rect 12438 9766 12440 9818
rect 12194 9764 12200 9766
rect 12256 9764 12280 9766
rect 12336 9764 12360 9766
rect 12416 9764 12440 9766
rect 12496 9764 12502 9766
rect 12194 9755 12502 9764
rect 12544 9654 12572 10746
rect 12636 10538 12664 11698
rect 12728 10538 12756 11698
rect 12820 10742 12848 12038
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12716 10532 12768 10538
rect 12716 10474 12768 10480
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12820 9110 12848 9522
rect 12808 9104 12860 9110
rect 12714 9072 12770 9081
rect 12808 9046 12860 9052
rect 12714 9007 12770 9016
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 12728 8906 12756 9007
rect 11888 8900 11940 8906
rect 11888 8842 11940 8848
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10796 7886 10824 8230
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10796 7478 10824 7822
rect 11624 7478 11652 8298
rect 11900 8090 11928 8842
rect 12194 8732 12502 8741
rect 12194 8730 12200 8732
rect 12256 8730 12280 8732
rect 12336 8730 12360 8732
rect 12416 8730 12440 8732
rect 12496 8730 12502 8732
rect 12256 8678 12258 8730
rect 12438 8678 12440 8730
rect 12194 8676 12200 8678
rect 12256 8676 12280 8678
rect 12336 8676 12360 8678
rect 12416 8676 12440 8678
rect 12496 8676 12502 8678
rect 12194 8667 12502 8676
rect 12728 8294 12756 8842
rect 12912 8378 12940 12310
rect 13004 11898 13032 14742
rect 13188 14385 13216 15914
rect 13174 14376 13230 14385
rect 13084 14340 13136 14346
rect 13174 14311 13230 14320
rect 13084 14282 13136 14288
rect 13096 14006 13124 14282
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 13096 13530 13124 13942
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 13096 12918 13124 13466
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 13096 12306 13124 12854
rect 13188 12646 13216 13806
rect 13280 12986 13308 16594
rect 13372 14618 13400 16759
rect 13464 16697 13492 17031
rect 13450 16688 13506 16697
rect 13450 16623 13452 16632
rect 13504 16623 13506 16632
rect 13452 16594 13504 16600
rect 13556 16250 13584 17682
rect 13648 16794 13676 17870
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13636 16788 13688 16794
rect 13636 16730 13688 16736
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13452 16176 13504 16182
rect 13452 16118 13504 16124
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13372 13530 13400 13874
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 13084 12300 13136 12306
rect 13084 12242 13136 12248
rect 13174 11928 13230 11937
rect 12992 11892 13044 11898
rect 13174 11863 13176 11872
rect 12992 11834 13044 11840
rect 13228 11863 13230 11872
rect 13176 11834 13228 11840
rect 13372 11642 13400 13194
rect 13464 12306 13492 16118
rect 13648 15450 13676 16730
rect 13832 16658 13860 16934
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13832 15473 13860 15982
rect 13818 15464 13874 15473
rect 13544 15428 13596 15434
rect 13648 15422 13768 15450
rect 13544 15370 13596 15376
rect 13556 15042 13584 15370
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13648 15162 13676 15302
rect 13636 15156 13688 15162
rect 13636 15098 13688 15104
rect 13740 15065 13768 15422
rect 13924 15450 13952 19200
rect 14292 19122 14320 19200
rect 14384 19122 14412 19230
rect 14292 19094 14412 19122
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14372 17128 14424 17134
rect 14370 17096 14372 17105
rect 14424 17096 14426 17105
rect 14370 17031 14426 17040
rect 14068 16892 14376 16901
rect 14068 16890 14074 16892
rect 14130 16890 14154 16892
rect 14210 16890 14234 16892
rect 14290 16890 14314 16892
rect 14370 16890 14376 16892
rect 14130 16838 14132 16890
rect 14312 16838 14314 16890
rect 14068 16836 14074 16838
rect 14130 16836 14154 16838
rect 14210 16836 14234 16838
rect 14290 16836 14314 16838
rect 14370 16836 14376 16838
rect 14068 16827 14376 16836
rect 14476 16250 14504 17138
rect 14464 16244 14516 16250
rect 14464 16186 14516 16192
rect 14068 15804 14376 15813
rect 14068 15802 14074 15804
rect 14130 15802 14154 15804
rect 14210 15802 14234 15804
rect 14290 15802 14314 15804
rect 14370 15802 14376 15804
rect 14130 15750 14132 15802
rect 14312 15750 14314 15802
rect 14068 15748 14074 15750
rect 14130 15748 14154 15750
rect 14210 15748 14234 15750
rect 14290 15748 14314 15750
rect 14370 15748 14376 15750
rect 14068 15739 14376 15748
rect 14280 15564 14332 15570
rect 14280 15506 14332 15512
rect 13924 15434 14044 15450
rect 13924 15428 14056 15434
rect 13924 15422 14004 15428
rect 13818 15399 13874 15408
rect 14004 15370 14056 15376
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 13726 15056 13782 15065
rect 13556 15014 13676 15042
rect 13542 14920 13598 14929
rect 13542 14855 13598 14864
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13556 11830 13584 14855
rect 13648 14414 13676 15014
rect 13726 14991 13782 15000
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13636 14408 13688 14414
rect 13636 14350 13688 14356
rect 13544 11824 13596 11830
rect 13544 11766 13596 11772
rect 13372 11614 13492 11642
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13372 10810 13400 11494
rect 13360 10804 13412 10810
rect 13360 10746 13412 10752
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13096 9722 13124 9862
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13174 8936 13230 8945
rect 13174 8871 13230 8880
rect 13188 8838 13216 8871
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 12820 8350 12940 8378
rect 13188 8362 13216 8774
rect 13176 8356 13228 8362
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 11702 7848 11758 7857
rect 12636 7818 12664 7958
rect 11702 7783 11758 7792
rect 12624 7812 12676 7818
rect 10784 7472 10836 7478
rect 10784 7414 10836 7420
rect 11612 7472 11664 7478
rect 11612 7414 11664 7420
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 10968 6384 11020 6390
rect 10966 6352 10968 6361
rect 11020 6352 11022 6361
rect 10966 6287 11022 6296
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 11164 5846 11192 7346
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11348 6730 11376 7142
rect 11426 6760 11482 6769
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 11336 6724 11388 6730
rect 11426 6695 11482 6704
rect 11336 6666 11388 6672
rect 11256 5914 11284 6666
rect 11244 5908 11296 5914
rect 11244 5850 11296 5856
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 11164 5574 11192 5782
rect 10324 5568 10376 5574
rect 10322 5536 10324 5545
rect 10968 5568 11020 5574
rect 10376 5536 10378 5545
rect 10968 5510 11020 5516
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 10322 5471 10378 5480
rect 10138 5335 10194 5344
rect 10232 5364 10284 5370
rect 10048 5306 10100 5312
rect 10232 5306 10284 5312
rect 10784 5364 10836 5370
rect 10784 5306 10836 5312
rect 9876 4576 9996 4604
rect 9876 4146 9904 4576
rect 9956 4480 10008 4486
rect 9956 4422 10008 4428
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9862 4040 9918 4049
rect 9862 3975 9864 3984
rect 9916 3975 9918 3984
rect 9864 3946 9916 3952
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9416 3454 9536 3482
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9324 3194 9352 3334
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8956 800 8984 2246
rect 9324 800 9352 2994
rect 9416 2922 9444 3334
rect 9404 2916 9456 2922
rect 9404 2858 9456 2864
rect 9508 2582 9536 3454
rect 9588 3460 9640 3466
rect 9588 3402 9640 3408
rect 9600 3058 9628 3402
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9692 2774 9720 2926
rect 9600 2746 9720 2774
rect 9496 2576 9548 2582
rect 9496 2518 9548 2524
rect 9600 2514 9628 2746
rect 9784 2650 9812 3878
rect 9968 3738 9996 4422
rect 10060 4185 10088 5306
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 10046 4176 10102 4185
rect 10046 4111 10102 4120
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 10152 3534 10180 5238
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 10244 4826 10272 5034
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10320 4924 10628 4933
rect 10320 4922 10326 4924
rect 10382 4922 10406 4924
rect 10462 4922 10486 4924
rect 10542 4922 10566 4924
rect 10622 4922 10628 4924
rect 10382 4870 10384 4922
rect 10564 4870 10566 4922
rect 10320 4868 10326 4870
rect 10382 4868 10406 4870
rect 10462 4868 10486 4870
rect 10542 4868 10566 4870
rect 10622 4868 10628 4870
rect 10320 4859 10628 4868
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10244 4214 10272 4558
rect 10324 4548 10376 4554
rect 10324 4490 10376 4496
rect 10336 4282 10364 4490
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10232 4208 10284 4214
rect 10232 4150 10284 4156
rect 10428 3924 10456 4762
rect 10506 4584 10562 4593
rect 10506 4519 10562 4528
rect 10520 4010 10548 4519
rect 10508 4004 10560 4010
rect 10508 3946 10560 3952
rect 10244 3896 10456 3924
rect 10140 3528 10192 3534
rect 10244 3505 10272 3896
rect 10320 3836 10628 3845
rect 10320 3834 10326 3836
rect 10382 3834 10406 3836
rect 10462 3834 10486 3836
rect 10542 3834 10566 3836
rect 10622 3834 10628 3836
rect 10382 3782 10384 3834
rect 10564 3782 10566 3834
rect 10320 3780 10326 3782
rect 10382 3780 10406 3782
rect 10462 3780 10486 3782
rect 10542 3780 10566 3782
rect 10622 3780 10628 3782
rect 10320 3771 10628 3780
rect 10600 3596 10652 3602
rect 10600 3538 10652 3544
rect 10140 3470 10192 3476
rect 10230 3496 10286 3505
rect 10230 3431 10286 3440
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 9954 3224 10010 3233
rect 10060 3194 10088 3334
rect 9954 3159 10010 3168
rect 10048 3188 10100 3194
rect 9864 3052 9916 3058
rect 9864 2994 9916 3000
rect 9876 2825 9904 2994
rect 9968 2990 9996 3159
rect 10048 3130 10100 3136
rect 10244 3126 10272 3431
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 10322 3088 10378 3097
rect 10322 3023 10378 3032
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 10336 2904 10364 3023
rect 10612 2922 10640 3538
rect 10244 2876 10364 2904
rect 10600 2916 10652 2922
rect 9862 2816 9918 2825
rect 9862 2751 9918 2760
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 9692 2038 9720 2314
rect 9876 2038 9904 2450
rect 10244 2310 10272 2876
rect 10600 2858 10652 2864
rect 10320 2748 10628 2757
rect 10320 2746 10326 2748
rect 10382 2746 10406 2748
rect 10462 2746 10486 2748
rect 10542 2746 10566 2748
rect 10622 2746 10628 2748
rect 10382 2694 10384 2746
rect 10564 2694 10566 2746
rect 10320 2692 10326 2694
rect 10382 2692 10406 2694
rect 10462 2692 10486 2694
rect 10542 2692 10566 2694
rect 10622 2692 10628 2694
rect 10320 2683 10628 2692
rect 10336 2514 10548 2530
rect 10324 2508 10548 2514
rect 10376 2502 10548 2508
rect 10324 2450 10376 2456
rect 10520 2394 10548 2502
rect 10704 2446 10732 4966
rect 10796 4826 10824 5306
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10796 3738 10824 4014
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10888 3126 10916 4966
rect 10980 4826 11008 5510
rect 11256 5166 11284 5850
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 11348 4758 11376 6666
rect 11440 6458 11468 6695
rect 11532 6458 11560 7278
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11716 6390 11744 7783
rect 12624 7754 12676 7760
rect 12194 7644 12502 7653
rect 12194 7642 12200 7644
rect 12256 7642 12280 7644
rect 12336 7642 12360 7644
rect 12416 7642 12440 7644
rect 12496 7642 12502 7644
rect 12256 7590 12258 7642
rect 12438 7590 12440 7642
rect 12194 7588 12200 7590
rect 12256 7588 12280 7590
rect 12336 7588 12360 7590
rect 12416 7588 12440 7590
rect 12496 7588 12502 7590
rect 12194 7579 12502 7588
rect 12728 7562 12756 8230
rect 12636 7534 12756 7562
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 11704 6384 11756 6390
rect 11704 6326 11756 6332
rect 11716 6202 11744 6326
rect 11532 6174 11744 6202
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11532 5352 11560 6174
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11440 5324 11560 5352
rect 11440 5166 11468 5324
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 10980 3534 11008 4558
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11150 4448 11206 4457
rect 11072 4282 11100 4422
rect 11348 4434 11376 4694
rect 11206 4406 11376 4434
rect 11150 4383 11206 4392
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 11164 4146 11192 4383
rect 11242 4312 11298 4321
rect 11242 4247 11298 4256
rect 11256 4214 11284 4247
rect 11244 4208 11296 4214
rect 11244 4150 11296 4156
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10876 3120 10928 3126
rect 10796 3080 10876 3108
rect 10692 2440 10744 2446
rect 10520 2378 10640 2394
rect 10692 2382 10744 2388
rect 10416 2372 10468 2378
rect 10520 2372 10652 2378
rect 10520 2366 10600 2372
rect 10416 2314 10468 2320
rect 10600 2314 10652 2320
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 9680 2032 9732 2038
rect 9680 1974 9732 1980
rect 9864 2032 9916 2038
rect 9864 1974 9916 1980
rect 9692 800 9720 1974
rect 10048 1556 10100 1562
rect 10048 1498 10100 1504
rect 10060 800 10088 1498
rect 10428 800 10456 2314
rect 10796 800 10824 3080
rect 10876 3062 10928 3068
rect 10980 2650 11008 3334
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 11072 1970 11100 3946
rect 11242 3768 11298 3777
rect 11242 3703 11298 3712
rect 11256 3602 11284 3703
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 11060 1964 11112 1970
rect 11060 1906 11112 1912
rect 11164 800 11192 3402
rect 11256 2378 11284 3402
rect 11334 3224 11390 3233
rect 11334 3159 11336 3168
rect 11388 3159 11390 3168
rect 11336 3130 11388 3136
rect 11440 3126 11468 5102
rect 11532 4826 11560 5170
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 11532 4282 11560 4422
rect 11520 4276 11572 4282
rect 11520 4218 11572 4224
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11428 3120 11480 3126
rect 11428 3062 11480 3068
rect 11440 2446 11468 3062
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 11244 2372 11296 2378
rect 11244 2314 11296 2320
rect 11532 800 11560 4082
rect 11624 2938 11652 6054
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11716 4078 11744 5510
rect 11808 4214 11836 5578
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11704 4072 11756 4078
rect 11756 4032 11836 4060
rect 11704 4014 11756 4020
rect 11624 2910 11744 2938
rect 11612 2848 11664 2854
rect 11612 2790 11664 2796
rect 11624 2038 11652 2790
rect 11716 2446 11744 2910
rect 11808 2854 11836 4032
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11900 2774 11928 6190
rect 11992 5574 12020 6598
rect 12084 6458 12112 6734
rect 12194 6556 12502 6565
rect 12194 6554 12200 6556
rect 12256 6554 12280 6556
rect 12336 6554 12360 6556
rect 12416 6554 12440 6556
rect 12496 6554 12502 6556
rect 12256 6502 12258 6554
rect 12438 6502 12440 6554
rect 12194 6500 12200 6502
rect 12256 6500 12280 6502
rect 12336 6500 12360 6502
rect 12416 6500 12440 6502
rect 12496 6500 12502 6502
rect 12194 6491 12502 6500
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12084 5710 12112 6394
rect 12176 6254 12204 6394
rect 12346 6352 12402 6361
rect 12346 6287 12348 6296
rect 12400 6287 12402 6296
rect 12348 6258 12400 6264
rect 12636 6254 12664 7534
rect 12716 7472 12768 7478
rect 12716 7414 12768 7420
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 12084 5370 12112 5646
rect 12176 5642 12204 6054
rect 12636 5846 12664 6190
rect 12728 5914 12756 7414
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12714 5808 12770 5817
rect 12714 5743 12770 5752
rect 12728 5710 12756 5743
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12164 5636 12216 5642
rect 12164 5578 12216 5584
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12194 5468 12502 5477
rect 12194 5466 12200 5468
rect 12256 5466 12280 5468
rect 12336 5466 12360 5468
rect 12416 5466 12440 5468
rect 12496 5466 12502 5468
rect 12256 5414 12258 5466
rect 12438 5414 12440 5466
rect 12194 5412 12200 5414
rect 12256 5412 12280 5414
rect 12336 5412 12360 5414
rect 12416 5412 12440 5414
rect 12496 5412 12502 5414
rect 12194 5403 12502 5412
rect 12072 5364 12124 5370
rect 12636 5352 12664 5510
rect 12072 5306 12124 5312
rect 12452 5324 12664 5352
rect 12256 5296 12308 5302
rect 12070 5264 12126 5273
rect 12070 5199 12126 5208
rect 12254 5264 12256 5273
rect 12308 5264 12310 5273
rect 12254 5199 12310 5208
rect 12084 5030 12112 5199
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12072 5024 12124 5030
rect 11978 4992 12034 5001
rect 12072 4966 12124 4972
rect 12164 5024 12216 5030
rect 12164 4966 12216 4972
rect 11978 4927 12034 4936
rect 11992 4282 12020 4927
rect 12070 4584 12126 4593
rect 12070 4519 12126 4528
rect 11980 4276 12032 4282
rect 12084 4264 12112 4519
rect 12176 4486 12204 4966
rect 12268 4622 12296 5102
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12452 4554 12480 5324
rect 12532 5160 12584 5166
rect 12532 5102 12584 5108
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12194 4380 12502 4389
rect 12194 4378 12200 4380
rect 12256 4378 12280 4380
rect 12336 4378 12360 4380
rect 12416 4378 12440 4380
rect 12496 4378 12502 4380
rect 12256 4326 12258 4378
rect 12438 4326 12440 4378
rect 12194 4324 12200 4326
rect 12256 4324 12280 4326
rect 12336 4324 12360 4326
rect 12416 4324 12440 4326
rect 12496 4324 12502 4326
rect 12194 4315 12502 4324
rect 12440 4276 12492 4282
rect 12084 4236 12204 4264
rect 11980 4218 12032 4224
rect 12176 4146 12204 4236
rect 12440 4218 12492 4224
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12072 4072 12124 4078
rect 11992 4032 12072 4060
rect 11992 3602 12020 4032
rect 12348 4072 12400 4078
rect 12072 4014 12124 4020
rect 12346 4040 12348 4049
rect 12400 4040 12402 4049
rect 12346 3975 12402 3984
rect 12072 3936 12124 3942
rect 12072 3878 12124 3884
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 12084 3194 12112 3878
rect 12452 3466 12480 4218
rect 12544 3738 12572 5102
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12636 3602 12664 4490
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12194 3292 12502 3301
rect 12194 3290 12200 3292
rect 12256 3290 12280 3292
rect 12336 3290 12360 3292
rect 12416 3290 12440 3292
rect 12496 3290 12502 3292
rect 12256 3238 12258 3290
rect 12438 3238 12440 3290
rect 12194 3236 12200 3238
rect 12256 3236 12280 3238
rect 12336 3236 12360 3238
rect 12416 3236 12440 3238
rect 12496 3236 12502 3238
rect 12194 3227 12502 3236
rect 12636 3194 12664 3334
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12728 3126 12756 5510
rect 12820 4690 12848 8350
rect 13176 8298 13228 8304
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12912 7478 12940 8026
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 6730 12940 7142
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 13004 6202 13032 8230
rect 13464 8090 13492 11614
rect 13648 9602 13676 14350
rect 13740 14074 13768 14894
rect 13832 14793 13860 15302
rect 13818 14784 13874 14793
rect 13818 14719 13874 14728
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13820 14000 13872 14006
rect 13818 13968 13820 13977
rect 13872 13968 13874 13977
rect 13818 13903 13874 13912
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13740 13530 13768 13806
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13832 12442 13860 12786
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13728 12096 13780 12102
rect 13726 12064 13728 12073
rect 13780 12064 13782 12073
rect 13726 11999 13782 12008
rect 13818 11928 13874 11937
rect 13818 11863 13820 11872
rect 13872 11863 13874 11872
rect 13820 11834 13872 11840
rect 13924 11642 13952 15302
rect 14292 15026 14320 15506
rect 14568 15502 14596 19230
rect 14646 19200 14702 20000
rect 15014 19200 15070 20000
rect 15382 19200 15438 20000
rect 15488 19230 15700 19258
rect 14660 17898 14688 19200
rect 14660 17870 14872 17898
rect 14646 16688 14702 16697
rect 14646 16623 14648 16632
rect 14700 16623 14702 16632
rect 14648 16594 14700 16600
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 14464 15428 14516 15434
rect 14464 15370 14516 15376
rect 14280 15020 14332 15026
rect 14280 14962 14332 14968
rect 14068 14716 14376 14725
rect 14068 14714 14074 14716
rect 14130 14714 14154 14716
rect 14210 14714 14234 14716
rect 14290 14714 14314 14716
rect 14370 14714 14376 14716
rect 14130 14662 14132 14714
rect 14312 14662 14314 14714
rect 14068 14660 14074 14662
rect 14130 14660 14154 14662
rect 14210 14660 14234 14662
rect 14290 14660 14314 14662
rect 14370 14660 14376 14662
rect 14068 14651 14376 14660
rect 14372 14544 14424 14550
rect 14278 14512 14334 14521
rect 14372 14486 14424 14492
rect 14278 14447 14334 14456
rect 14292 14278 14320 14447
rect 14280 14272 14332 14278
rect 14278 14240 14280 14249
rect 14332 14240 14334 14249
rect 14278 14175 14334 14184
rect 14384 13734 14412 14486
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14068 13628 14376 13637
rect 14068 13626 14074 13628
rect 14130 13626 14154 13628
rect 14210 13626 14234 13628
rect 14290 13626 14314 13628
rect 14370 13626 14376 13628
rect 14130 13574 14132 13626
rect 14312 13574 14314 13626
rect 14068 13572 14074 13574
rect 14130 13572 14154 13574
rect 14210 13572 14234 13574
rect 14290 13572 14314 13574
rect 14370 13572 14376 13574
rect 14068 13563 14376 13572
rect 14094 13288 14150 13297
rect 14094 13223 14150 13232
rect 14372 13252 14424 13258
rect 14108 13190 14136 13223
rect 14372 13194 14424 13200
rect 14096 13184 14148 13190
rect 14096 13126 14148 13132
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14200 12714 14228 13126
rect 14384 12918 14412 13194
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 14068 12540 14376 12549
rect 14068 12538 14074 12540
rect 14130 12538 14154 12540
rect 14210 12538 14234 12540
rect 14290 12538 14314 12540
rect 14370 12538 14376 12540
rect 14130 12486 14132 12538
rect 14312 12486 14314 12538
rect 14068 12484 14074 12486
rect 14130 12484 14154 12486
rect 14210 12484 14234 12486
rect 14290 12484 14314 12486
rect 14370 12484 14376 12486
rect 14068 12475 14376 12484
rect 14370 12336 14426 12345
rect 14370 12271 14426 12280
rect 13832 11626 13952 11642
rect 13820 11620 13952 11626
rect 13872 11614 13952 11620
rect 13820 11562 13872 11568
rect 13912 11552 13964 11558
rect 14384 11540 14412 12271
rect 14476 11898 14504 15370
rect 14556 15360 14608 15366
rect 14554 15328 14556 15337
rect 14608 15328 14610 15337
rect 14554 15263 14610 15272
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 14568 13326 14596 15098
rect 14648 13796 14700 13802
rect 14648 13738 14700 13744
rect 14660 13394 14688 13738
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14752 13138 14780 15438
rect 14844 15094 14872 17870
rect 15028 15570 15056 19200
rect 15396 19122 15424 19200
rect 15488 19122 15516 19230
rect 15396 19094 15516 19122
rect 15672 18034 15700 19230
rect 15750 19200 15806 20000
rect 16118 19200 16174 20000
rect 15764 18170 15792 19200
rect 15764 18142 15884 18170
rect 15672 18006 15792 18034
rect 15658 17912 15714 17921
rect 15658 17847 15714 17856
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 14924 15428 14976 15434
rect 14924 15370 14976 15376
rect 14832 15088 14884 15094
rect 14832 15030 14884 15036
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14568 13110 14780 13138
rect 14568 12306 14596 13110
rect 14738 13016 14794 13025
rect 14738 12951 14740 12960
rect 14792 12951 14794 12960
rect 14740 12922 14792 12928
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14556 12300 14608 12306
rect 14556 12242 14608 12248
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14660 11694 14688 12174
rect 14752 11898 14780 12786
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14384 11512 14504 11540
rect 13912 11494 13964 11500
rect 13556 9574 13676 9602
rect 13820 9580 13872 9586
rect 13556 8498 13584 9574
rect 13820 9522 13872 9528
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13648 9178 13676 9454
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13740 8634 13768 8774
rect 13832 8634 13860 9522
rect 13924 9194 13952 11494
rect 14068 11452 14376 11461
rect 14068 11450 14074 11452
rect 14130 11450 14154 11452
rect 14210 11450 14234 11452
rect 14290 11450 14314 11452
rect 14370 11450 14376 11452
rect 14130 11398 14132 11450
rect 14312 11398 14314 11450
rect 14068 11396 14074 11398
rect 14130 11396 14154 11398
rect 14210 11396 14234 11398
rect 14290 11396 14314 11398
rect 14370 11396 14376 11398
rect 14068 11387 14376 11396
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14108 10742 14136 10950
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14068 10364 14376 10373
rect 14068 10362 14074 10364
rect 14130 10362 14154 10364
rect 14210 10362 14234 10364
rect 14290 10362 14314 10364
rect 14370 10362 14376 10364
rect 14130 10310 14132 10362
rect 14312 10310 14314 10362
rect 14068 10308 14074 10310
rect 14130 10308 14154 10310
rect 14210 10308 14234 10310
rect 14290 10308 14314 10310
rect 14370 10308 14376 10310
rect 14068 10299 14376 10308
rect 14476 9994 14504 11512
rect 14660 11218 14688 11630
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14554 11112 14610 11121
rect 14554 11047 14556 11056
rect 14608 11047 14610 11056
rect 14556 11018 14608 11024
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14280 9988 14332 9994
rect 14280 9930 14332 9936
rect 14464 9988 14516 9994
rect 14464 9930 14516 9936
rect 14292 9722 14320 9930
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14568 9722 14596 9862
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14068 9276 14376 9285
rect 14068 9274 14074 9276
rect 14130 9274 14154 9276
rect 14210 9274 14234 9276
rect 14290 9274 14314 9276
rect 14370 9274 14376 9276
rect 14130 9222 14132 9274
rect 14312 9222 14314 9274
rect 14068 9220 14074 9222
rect 14130 9220 14154 9222
rect 14210 9220 14234 9222
rect 14290 9220 14314 9222
rect 14370 9220 14376 9222
rect 14068 9211 14376 9220
rect 13924 9166 14044 9194
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13924 8430 13952 9046
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13084 7812 13136 7818
rect 13084 7754 13136 7760
rect 13096 7002 13124 7754
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13464 7546 13492 7686
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 13096 6254 13124 6938
rect 12912 6174 13032 6202
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 12808 4684 12860 4690
rect 12808 4626 12860 4632
rect 12820 4486 12848 4626
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12912 4282 12940 6174
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 12900 4276 12952 4282
rect 12900 4218 12952 4224
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12820 3194 12848 3878
rect 12912 3534 12940 3878
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12716 3120 12768 3126
rect 11978 3088 12034 3097
rect 12716 3062 12768 3068
rect 11978 3023 12034 3032
rect 11992 2990 12020 3023
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 11900 2746 12020 2774
rect 11992 2446 12020 2746
rect 11704 2440 11756 2446
rect 11980 2440 12032 2446
rect 11704 2382 11756 2388
rect 11900 2388 11980 2394
rect 11900 2382 12032 2388
rect 11612 2032 11664 2038
rect 11612 1974 11664 1980
rect 11716 1562 11744 2382
rect 11900 2366 12020 2382
rect 11704 1556 11756 1562
rect 11704 1498 11756 1504
rect 11900 800 11928 2366
rect 12084 2088 12112 2790
rect 13004 2774 13032 6054
rect 13188 5352 13216 7142
rect 13372 6730 13400 7346
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 13360 6724 13412 6730
rect 13360 6666 13412 6672
rect 13280 5930 13308 6666
rect 13464 6186 13492 7278
rect 13452 6180 13504 6186
rect 13452 6122 13504 6128
rect 13280 5902 13492 5930
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13268 5568 13320 5574
rect 13268 5510 13320 5516
rect 13096 5324 13216 5352
rect 13096 3738 13124 5324
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 13188 4486 13216 5170
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13280 4146 13308 5510
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 13188 3602 13216 4014
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13188 2854 13216 3334
rect 13280 2990 13308 4082
rect 13372 4078 13400 5714
rect 13464 5642 13492 5902
rect 13452 5636 13504 5642
rect 13452 5578 13504 5584
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13464 4758 13492 5102
rect 13452 4752 13504 4758
rect 13452 4694 13504 4700
rect 13360 4072 13412 4078
rect 13412 4032 13492 4060
rect 13360 4014 13412 4020
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 12912 2746 13032 2774
rect 12912 2446 12940 2746
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 12194 2204 12502 2213
rect 12194 2202 12200 2204
rect 12256 2202 12280 2204
rect 12336 2202 12360 2204
rect 12416 2202 12440 2204
rect 12496 2202 12502 2204
rect 12256 2150 12258 2202
rect 12438 2150 12440 2202
rect 12194 2148 12200 2150
rect 12256 2148 12280 2150
rect 12336 2148 12360 2150
rect 12416 2148 12440 2150
rect 12496 2148 12502 2150
rect 12194 2139 12502 2148
rect 12084 2060 12296 2088
rect 12268 800 12296 2060
rect 12636 800 12664 2382
rect 13084 2372 13136 2378
rect 13084 2314 13136 2320
rect 13096 2258 13124 2314
rect 13004 2230 13124 2258
rect 13004 800 13032 2230
rect 13372 800 13400 3674
rect 13464 2854 13492 4032
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 13556 2446 13584 7686
rect 13648 6866 13676 7822
rect 13832 7290 13860 8298
rect 14016 8242 14044 9166
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 13924 8214 14044 8242
rect 13924 7970 13952 8214
rect 14068 8188 14376 8197
rect 14068 8186 14074 8188
rect 14130 8186 14154 8188
rect 14210 8186 14234 8188
rect 14290 8186 14314 8188
rect 14370 8186 14376 8188
rect 14130 8134 14132 8186
rect 14312 8134 14314 8186
rect 14068 8132 14074 8134
rect 14130 8132 14154 8134
rect 14210 8132 14234 8134
rect 14290 8132 14314 8134
rect 14370 8132 14376 8134
rect 14068 8123 14376 8132
rect 14476 8090 14504 8774
rect 14568 8634 14596 8774
rect 14660 8634 14688 10950
rect 14844 10146 14872 14894
rect 14936 12850 14964 15370
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14924 12708 14976 12714
rect 14924 12650 14976 12656
rect 14936 12306 14964 12650
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 15028 11014 15056 14350
rect 15120 13258 15148 17002
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 15120 13161 15148 13194
rect 15106 13152 15162 13161
rect 15106 13087 15162 13096
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 15120 10826 15148 12922
rect 15212 12850 15240 17070
rect 15304 16658 15332 17750
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15292 16652 15344 16658
rect 15292 16594 15344 16600
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15304 11898 15332 15506
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15212 11218 15240 11494
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15200 11212 15252 11218
rect 15200 11154 15252 11160
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 14752 10118 14872 10146
rect 15028 10798 15148 10826
rect 14556 8628 14608 8634
rect 14556 8570 14608 8576
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14556 8424 14608 8430
rect 14556 8366 14608 8372
rect 14568 8294 14596 8366
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14464 8084 14516 8090
rect 14464 8026 14516 8032
rect 13924 7942 14044 7970
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13740 7262 13860 7290
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13648 5114 13676 6598
rect 13740 6338 13768 7262
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13832 6458 13860 7142
rect 13924 6882 13952 7822
rect 14016 7206 14044 7942
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 14384 7342 14412 7754
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14068 7100 14376 7109
rect 14068 7098 14074 7100
rect 14130 7098 14154 7100
rect 14210 7098 14234 7100
rect 14290 7098 14314 7100
rect 14370 7098 14376 7100
rect 14130 7046 14132 7098
rect 14312 7046 14314 7098
rect 14068 7044 14074 7046
rect 14130 7044 14154 7046
rect 14210 7044 14234 7046
rect 14290 7044 14314 7046
rect 14370 7044 14376 7046
rect 14068 7035 14376 7044
rect 13924 6854 14044 6882
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13740 6310 13860 6338
rect 13726 6216 13782 6225
rect 13726 6151 13728 6160
rect 13780 6151 13782 6160
rect 13728 6122 13780 6128
rect 13740 5914 13768 6122
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13740 5370 13768 5850
rect 13832 5574 13860 6310
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13648 5086 13768 5114
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13648 4690 13676 4966
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13740 4026 13768 5086
rect 13832 4282 13860 5510
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 13648 3998 13768 4026
rect 13648 3398 13676 3998
rect 13820 3936 13872 3942
rect 13726 3904 13782 3913
rect 13820 3878 13872 3884
rect 13726 3839 13782 3848
rect 13740 3670 13768 3839
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13648 2990 13676 3334
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13544 2440 13596 2446
rect 13544 2382 13596 2388
rect 13740 800 13768 3470
rect 13832 3058 13860 3878
rect 13924 3466 13952 6734
rect 14016 6304 14044 6854
rect 14096 6316 14148 6322
rect 14016 6276 14096 6304
rect 14096 6258 14148 6264
rect 14108 6225 14136 6258
rect 14094 6216 14150 6225
rect 14094 6151 14150 6160
rect 14068 6012 14376 6021
rect 14068 6010 14074 6012
rect 14130 6010 14154 6012
rect 14210 6010 14234 6012
rect 14290 6010 14314 6012
rect 14370 6010 14376 6012
rect 14130 5958 14132 6010
rect 14312 5958 14314 6010
rect 14068 5956 14074 5958
rect 14130 5956 14154 5958
rect 14210 5956 14234 5958
rect 14290 5956 14314 5958
rect 14370 5956 14376 5958
rect 14068 5947 14376 5956
rect 14188 5704 14240 5710
rect 14188 5646 14240 5652
rect 14200 5370 14228 5646
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14108 5137 14136 5170
rect 14292 5166 14320 5578
rect 14476 5250 14504 7686
rect 14568 7478 14596 8230
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14568 7002 14596 7142
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14568 6458 14596 6598
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14660 6236 14688 8434
rect 14752 7750 14780 10118
rect 15028 10062 15056 10798
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15016 10056 15068 10062
rect 15014 10024 15016 10033
rect 15068 10024 15070 10033
rect 14832 9988 14884 9994
rect 15014 9959 15070 9968
rect 14832 9930 14884 9936
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14752 6798 14780 7142
rect 14740 6792 14792 6798
rect 14740 6734 14792 6740
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14752 6390 14780 6598
rect 14844 6458 14872 9930
rect 15014 9752 15070 9761
rect 15014 9687 15070 9696
rect 15028 9654 15056 9687
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 14936 9178 14964 9522
rect 14924 9172 14976 9178
rect 14924 9114 14976 9120
rect 15120 9042 15148 10066
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14936 8430 14964 8910
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14936 7954 14964 8366
rect 15212 8362 15240 11018
rect 15304 10470 15332 11290
rect 15396 11082 15424 17138
rect 15568 16516 15620 16522
rect 15568 16458 15620 16464
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15488 16046 15516 16390
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15488 14414 15516 15982
rect 15580 15162 15608 16458
rect 15672 16182 15700 17847
rect 15660 16176 15712 16182
rect 15660 16118 15712 16124
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15488 14006 15516 14214
rect 15476 14000 15528 14006
rect 15476 13942 15528 13948
rect 15566 13968 15622 13977
rect 15672 13954 15700 14962
rect 15764 14346 15792 18006
rect 15856 16998 15884 18142
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 16028 16992 16080 16998
rect 16028 16934 16080 16940
rect 15844 15088 15896 15094
rect 15844 15030 15896 15036
rect 15752 14340 15804 14346
rect 15752 14282 15804 14288
rect 15672 13926 15792 13954
rect 15566 13903 15622 13912
rect 15476 13728 15528 13734
rect 15476 13670 15528 13676
rect 15488 13258 15516 13670
rect 15476 13252 15528 13258
rect 15476 13194 15528 13200
rect 15580 12850 15608 13903
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15580 12442 15608 12786
rect 15672 12714 15700 13806
rect 15764 13326 15792 13926
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15660 12708 15712 12714
rect 15660 12650 15712 12656
rect 15764 12594 15792 13262
rect 15672 12566 15792 12594
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15566 10024 15622 10033
rect 15566 9959 15622 9968
rect 15580 9926 15608 9959
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15672 9674 15700 12566
rect 15750 12472 15806 12481
rect 15750 12407 15806 12416
rect 15764 11830 15792 12407
rect 15856 12374 15884 15030
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15844 12368 15896 12374
rect 15844 12310 15896 12316
rect 15948 12306 15976 14282
rect 15936 12300 15988 12306
rect 15936 12242 15988 12248
rect 15752 11824 15804 11830
rect 15752 11766 15804 11772
rect 16040 11762 16068 16934
rect 16132 12986 16160 19200
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15488 9646 15700 9674
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15304 8974 15332 9454
rect 15396 8974 15424 9590
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15396 8634 15424 8910
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15200 8356 15252 8362
rect 15200 8298 15252 8304
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 15016 7744 15068 7750
rect 14936 7704 15016 7732
rect 14936 6798 14964 7704
rect 15016 7686 15068 7692
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 15028 6934 15056 7482
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 15016 6928 15068 6934
rect 15016 6870 15068 6876
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14740 6384 14792 6390
rect 14740 6326 14792 6332
rect 14660 6208 14872 6236
rect 14646 5808 14702 5817
rect 14646 5743 14702 5752
rect 14660 5642 14688 5743
rect 14648 5636 14700 5642
rect 14648 5578 14700 5584
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14476 5222 14596 5250
rect 14280 5160 14332 5166
rect 14094 5128 14150 5137
rect 14280 5102 14332 5108
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14094 5063 14150 5072
rect 14068 4924 14376 4933
rect 14068 4922 14074 4924
rect 14130 4922 14154 4924
rect 14210 4922 14234 4924
rect 14290 4922 14314 4924
rect 14370 4922 14376 4924
rect 14130 4870 14132 4922
rect 14312 4870 14314 4922
rect 14068 4868 14074 4870
rect 14130 4868 14154 4870
rect 14210 4868 14234 4870
rect 14290 4868 14314 4870
rect 14370 4868 14376 4870
rect 14068 4859 14376 4868
rect 14476 4622 14504 5102
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14464 4480 14516 4486
rect 14462 4448 14464 4457
rect 14516 4448 14518 4457
rect 14462 4383 14518 4392
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14068 3836 14376 3845
rect 14068 3834 14074 3836
rect 14130 3834 14154 3836
rect 14210 3834 14234 3836
rect 14290 3834 14314 3836
rect 14370 3834 14376 3836
rect 14130 3782 14132 3834
rect 14312 3782 14314 3834
rect 14068 3780 14074 3782
rect 14130 3780 14154 3782
rect 14210 3780 14234 3782
rect 14290 3780 14314 3782
rect 14370 3780 14376 3782
rect 14068 3771 14376 3780
rect 14370 3496 14426 3505
rect 13912 3460 13964 3466
rect 14370 3431 14426 3440
rect 13912 3402 13964 3408
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 13818 2952 13874 2961
rect 13818 2887 13820 2896
rect 13872 2887 13874 2896
rect 13820 2858 13872 2864
rect 13924 2530 13952 3402
rect 14094 3088 14150 3097
rect 14094 3023 14096 3032
rect 14148 3023 14150 3032
rect 14096 2994 14148 3000
rect 14384 2990 14412 3431
rect 14476 3398 14504 4218
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14568 3058 14596 5222
rect 14648 5092 14700 5098
rect 14648 5034 14700 5040
rect 14660 4690 14688 5034
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14660 4078 14688 4626
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14568 2774 14596 2994
rect 14068 2748 14376 2757
rect 14068 2746 14074 2748
rect 14130 2746 14154 2748
rect 14210 2746 14234 2748
rect 14290 2746 14314 2748
rect 14370 2746 14376 2748
rect 14130 2694 14132 2746
rect 14312 2694 14314 2746
rect 14068 2692 14074 2694
rect 14130 2692 14154 2694
rect 14210 2692 14234 2694
rect 14290 2692 14314 2694
rect 14370 2692 14376 2694
rect 14068 2683 14376 2692
rect 14476 2746 14596 2774
rect 14370 2544 14426 2553
rect 13924 2502 14136 2530
rect 14108 800 14136 2502
rect 14370 2479 14426 2488
rect 14384 2446 14412 2479
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 14476 800 14504 2746
rect 14660 2145 14688 3878
rect 14752 3534 14780 5510
rect 14844 4826 14872 6208
rect 14936 5953 14964 6734
rect 15028 6390 15056 6870
rect 15016 6384 15068 6390
rect 15016 6326 15068 6332
rect 14922 5944 14978 5953
rect 14922 5879 14978 5888
rect 15120 5778 15148 7346
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15106 5536 15162 5545
rect 15106 5471 15162 5480
rect 15014 5400 15070 5409
rect 15120 5370 15148 5471
rect 15014 5335 15070 5344
rect 15108 5364 15160 5370
rect 15028 5302 15056 5335
rect 15108 5306 15160 5312
rect 15016 5296 15068 5302
rect 15016 5238 15068 5244
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14844 4049 14872 4082
rect 14830 4040 14886 4049
rect 14830 3975 14886 3984
rect 14936 3670 14964 5170
rect 14924 3664 14976 3670
rect 14924 3606 14976 3612
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14646 2136 14702 2145
rect 14646 2071 14702 2080
rect 14844 800 14872 3538
rect 15028 3534 15056 5238
rect 15108 5024 15160 5030
rect 15108 4966 15160 4972
rect 15120 4622 15148 4966
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 15120 3738 15148 4558
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 15016 3528 15068 3534
rect 15016 3470 15068 3476
rect 15016 3392 15068 3398
rect 15016 3334 15068 3340
rect 15028 2650 15056 3334
rect 15016 2644 15068 2650
rect 15016 2586 15068 2592
rect 15212 2514 15240 8298
rect 15396 7546 15424 8570
rect 15488 8566 15516 9646
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 15488 7834 15516 8502
rect 15488 7806 15608 7834
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15292 6724 15344 6730
rect 15292 6666 15344 6672
rect 15304 5273 15332 6666
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 15396 5914 15424 6258
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15290 5264 15346 5273
rect 15290 5199 15346 5208
rect 15396 4622 15424 5510
rect 15488 5352 15516 7686
rect 15580 7274 15608 7806
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15568 6112 15620 6118
rect 15566 6080 15568 6089
rect 15620 6080 15622 6089
rect 15566 6015 15622 6024
rect 15568 5704 15620 5710
rect 15566 5672 15568 5681
rect 15620 5672 15622 5681
rect 15566 5607 15622 5616
rect 15488 5324 15608 5352
rect 15476 5228 15528 5234
rect 15476 5170 15528 5176
rect 15384 4616 15436 4622
rect 15304 4576 15384 4604
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15304 2394 15332 4576
rect 15384 4558 15436 4564
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15396 4185 15424 4422
rect 15382 4176 15438 4185
rect 15382 4111 15438 4120
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 15212 2366 15332 2394
rect 15212 800 15240 2366
rect 15396 2106 15424 2790
rect 15488 2514 15516 5170
rect 15580 3602 15608 5324
rect 15672 4146 15700 7686
rect 15844 7540 15896 7546
rect 15844 7482 15896 7488
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 15672 2774 15700 4082
rect 15764 4078 15792 6394
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 15856 3058 15884 7482
rect 15948 5642 15976 10406
rect 15936 5636 15988 5642
rect 15936 5578 15988 5584
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15580 2746 15700 2774
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15384 2100 15436 2106
rect 15384 2042 15436 2048
rect 15580 800 15608 2746
rect 15948 800 15976 4966
rect 16040 4486 16068 11086
rect 16224 10062 16252 14350
rect 16316 11354 16344 16730
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16408 12481 16436 16186
rect 16394 12472 16450 12481
rect 16394 12407 16450 12416
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16028 4480 16080 4486
rect 16028 4422 16080 4428
rect 8680 734 8892 762
rect 8942 0 8998 800
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 10046 0 10102 800
rect 10414 0 10470 800
rect 10782 0 10838 800
rect 11150 0 11206 800
rect 11518 0 11574 800
rect 11886 0 11942 800
rect 12254 0 12310 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 15934 0 15990 800
<< via2 >>
rect 1306 18536 1362 18592
rect 2318 17584 2374 17640
rect 2778 19080 2834 19136
rect 1950 16668 1952 16688
rect 1952 16668 2004 16688
rect 2004 16668 2006 16688
rect 1950 16632 2006 16668
rect 1490 15680 1546 15736
rect 2318 16108 2374 16144
rect 2318 16088 2320 16108
rect 2320 16088 2372 16108
rect 2372 16088 2374 16108
rect 2830 16890 2886 16892
rect 2910 16890 2966 16892
rect 2990 16890 3046 16892
rect 3070 16890 3126 16892
rect 2830 16838 2876 16890
rect 2876 16838 2886 16890
rect 2910 16838 2940 16890
rect 2940 16838 2952 16890
rect 2952 16838 2966 16890
rect 2990 16838 3004 16890
rect 3004 16838 3016 16890
rect 3016 16838 3046 16890
rect 3070 16838 3080 16890
rect 3080 16838 3126 16890
rect 2830 16836 2886 16838
rect 2910 16836 2966 16838
rect 2990 16836 3046 16838
rect 3070 16836 3126 16838
rect 2042 15408 2098 15464
rect 2134 15308 2136 15328
rect 2136 15308 2188 15328
rect 2188 15308 2190 15328
rect 2134 15272 2190 15308
rect 2410 15308 2412 15328
rect 2412 15308 2464 15328
rect 2464 15308 2466 15328
rect 2410 15272 2466 15308
rect 1950 15020 2006 15056
rect 1950 15000 1952 15020
rect 1952 15000 2004 15020
rect 2004 15000 2006 15020
rect 1490 14764 1492 14784
rect 1492 14764 1544 14784
rect 1544 14764 1546 14784
rect 1490 14728 1546 14764
rect 1950 13912 2006 13968
rect 1490 13796 1546 13832
rect 1490 13776 1492 13796
rect 1492 13776 1544 13796
rect 1544 13776 1546 13796
rect 1490 12824 1546 12880
rect 1490 11892 1546 11928
rect 1490 11872 1492 11892
rect 1492 11872 1544 11892
rect 1544 11872 1546 11892
rect 1490 10956 1492 10976
rect 1492 10956 1544 10976
rect 1544 10956 1546 10976
rect 1490 10920 1546 10956
rect 1490 9968 1546 10024
rect 1582 9560 1638 9616
rect 1490 9016 1546 9072
rect 1490 8084 1546 8120
rect 1490 8064 1492 8084
rect 1492 8064 1544 8084
rect 1544 8064 1546 8084
rect 1490 7148 1492 7168
rect 1492 7148 1544 7168
rect 1544 7148 1546 7168
rect 1490 7112 1546 7148
rect 1490 6180 1546 6216
rect 1490 6160 1492 6180
rect 1492 6160 1544 6180
rect 1544 6160 1546 6180
rect 2686 16360 2742 16416
rect 3146 16360 3202 16416
rect 2830 15802 2886 15804
rect 2910 15802 2966 15804
rect 2990 15802 3046 15804
rect 3070 15802 3126 15804
rect 2830 15750 2876 15802
rect 2876 15750 2886 15802
rect 2910 15750 2940 15802
rect 2940 15750 2952 15802
rect 2952 15750 2966 15802
rect 2990 15750 3004 15802
rect 3004 15750 3016 15802
rect 3016 15750 3046 15802
rect 3070 15750 3080 15802
rect 3080 15750 3126 15802
rect 2830 15748 2886 15750
rect 2910 15748 2966 15750
rect 2990 15748 3046 15750
rect 3070 15748 3126 15750
rect 3054 14864 3110 14920
rect 3422 15544 3478 15600
rect 2830 14714 2886 14716
rect 2910 14714 2966 14716
rect 2990 14714 3046 14716
rect 3070 14714 3126 14716
rect 2830 14662 2876 14714
rect 2876 14662 2886 14714
rect 2910 14662 2940 14714
rect 2940 14662 2952 14714
rect 2952 14662 2966 14714
rect 2990 14662 3004 14714
rect 3004 14662 3016 14714
rect 3016 14662 3046 14714
rect 3070 14662 3080 14714
rect 3080 14662 3126 14714
rect 2830 14660 2886 14662
rect 2910 14660 2966 14662
rect 2990 14660 3046 14662
rect 3070 14660 3126 14662
rect 2830 13626 2886 13628
rect 2910 13626 2966 13628
rect 2990 13626 3046 13628
rect 3070 13626 3126 13628
rect 2830 13574 2876 13626
rect 2876 13574 2886 13626
rect 2910 13574 2940 13626
rect 2940 13574 2952 13626
rect 2952 13574 2966 13626
rect 2990 13574 3004 13626
rect 3004 13574 3016 13626
rect 3016 13574 3046 13626
rect 3070 13574 3080 13626
rect 3080 13574 3126 13626
rect 2830 13572 2886 13574
rect 2910 13572 2966 13574
rect 2990 13572 3046 13574
rect 3070 13572 3126 13574
rect 2686 13232 2742 13288
rect 2830 12538 2886 12540
rect 2910 12538 2966 12540
rect 2990 12538 3046 12540
rect 3070 12538 3126 12540
rect 2830 12486 2876 12538
rect 2876 12486 2886 12538
rect 2910 12486 2940 12538
rect 2940 12486 2952 12538
rect 2952 12486 2966 12538
rect 2990 12486 3004 12538
rect 3004 12486 3016 12538
rect 3016 12486 3046 12538
rect 3070 12486 3080 12538
rect 3080 12486 3126 12538
rect 2830 12484 2886 12486
rect 2910 12484 2966 12486
rect 2990 12484 3046 12486
rect 3070 12484 3126 12486
rect 3238 12552 3294 12608
rect 2830 11450 2886 11452
rect 2910 11450 2966 11452
rect 2990 11450 3046 11452
rect 3070 11450 3126 11452
rect 2830 11398 2876 11450
rect 2876 11398 2886 11450
rect 2910 11398 2940 11450
rect 2940 11398 2952 11450
rect 2952 11398 2966 11450
rect 2990 11398 3004 11450
rect 3004 11398 3016 11450
rect 3016 11398 3046 11450
rect 3070 11398 3080 11450
rect 3080 11398 3126 11450
rect 2830 11396 2886 11398
rect 2910 11396 2966 11398
rect 2990 11396 3046 11398
rect 3070 11396 3126 11398
rect 3238 11328 3294 11384
rect 2830 10362 2886 10364
rect 2910 10362 2966 10364
rect 2990 10362 3046 10364
rect 3070 10362 3126 10364
rect 2830 10310 2876 10362
rect 2876 10310 2886 10362
rect 2910 10310 2940 10362
rect 2940 10310 2952 10362
rect 2952 10310 2966 10362
rect 2990 10310 3004 10362
rect 3004 10310 3016 10362
rect 3016 10310 3046 10362
rect 3070 10310 3080 10362
rect 3080 10310 3126 10362
rect 2830 10308 2886 10310
rect 2910 10308 2966 10310
rect 2990 10308 3046 10310
rect 3070 10308 3126 10310
rect 2830 9274 2886 9276
rect 2910 9274 2966 9276
rect 2990 9274 3046 9276
rect 3070 9274 3126 9276
rect 2830 9222 2876 9274
rect 2876 9222 2886 9274
rect 2910 9222 2940 9274
rect 2940 9222 2952 9274
rect 2952 9222 2966 9274
rect 2990 9222 3004 9274
rect 3004 9222 3016 9274
rect 3016 9222 3046 9274
rect 3070 9222 3080 9274
rect 3080 9222 3126 9274
rect 2830 9220 2886 9222
rect 2910 9220 2966 9222
rect 2990 9220 3046 9222
rect 3070 9220 3126 9222
rect 3606 15272 3662 15328
rect 4704 17434 4760 17436
rect 4784 17434 4840 17436
rect 4864 17434 4920 17436
rect 4944 17434 5000 17436
rect 4704 17382 4750 17434
rect 4750 17382 4760 17434
rect 4784 17382 4814 17434
rect 4814 17382 4826 17434
rect 4826 17382 4840 17434
rect 4864 17382 4878 17434
rect 4878 17382 4890 17434
rect 4890 17382 4920 17434
rect 4944 17382 4954 17434
rect 4954 17382 5000 17434
rect 4704 17380 4760 17382
rect 4784 17380 4840 17382
rect 4864 17380 4920 17382
rect 4944 17380 5000 17382
rect 3882 15272 3938 15328
rect 3514 14864 3570 14920
rect 3422 14048 3478 14104
rect 2134 6604 2136 6624
rect 2136 6604 2188 6624
rect 2188 6604 2190 6624
rect 2134 6568 2190 6604
rect 2318 7268 2374 7304
rect 2318 7248 2320 7268
rect 2320 7248 2372 7268
rect 2372 7248 2374 7268
rect 1490 5208 1546 5264
rect 1490 4256 1546 4312
rect 1582 3984 1638 4040
rect 1858 3612 1860 3632
rect 1860 3612 1912 3632
rect 1912 3612 1914 3632
rect 1858 3576 1914 3612
rect 1582 3340 1584 3360
rect 1584 3340 1636 3360
rect 1636 3340 1638 3360
rect 1582 3304 1638 3340
rect 2830 8186 2886 8188
rect 2910 8186 2966 8188
rect 2990 8186 3046 8188
rect 3070 8186 3126 8188
rect 2830 8134 2876 8186
rect 2876 8134 2886 8186
rect 2910 8134 2940 8186
rect 2940 8134 2952 8186
rect 2952 8134 2966 8186
rect 2990 8134 3004 8186
rect 3004 8134 3016 8186
rect 3016 8134 3046 8186
rect 3070 8134 3080 8186
rect 3080 8134 3126 8186
rect 2830 8132 2886 8134
rect 2910 8132 2966 8134
rect 2990 8132 3046 8134
rect 3070 8132 3126 8134
rect 4066 15988 4068 16008
rect 4068 15988 4120 16008
rect 4120 15988 4122 16008
rect 4066 15952 4122 15988
rect 4710 17196 4766 17232
rect 4710 17176 4712 17196
rect 4712 17176 4764 17196
rect 4764 17176 4766 17196
rect 4526 16532 4528 16552
rect 4528 16532 4580 16552
rect 4580 16532 4582 16552
rect 4526 16496 4582 16532
rect 4342 15544 4398 15600
rect 5446 17040 5502 17096
rect 4704 16346 4760 16348
rect 4784 16346 4840 16348
rect 4864 16346 4920 16348
rect 4944 16346 5000 16348
rect 4704 16294 4750 16346
rect 4750 16294 4760 16346
rect 4784 16294 4814 16346
rect 4814 16294 4826 16346
rect 4826 16294 4840 16346
rect 4864 16294 4878 16346
rect 4878 16294 4890 16346
rect 4890 16294 4920 16346
rect 4944 16294 4954 16346
rect 4954 16294 5000 16346
rect 4704 16292 4760 16294
rect 4784 16292 4840 16294
rect 4864 16292 4920 16294
rect 4944 16292 5000 16294
rect 4618 15680 4674 15736
rect 4704 15258 4760 15260
rect 4784 15258 4840 15260
rect 4864 15258 4920 15260
rect 4944 15258 5000 15260
rect 4704 15206 4750 15258
rect 4750 15206 4760 15258
rect 4784 15206 4814 15258
rect 4814 15206 4826 15258
rect 4826 15206 4840 15258
rect 4864 15206 4878 15258
rect 4878 15206 4890 15258
rect 4890 15206 4920 15258
rect 4944 15206 4954 15258
rect 4954 15206 5000 15258
rect 4704 15204 4760 15206
rect 4784 15204 4840 15206
rect 4864 15204 4920 15206
rect 4944 15204 5000 15206
rect 4250 14456 4306 14512
rect 4250 13948 4252 13968
rect 4252 13948 4304 13968
rect 4304 13948 4306 13968
rect 4250 13912 4306 13948
rect 4158 13812 4160 13832
rect 4160 13812 4212 13832
rect 4212 13812 4214 13832
rect 4158 13776 4214 13812
rect 3882 12180 3884 12200
rect 3884 12180 3936 12200
rect 3936 12180 3938 12200
rect 3882 12144 3938 12180
rect 2830 7098 2886 7100
rect 2910 7098 2966 7100
rect 2990 7098 3046 7100
rect 3070 7098 3126 7100
rect 2830 7046 2876 7098
rect 2876 7046 2886 7098
rect 2910 7046 2940 7098
rect 2940 7046 2952 7098
rect 2952 7046 2966 7098
rect 2990 7046 3004 7098
rect 3004 7046 3016 7098
rect 3016 7046 3046 7098
rect 3070 7046 3080 7098
rect 3080 7046 3126 7098
rect 2830 7044 2886 7046
rect 2910 7044 2966 7046
rect 2990 7044 3046 7046
rect 3070 7044 3126 7046
rect 3606 7792 3662 7848
rect 2502 5616 2558 5672
rect 2502 5228 2558 5264
rect 2502 5208 2504 5228
rect 2504 5208 2556 5228
rect 2556 5208 2558 5228
rect 2778 6196 2780 6216
rect 2780 6196 2832 6216
rect 2832 6196 2834 6216
rect 2778 6160 2834 6196
rect 2830 6010 2886 6012
rect 2910 6010 2966 6012
rect 2990 6010 3046 6012
rect 3070 6010 3126 6012
rect 2830 5958 2876 6010
rect 2876 5958 2886 6010
rect 2910 5958 2940 6010
rect 2940 5958 2952 6010
rect 2952 5958 2966 6010
rect 2990 5958 3004 6010
rect 3004 5958 3016 6010
rect 3016 5958 3046 6010
rect 3070 5958 3080 6010
rect 3080 5958 3126 6010
rect 2830 5956 2886 5958
rect 2910 5956 2966 5958
rect 2990 5956 3046 5958
rect 3070 5956 3126 5958
rect 3146 5072 3202 5128
rect 2830 4922 2886 4924
rect 2910 4922 2966 4924
rect 2990 4922 3046 4924
rect 3070 4922 3126 4924
rect 2830 4870 2876 4922
rect 2876 4870 2886 4922
rect 2910 4870 2940 4922
rect 2940 4870 2952 4922
rect 2952 4870 2966 4922
rect 2990 4870 3004 4922
rect 3004 4870 3016 4922
rect 3016 4870 3046 4922
rect 3070 4870 3080 4922
rect 3080 4870 3126 4922
rect 2830 4868 2886 4870
rect 2910 4868 2966 4870
rect 2990 4868 3046 4870
rect 3070 4868 3126 4870
rect 3054 4664 3110 4720
rect 2778 4528 2834 4584
rect 3606 6160 3662 6216
rect 3330 5480 3386 5536
rect 2830 3834 2886 3836
rect 2910 3834 2966 3836
rect 2990 3834 3046 3836
rect 3070 3834 3126 3836
rect 2830 3782 2876 3834
rect 2876 3782 2886 3834
rect 2910 3782 2940 3834
rect 2940 3782 2952 3834
rect 2952 3782 2966 3834
rect 2990 3782 3004 3834
rect 3004 3782 3016 3834
rect 3016 3782 3046 3834
rect 3070 3782 3080 3834
rect 3080 3782 3126 3834
rect 2830 3780 2886 3782
rect 2910 3780 2966 3782
rect 2990 3780 3046 3782
rect 3070 3780 3126 3782
rect 4704 14170 4760 14172
rect 4784 14170 4840 14172
rect 4864 14170 4920 14172
rect 4944 14170 5000 14172
rect 4704 14118 4750 14170
rect 4750 14118 4760 14170
rect 4784 14118 4814 14170
rect 4814 14118 4826 14170
rect 4826 14118 4840 14170
rect 4864 14118 4878 14170
rect 4878 14118 4890 14170
rect 4890 14118 4920 14170
rect 4944 14118 4954 14170
rect 4954 14118 5000 14170
rect 4704 14116 4760 14118
rect 4784 14116 4840 14118
rect 4864 14116 4920 14118
rect 4944 14116 5000 14118
rect 5262 14184 5318 14240
rect 5630 15000 5686 15056
rect 6090 15952 6146 16008
rect 4704 13082 4760 13084
rect 4784 13082 4840 13084
rect 4864 13082 4920 13084
rect 4944 13082 5000 13084
rect 4704 13030 4750 13082
rect 4750 13030 4760 13082
rect 4784 13030 4814 13082
rect 4814 13030 4826 13082
rect 4826 13030 4840 13082
rect 4864 13030 4878 13082
rect 4878 13030 4890 13082
rect 4890 13030 4920 13082
rect 4944 13030 4954 13082
rect 4954 13030 5000 13082
rect 4704 13028 4760 13030
rect 4784 13028 4840 13030
rect 4864 13028 4920 13030
rect 4944 13028 5000 13030
rect 4704 11994 4760 11996
rect 4784 11994 4840 11996
rect 4864 11994 4920 11996
rect 4944 11994 5000 11996
rect 4704 11942 4750 11994
rect 4750 11942 4760 11994
rect 4784 11942 4814 11994
rect 4814 11942 4826 11994
rect 4826 11942 4840 11994
rect 4864 11942 4878 11994
rect 4878 11942 4890 11994
rect 4890 11942 4920 11994
rect 4944 11942 4954 11994
rect 4954 11942 5000 11994
rect 4704 11940 4760 11942
rect 4784 11940 4840 11942
rect 4864 11940 4920 11942
rect 4944 11940 5000 11942
rect 4704 10906 4760 10908
rect 4784 10906 4840 10908
rect 4864 10906 4920 10908
rect 4944 10906 5000 10908
rect 4704 10854 4750 10906
rect 4750 10854 4760 10906
rect 4784 10854 4814 10906
rect 4814 10854 4826 10906
rect 4826 10854 4840 10906
rect 4864 10854 4878 10906
rect 4878 10854 4890 10906
rect 4890 10854 4920 10906
rect 4944 10854 4954 10906
rect 4954 10854 5000 10906
rect 4704 10852 4760 10854
rect 4784 10852 4840 10854
rect 4864 10852 4920 10854
rect 4944 10852 5000 10854
rect 3974 5616 4030 5672
rect 3790 4936 3846 4992
rect 3238 2896 3294 2952
rect 2830 2746 2886 2748
rect 2910 2746 2966 2748
rect 2990 2746 3046 2748
rect 3070 2746 3126 2748
rect 2830 2694 2876 2746
rect 2876 2694 2886 2746
rect 2910 2694 2940 2746
rect 2940 2694 2952 2746
rect 2952 2694 2966 2746
rect 2990 2694 3004 2746
rect 3004 2694 3016 2746
rect 3016 2694 3046 2746
rect 3070 2694 3080 2746
rect 3080 2694 3126 2746
rect 2830 2692 2886 2694
rect 2910 2692 2966 2694
rect 2990 2692 3046 2694
rect 3070 2692 3126 2694
rect 2502 1400 2558 1456
rect 4158 3576 4214 3632
rect 4704 9818 4760 9820
rect 4784 9818 4840 9820
rect 4864 9818 4920 9820
rect 4944 9818 5000 9820
rect 4704 9766 4750 9818
rect 4750 9766 4760 9818
rect 4784 9766 4814 9818
rect 4814 9766 4826 9818
rect 4826 9766 4840 9818
rect 4864 9766 4878 9818
rect 4878 9766 4890 9818
rect 4890 9766 4920 9818
rect 4944 9766 4954 9818
rect 4954 9766 5000 9818
rect 4704 9764 4760 9766
rect 4784 9764 4840 9766
rect 4864 9764 4920 9766
rect 4944 9764 5000 9766
rect 4704 8730 4760 8732
rect 4784 8730 4840 8732
rect 4864 8730 4920 8732
rect 4944 8730 5000 8732
rect 4704 8678 4750 8730
rect 4750 8678 4760 8730
rect 4784 8678 4814 8730
rect 4814 8678 4826 8730
rect 4826 8678 4840 8730
rect 4864 8678 4878 8730
rect 4878 8678 4890 8730
rect 4890 8678 4920 8730
rect 4944 8678 4954 8730
rect 4954 8678 5000 8730
rect 4704 8676 4760 8678
rect 4784 8676 4840 8678
rect 4864 8676 4920 8678
rect 4944 8676 5000 8678
rect 4704 7642 4760 7644
rect 4784 7642 4840 7644
rect 4864 7642 4920 7644
rect 4944 7642 5000 7644
rect 4704 7590 4750 7642
rect 4750 7590 4760 7642
rect 4784 7590 4814 7642
rect 4814 7590 4826 7642
rect 4826 7590 4840 7642
rect 4864 7590 4878 7642
rect 4878 7590 4890 7642
rect 4890 7590 4920 7642
rect 4944 7590 4954 7642
rect 4954 7590 5000 7642
rect 4704 7588 4760 7590
rect 4784 7588 4840 7590
rect 4864 7588 4920 7590
rect 4944 7588 5000 7590
rect 4704 6554 4760 6556
rect 4784 6554 4840 6556
rect 4864 6554 4920 6556
rect 4944 6554 5000 6556
rect 4704 6502 4750 6554
rect 4750 6502 4760 6554
rect 4784 6502 4814 6554
rect 4814 6502 4826 6554
rect 4826 6502 4840 6554
rect 4864 6502 4878 6554
rect 4878 6502 4890 6554
rect 4890 6502 4920 6554
rect 4944 6502 4954 6554
rect 4954 6502 5000 6554
rect 4704 6500 4760 6502
rect 4784 6500 4840 6502
rect 4864 6500 4920 6502
rect 4944 6500 5000 6502
rect 6182 15136 6238 15192
rect 6578 16890 6634 16892
rect 6658 16890 6714 16892
rect 6738 16890 6794 16892
rect 6818 16890 6874 16892
rect 6578 16838 6624 16890
rect 6624 16838 6634 16890
rect 6658 16838 6688 16890
rect 6688 16838 6700 16890
rect 6700 16838 6714 16890
rect 6738 16838 6752 16890
rect 6752 16838 6764 16890
rect 6764 16838 6794 16890
rect 6818 16838 6828 16890
rect 6828 16838 6874 16890
rect 6578 16836 6634 16838
rect 6658 16836 6714 16838
rect 6738 16836 6794 16838
rect 6818 16836 6874 16838
rect 7102 16632 7158 16688
rect 6578 15802 6634 15804
rect 6658 15802 6714 15804
rect 6738 15802 6794 15804
rect 6818 15802 6874 15804
rect 6578 15750 6624 15802
rect 6624 15750 6634 15802
rect 6658 15750 6688 15802
rect 6688 15750 6700 15802
rect 6700 15750 6714 15802
rect 6738 15750 6752 15802
rect 6752 15750 6764 15802
rect 6764 15750 6794 15802
rect 6818 15750 6828 15802
rect 6828 15750 6874 15802
rect 6578 15748 6634 15750
rect 6658 15748 6714 15750
rect 6738 15748 6794 15750
rect 6818 15748 6874 15750
rect 6918 15000 6974 15056
rect 6578 14714 6634 14716
rect 6658 14714 6714 14716
rect 6738 14714 6794 14716
rect 6818 14714 6874 14716
rect 6578 14662 6624 14714
rect 6624 14662 6634 14714
rect 6658 14662 6688 14714
rect 6688 14662 6700 14714
rect 6700 14662 6714 14714
rect 6738 14662 6752 14714
rect 6752 14662 6764 14714
rect 6764 14662 6794 14714
rect 6818 14662 6828 14714
rect 6828 14662 6874 14714
rect 6578 14660 6634 14662
rect 6658 14660 6714 14662
rect 6738 14660 6794 14662
rect 6818 14660 6874 14662
rect 6578 13626 6634 13628
rect 6658 13626 6714 13628
rect 6738 13626 6794 13628
rect 6818 13626 6874 13628
rect 6578 13574 6624 13626
rect 6624 13574 6634 13626
rect 6658 13574 6688 13626
rect 6688 13574 6700 13626
rect 6700 13574 6714 13626
rect 6738 13574 6752 13626
rect 6752 13574 6764 13626
rect 6764 13574 6794 13626
rect 6818 13574 6828 13626
rect 6828 13574 6874 13626
rect 6578 13572 6634 13574
rect 6658 13572 6714 13574
rect 6738 13572 6794 13574
rect 6818 13572 6874 13574
rect 6578 12538 6634 12540
rect 6658 12538 6714 12540
rect 6738 12538 6794 12540
rect 6818 12538 6874 12540
rect 6578 12486 6624 12538
rect 6624 12486 6634 12538
rect 6658 12486 6688 12538
rect 6688 12486 6700 12538
rect 6700 12486 6714 12538
rect 6738 12486 6752 12538
rect 6752 12486 6764 12538
rect 6764 12486 6794 12538
rect 6818 12486 6828 12538
rect 6828 12486 6874 12538
rect 6578 12484 6634 12486
rect 6658 12484 6714 12486
rect 6738 12484 6794 12486
rect 6818 12484 6874 12486
rect 6578 11450 6634 11452
rect 6658 11450 6714 11452
rect 6738 11450 6794 11452
rect 6818 11450 6874 11452
rect 6578 11398 6624 11450
rect 6624 11398 6634 11450
rect 6658 11398 6688 11450
rect 6688 11398 6700 11450
rect 6700 11398 6714 11450
rect 6738 11398 6752 11450
rect 6752 11398 6764 11450
rect 6764 11398 6794 11450
rect 6818 11398 6828 11450
rect 6828 11398 6874 11450
rect 6578 11396 6634 11398
rect 6658 11396 6714 11398
rect 6738 11396 6794 11398
rect 6818 11396 6874 11398
rect 8452 17434 8508 17436
rect 8532 17434 8588 17436
rect 8612 17434 8668 17436
rect 8692 17434 8748 17436
rect 8452 17382 8498 17434
rect 8498 17382 8508 17434
rect 8532 17382 8562 17434
rect 8562 17382 8574 17434
rect 8574 17382 8588 17434
rect 8612 17382 8626 17434
rect 8626 17382 8638 17434
rect 8638 17382 8668 17434
rect 8692 17382 8702 17434
rect 8702 17382 8748 17434
rect 8452 17380 8508 17382
rect 8532 17380 8588 17382
rect 8612 17380 8668 17382
rect 8692 17380 8748 17382
rect 7562 16632 7618 16688
rect 7746 16496 7802 16552
rect 7194 14320 7250 14376
rect 7194 13912 7250 13968
rect 6578 10362 6634 10364
rect 6658 10362 6714 10364
rect 6738 10362 6794 10364
rect 6818 10362 6874 10364
rect 6578 10310 6624 10362
rect 6624 10310 6634 10362
rect 6658 10310 6688 10362
rect 6688 10310 6700 10362
rect 6700 10310 6714 10362
rect 6738 10310 6752 10362
rect 6752 10310 6764 10362
rect 6764 10310 6794 10362
rect 6818 10310 6828 10362
rect 6828 10310 6874 10362
rect 6578 10308 6634 10310
rect 6658 10308 6714 10310
rect 6738 10308 6794 10310
rect 6818 10308 6874 10310
rect 7654 15816 7710 15872
rect 8206 15136 8262 15192
rect 7746 14592 7802 14648
rect 8942 17176 8998 17232
rect 9310 16768 9366 16824
rect 9126 16532 9128 16552
rect 9128 16532 9180 16552
rect 9180 16532 9182 16552
rect 9126 16496 9182 16532
rect 8452 16346 8508 16348
rect 8532 16346 8588 16348
rect 8612 16346 8668 16348
rect 8692 16346 8748 16348
rect 8452 16294 8498 16346
rect 8498 16294 8508 16346
rect 8532 16294 8562 16346
rect 8562 16294 8574 16346
rect 8574 16294 8588 16346
rect 8612 16294 8626 16346
rect 8626 16294 8638 16346
rect 8638 16294 8668 16346
rect 8692 16294 8702 16346
rect 8702 16294 8748 16346
rect 8452 16292 8508 16294
rect 8532 16292 8588 16294
rect 8612 16292 8668 16294
rect 8692 16292 8748 16294
rect 8452 15258 8508 15260
rect 8532 15258 8588 15260
rect 8612 15258 8668 15260
rect 8692 15258 8748 15260
rect 8452 15206 8498 15258
rect 8498 15206 8508 15258
rect 8532 15206 8562 15258
rect 8562 15206 8574 15258
rect 8574 15206 8588 15258
rect 8612 15206 8626 15258
rect 8626 15206 8638 15258
rect 8638 15206 8668 15258
rect 8692 15206 8702 15258
rect 8702 15206 8748 15258
rect 8452 15204 8508 15206
rect 8532 15204 8588 15206
rect 8612 15204 8668 15206
rect 8692 15204 8748 15206
rect 8574 14764 8576 14784
rect 8576 14764 8628 14784
rect 8628 14764 8630 14784
rect 8574 14728 8630 14764
rect 8574 14592 8630 14648
rect 8850 15000 8906 15056
rect 6578 9274 6634 9276
rect 6658 9274 6714 9276
rect 6738 9274 6794 9276
rect 6818 9274 6874 9276
rect 6578 9222 6624 9274
rect 6624 9222 6634 9274
rect 6658 9222 6688 9274
rect 6688 9222 6700 9274
rect 6700 9222 6714 9274
rect 6738 9222 6752 9274
rect 6752 9222 6764 9274
rect 6764 9222 6794 9274
rect 6818 9222 6828 9274
rect 6828 9222 6874 9274
rect 6578 9220 6634 9222
rect 6658 9220 6714 9222
rect 6738 9220 6794 9222
rect 6818 9220 6874 9222
rect 5078 5752 5134 5808
rect 4704 5466 4760 5468
rect 4784 5466 4840 5468
rect 4864 5466 4920 5468
rect 4944 5466 5000 5468
rect 4704 5414 4750 5466
rect 4750 5414 4760 5466
rect 4784 5414 4814 5466
rect 4814 5414 4826 5466
rect 4826 5414 4840 5466
rect 4864 5414 4878 5466
rect 4878 5414 4890 5466
rect 4890 5414 4920 5466
rect 4944 5414 4954 5466
rect 4954 5414 5000 5466
rect 4704 5412 4760 5414
rect 4784 5412 4840 5414
rect 4864 5412 4920 5414
rect 4944 5412 5000 5414
rect 4066 3476 4068 3496
rect 4068 3476 4120 3496
rect 4120 3476 4122 3496
rect 4066 3440 4122 3476
rect 4434 3576 4490 3632
rect 4802 4528 4858 4584
rect 4704 4378 4760 4380
rect 4784 4378 4840 4380
rect 4864 4378 4920 4380
rect 4944 4378 5000 4380
rect 4704 4326 4750 4378
rect 4750 4326 4760 4378
rect 4784 4326 4814 4378
rect 4814 4326 4826 4378
rect 4826 4326 4840 4378
rect 4864 4326 4878 4378
rect 4878 4326 4890 4378
rect 4890 4326 4920 4378
rect 4944 4326 4954 4378
rect 4954 4326 5000 4378
rect 4704 4324 4760 4326
rect 4784 4324 4840 4326
rect 4864 4324 4920 4326
rect 4944 4324 5000 4326
rect 4704 3290 4760 3292
rect 4784 3290 4840 3292
rect 4864 3290 4920 3292
rect 4944 3290 5000 3292
rect 4704 3238 4750 3290
rect 4750 3238 4760 3290
rect 4784 3238 4814 3290
rect 4814 3238 4826 3290
rect 4826 3238 4840 3290
rect 4864 3238 4878 3290
rect 4878 3238 4890 3290
rect 4890 3238 4920 3290
rect 4944 3238 4954 3290
rect 4954 3238 5000 3290
rect 4704 3236 4760 3238
rect 4784 3236 4840 3238
rect 4864 3236 4920 3238
rect 4944 3236 5000 3238
rect 6578 8186 6634 8188
rect 6658 8186 6714 8188
rect 6738 8186 6794 8188
rect 6818 8186 6874 8188
rect 6578 8134 6624 8186
rect 6624 8134 6634 8186
rect 6658 8134 6688 8186
rect 6688 8134 6700 8186
rect 6700 8134 6714 8186
rect 6738 8134 6752 8186
rect 6752 8134 6764 8186
rect 6764 8134 6794 8186
rect 6818 8134 6828 8186
rect 6828 8134 6874 8186
rect 6578 8132 6634 8134
rect 6658 8132 6714 8134
rect 6738 8132 6794 8134
rect 6818 8132 6874 8134
rect 7286 7248 7342 7304
rect 6578 7098 6634 7100
rect 6658 7098 6714 7100
rect 6738 7098 6794 7100
rect 6818 7098 6874 7100
rect 6578 7046 6624 7098
rect 6624 7046 6634 7098
rect 6658 7046 6688 7098
rect 6688 7046 6700 7098
rect 6700 7046 6714 7098
rect 6738 7046 6752 7098
rect 6752 7046 6764 7098
rect 6764 7046 6794 7098
rect 6818 7046 6828 7098
rect 6828 7046 6874 7098
rect 6578 7044 6634 7046
rect 6658 7044 6714 7046
rect 6738 7044 6794 7046
rect 6818 7044 6874 7046
rect 5630 4664 5686 4720
rect 5446 4392 5502 4448
rect 5446 3984 5502 4040
rect 5538 3576 5594 3632
rect 5538 3340 5540 3360
rect 5540 3340 5592 3360
rect 5592 3340 5594 3360
rect 5538 3304 5594 3340
rect 6366 6160 6422 6216
rect 6090 4936 6146 4992
rect 6090 3304 6146 3360
rect 3606 2372 3662 2408
rect 3606 2352 3608 2372
rect 3608 2352 3660 2372
rect 3660 2352 3662 2372
rect 4704 2202 4760 2204
rect 4784 2202 4840 2204
rect 4864 2202 4920 2204
rect 4944 2202 5000 2204
rect 4704 2150 4750 2202
rect 4750 2150 4760 2202
rect 4784 2150 4814 2202
rect 4814 2150 4826 2202
rect 4826 2150 4840 2202
rect 4864 2150 4878 2202
rect 4878 2150 4890 2202
rect 4890 2150 4920 2202
rect 4944 2150 4954 2202
rect 4954 2150 5000 2202
rect 4704 2148 4760 2150
rect 4784 2148 4840 2150
rect 4864 2148 4920 2150
rect 4944 2148 5000 2150
rect 6578 6010 6634 6012
rect 6658 6010 6714 6012
rect 6738 6010 6794 6012
rect 6818 6010 6874 6012
rect 6578 5958 6624 6010
rect 6624 5958 6634 6010
rect 6658 5958 6688 6010
rect 6688 5958 6700 6010
rect 6700 5958 6714 6010
rect 6738 5958 6752 6010
rect 6752 5958 6764 6010
rect 6764 5958 6794 6010
rect 6818 5958 6828 6010
rect 6828 5958 6874 6010
rect 6578 5956 6634 5958
rect 6658 5956 6714 5958
rect 6738 5956 6794 5958
rect 6818 5956 6874 5958
rect 6578 4922 6634 4924
rect 6658 4922 6714 4924
rect 6738 4922 6794 4924
rect 6818 4922 6874 4924
rect 6578 4870 6624 4922
rect 6624 4870 6634 4922
rect 6658 4870 6688 4922
rect 6688 4870 6700 4922
rect 6700 4870 6714 4922
rect 6738 4870 6752 4922
rect 6752 4870 6764 4922
rect 6764 4870 6794 4922
rect 6818 4870 6828 4922
rect 6828 4870 6874 4922
rect 6578 4868 6634 4870
rect 6658 4868 6714 4870
rect 6738 4868 6794 4870
rect 6818 4868 6874 4870
rect 6826 4528 6882 4584
rect 6578 3834 6634 3836
rect 6658 3834 6714 3836
rect 6738 3834 6794 3836
rect 6818 3834 6874 3836
rect 6578 3782 6624 3834
rect 6624 3782 6634 3834
rect 6658 3782 6688 3834
rect 6688 3782 6700 3834
rect 6700 3782 6714 3834
rect 6738 3782 6752 3834
rect 6752 3782 6764 3834
rect 6764 3782 6794 3834
rect 6818 3782 6828 3834
rect 6828 3782 6874 3834
rect 6578 3780 6634 3782
rect 6658 3780 6714 3782
rect 6738 3780 6794 3782
rect 6818 3780 6874 3782
rect 7746 9424 7802 9480
rect 7562 5888 7618 5944
rect 8452 14170 8508 14172
rect 8532 14170 8588 14172
rect 8612 14170 8668 14172
rect 8692 14170 8748 14172
rect 8452 14118 8498 14170
rect 8498 14118 8508 14170
rect 8532 14118 8562 14170
rect 8562 14118 8574 14170
rect 8574 14118 8588 14170
rect 8612 14118 8626 14170
rect 8626 14118 8638 14170
rect 8638 14118 8668 14170
rect 8692 14118 8702 14170
rect 8702 14118 8748 14170
rect 8452 14116 8508 14118
rect 8532 14116 8588 14118
rect 8612 14116 8668 14118
rect 8692 14116 8748 14118
rect 8452 13082 8508 13084
rect 8532 13082 8588 13084
rect 8612 13082 8668 13084
rect 8692 13082 8748 13084
rect 8452 13030 8498 13082
rect 8498 13030 8508 13082
rect 8532 13030 8562 13082
rect 8562 13030 8574 13082
rect 8574 13030 8588 13082
rect 8612 13030 8626 13082
rect 8626 13030 8638 13082
rect 8638 13030 8668 13082
rect 8692 13030 8702 13082
rect 8702 13030 8748 13082
rect 8452 13028 8508 13030
rect 8532 13028 8588 13030
rect 8612 13028 8668 13030
rect 8692 13028 8748 13030
rect 9402 13776 9458 13832
rect 8452 11994 8508 11996
rect 8532 11994 8588 11996
rect 8612 11994 8668 11996
rect 8692 11994 8748 11996
rect 8452 11942 8498 11994
rect 8498 11942 8508 11994
rect 8532 11942 8562 11994
rect 8562 11942 8574 11994
rect 8574 11942 8588 11994
rect 8612 11942 8626 11994
rect 8626 11942 8638 11994
rect 8638 11942 8668 11994
rect 8692 11942 8702 11994
rect 8702 11942 8748 11994
rect 8452 11940 8508 11942
rect 8532 11940 8588 11942
rect 8612 11940 8668 11942
rect 8692 11940 8748 11942
rect 8452 10906 8508 10908
rect 8532 10906 8588 10908
rect 8612 10906 8668 10908
rect 8692 10906 8748 10908
rect 8452 10854 8498 10906
rect 8498 10854 8508 10906
rect 8532 10854 8562 10906
rect 8562 10854 8574 10906
rect 8574 10854 8588 10906
rect 8612 10854 8626 10906
rect 8626 10854 8638 10906
rect 8638 10854 8668 10906
rect 8692 10854 8702 10906
rect 8702 10854 8748 10906
rect 8452 10852 8508 10854
rect 8532 10852 8588 10854
rect 8612 10852 8668 10854
rect 8692 10852 8748 10854
rect 8452 9818 8508 9820
rect 8532 9818 8588 9820
rect 8612 9818 8668 9820
rect 8692 9818 8748 9820
rect 8452 9766 8498 9818
rect 8498 9766 8508 9818
rect 8532 9766 8562 9818
rect 8562 9766 8574 9818
rect 8574 9766 8588 9818
rect 8612 9766 8626 9818
rect 8626 9766 8638 9818
rect 8638 9766 8668 9818
rect 8692 9766 8702 9818
rect 8702 9766 8748 9818
rect 8452 9764 8508 9766
rect 8532 9764 8588 9766
rect 8612 9764 8668 9766
rect 8692 9764 8748 9766
rect 7378 4800 7434 4856
rect 7286 4256 7342 4312
rect 7102 3576 7158 3632
rect 6578 2746 6634 2748
rect 6658 2746 6714 2748
rect 6738 2746 6794 2748
rect 6818 2746 6874 2748
rect 6578 2694 6624 2746
rect 6624 2694 6634 2746
rect 6658 2694 6688 2746
rect 6688 2694 6700 2746
rect 6700 2694 6714 2746
rect 6738 2694 6752 2746
rect 6752 2694 6764 2746
rect 6764 2694 6794 2746
rect 6818 2694 6828 2746
rect 6828 2694 6874 2746
rect 6578 2692 6634 2694
rect 6658 2692 6714 2694
rect 6738 2692 6794 2694
rect 6818 2692 6874 2694
rect 7194 2760 7250 2816
rect 7746 5344 7802 5400
rect 8022 5344 8078 5400
rect 8452 8730 8508 8732
rect 8532 8730 8588 8732
rect 8612 8730 8668 8732
rect 8692 8730 8748 8732
rect 8452 8678 8498 8730
rect 8498 8678 8508 8730
rect 8532 8678 8562 8730
rect 8562 8678 8574 8730
rect 8574 8678 8588 8730
rect 8612 8678 8626 8730
rect 8626 8678 8638 8730
rect 8638 8678 8668 8730
rect 8692 8678 8702 8730
rect 8702 8678 8748 8730
rect 8452 8676 8508 8678
rect 8532 8676 8588 8678
rect 8612 8676 8668 8678
rect 8692 8676 8748 8678
rect 8452 7642 8508 7644
rect 8532 7642 8588 7644
rect 8612 7642 8668 7644
rect 8692 7642 8748 7644
rect 8452 7590 8498 7642
rect 8498 7590 8508 7642
rect 8532 7590 8562 7642
rect 8562 7590 8574 7642
rect 8574 7590 8588 7642
rect 8612 7590 8626 7642
rect 8626 7590 8638 7642
rect 8638 7590 8668 7642
rect 8692 7590 8702 7642
rect 8702 7590 8748 7642
rect 8452 7588 8508 7590
rect 8532 7588 8588 7590
rect 8612 7588 8668 7590
rect 8692 7588 8748 7590
rect 8452 6554 8508 6556
rect 8532 6554 8588 6556
rect 8612 6554 8668 6556
rect 8692 6554 8748 6556
rect 8452 6502 8498 6554
rect 8498 6502 8508 6554
rect 8532 6502 8562 6554
rect 8562 6502 8574 6554
rect 8574 6502 8588 6554
rect 8612 6502 8626 6554
rect 8626 6502 8638 6554
rect 8638 6502 8668 6554
rect 8692 6502 8702 6554
rect 8702 6502 8748 6554
rect 8452 6500 8508 6502
rect 8532 6500 8588 6502
rect 8612 6500 8668 6502
rect 8692 6500 8748 6502
rect 8452 5466 8508 5468
rect 8532 5466 8588 5468
rect 8612 5466 8668 5468
rect 8692 5466 8748 5468
rect 8452 5414 8498 5466
rect 8498 5414 8508 5466
rect 8532 5414 8562 5466
rect 8562 5414 8574 5466
rect 8574 5414 8588 5466
rect 8612 5414 8626 5466
rect 8626 5414 8638 5466
rect 8638 5414 8668 5466
rect 8692 5414 8702 5466
rect 8702 5414 8748 5466
rect 8452 5412 8508 5414
rect 8532 5412 8588 5414
rect 8612 5412 8668 5414
rect 8692 5412 8748 5414
rect 8114 4800 8170 4856
rect 7930 3340 7932 3360
rect 7932 3340 7984 3360
rect 7984 3340 7986 3360
rect 7930 3304 7986 3340
rect 7746 2896 7802 2952
rect 9678 14592 9734 14648
rect 10046 17176 10102 17232
rect 10326 16890 10382 16892
rect 10406 16890 10462 16892
rect 10486 16890 10542 16892
rect 10566 16890 10622 16892
rect 10326 16838 10372 16890
rect 10372 16838 10382 16890
rect 10406 16838 10436 16890
rect 10436 16838 10448 16890
rect 10448 16838 10462 16890
rect 10486 16838 10500 16890
rect 10500 16838 10512 16890
rect 10512 16838 10542 16890
rect 10566 16838 10576 16890
rect 10576 16838 10622 16890
rect 10326 16836 10382 16838
rect 10406 16836 10462 16838
rect 10486 16836 10542 16838
rect 10566 16836 10622 16838
rect 9954 15988 9956 16008
rect 9956 15988 10008 16008
rect 10008 15988 10010 16008
rect 9954 15952 10010 15988
rect 9862 15680 9918 15736
rect 9862 14320 9918 14376
rect 9954 14220 9956 14240
rect 9956 14220 10008 14240
rect 10008 14220 10010 14240
rect 9954 14184 10010 14220
rect 10690 16360 10746 16416
rect 10690 15952 10746 16008
rect 10326 15802 10382 15804
rect 10406 15802 10462 15804
rect 10486 15802 10542 15804
rect 10566 15802 10622 15804
rect 10326 15750 10372 15802
rect 10372 15750 10382 15802
rect 10406 15750 10436 15802
rect 10436 15750 10448 15802
rect 10448 15750 10462 15802
rect 10486 15750 10500 15802
rect 10500 15750 10512 15802
rect 10512 15750 10542 15802
rect 10566 15750 10576 15802
rect 10576 15750 10622 15802
rect 10326 15748 10382 15750
rect 10406 15748 10462 15750
rect 10486 15748 10542 15750
rect 10566 15748 10622 15750
rect 10326 14714 10382 14716
rect 10406 14714 10462 14716
rect 10486 14714 10542 14716
rect 10566 14714 10622 14716
rect 10326 14662 10372 14714
rect 10372 14662 10382 14714
rect 10406 14662 10436 14714
rect 10436 14662 10448 14714
rect 10448 14662 10462 14714
rect 10486 14662 10500 14714
rect 10500 14662 10512 14714
rect 10512 14662 10542 14714
rect 10566 14662 10576 14714
rect 10576 14662 10622 14714
rect 10326 14660 10382 14662
rect 10406 14660 10462 14662
rect 10486 14660 10542 14662
rect 10566 14660 10622 14662
rect 10782 15136 10838 15192
rect 10782 14728 10838 14784
rect 10326 13626 10382 13628
rect 10406 13626 10462 13628
rect 10486 13626 10542 13628
rect 10566 13626 10622 13628
rect 10326 13574 10372 13626
rect 10372 13574 10382 13626
rect 10406 13574 10436 13626
rect 10436 13574 10448 13626
rect 10448 13574 10462 13626
rect 10486 13574 10500 13626
rect 10500 13574 10512 13626
rect 10512 13574 10542 13626
rect 10566 13574 10576 13626
rect 10576 13574 10622 13626
rect 10326 13572 10382 13574
rect 10406 13572 10462 13574
rect 10486 13572 10542 13574
rect 10566 13572 10622 13574
rect 10598 12980 10654 13016
rect 10598 12960 10600 12980
rect 10600 12960 10652 12980
rect 10652 12960 10654 12980
rect 10326 12538 10382 12540
rect 10406 12538 10462 12540
rect 10486 12538 10542 12540
rect 10566 12538 10622 12540
rect 10326 12486 10372 12538
rect 10372 12486 10382 12538
rect 10406 12486 10436 12538
rect 10436 12486 10448 12538
rect 10448 12486 10462 12538
rect 10486 12486 10500 12538
rect 10500 12486 10512 12538
rect 10512 12486 10542 12538
rect 10566 12486 10576 12538
rect 10576 12486 10622 12538
rect 10326 12484 10382 12486
rect 10406 12484 10462 12486
rect 10486 12484 10542 12486
rect 10566 12484 10622 12486
rect 10326 11450 10382 11452
rect 10406 11450 10462 11452
rect 10486 11450 10542 11452
rect 10566 11450 10622 11452
rect 10326 11398 10372 11450
rect 10372 11398 10382 11450
rect 10406 11398 10436 11450
rect 10436 11398 10448 11450
rect 10448 11398 10462 11450
rect 10486 11398 10500 11450
rect 10500 11398 10512 11450
rect 10512 11398 10542 11450
rect 10566 11398 10576 11450
rect 10576 11398 10622 11450
rect 10326 11396 10382 11398
rect 10406 11396 10462 11398
rect 10486 11396 10542 11398
rect 10566 11396 10622 11398
rect 10782 12552 10838 12608
rect 9126 5888 9182 5944
rect 9218 5752 9274 5808
rect 8452 4378 8508 4380
rect 8532 4378 8588 4380
rect 8612 4378 8668 4380
rect 8692 4378 8748 4380
rect 8452 4326 8498 4378
rect 8498 4326 8508 4378
rect 8532 4326 8562 4378
rect 8562 4326 8574 4378
rect 8574 4326 8588 4378
rect 8612 4326 8626 4378
rect 8626 4326 8638 4378
rect 8638 4326 8668 4378
rect 8692 4326 8702 4378
rect 8702 4326 8748 4378
rect 8452 4324 8508 4326
rect 8532 4324 8588 4326
rect 8612 4324 8668 4326
rect 8692 4324 8748 4326
rect 8452 3290 8508 3292
rect 8532 3290 8588 3292
rect 8612 3290 8668 3292
rect 8692 3290 8748 3292
rect 8452 3238 8498 3290
rect 8498 3238 8508 3290
rect 8532 3238 8562 3290
rect 8562 3238 8574 3290
rect 8574 3238 8588 3290
rect 8612 3238 8626 3290
rect 8626 3238 8638 3290
rect 8638 3238 8668 3290
rect 8692 3238 8702 3290
rect 8702 3238 8748 3290
rect 8452 3236 8508 3238
rect 8532 3236 8588 3238
rect 8612 3236 8668 3238
rect 8692 3236 8748 3238
rect 8452 2202 8508 2204
rect 8532 2202 8588 2204
rect 8612 2202 8668 2204
rect 8692 2202 8748 2204
rect 8452 2150 8498 2202
rect 8498 2150 8508 2202
rect 8532 2150 8562 2202
rect 8562 2150 8574 2202
rect 8574 2150 8588 2202
rect 8612 2150 8626 2202
rect 8626 2150 8638 2202
rect 8638 2150 8668 2202
rect 8692 2150 8702 2202
rect 8702 2150 8748 2202
rect 8452 2148 8508 2150
rect 8532 2148 8588 2150
rect 8612 2148 8668 2150
rect 8692 2148 8748 2150
rect 9402 3712 9458 3768
rect 9862 4800 9918 4856
rect 10138 5344 10194 5400
rect 11150 17040 11206 17096
rect 11150 16632 11206 16688
rect 11150 16088 11206 16144
rect 10966 15036 10968 15056
rect 10968 15036 11020 15056
rect 11020 15036 11022 15056
rect 10966 15000 11022 15036
rect 10966 14048 11022 14104
rect 11150 15136 11206 15192
rect 11426 12724 11428 12744
rect 11428 12724 11480 12744
rect 11480 12724 11482 12744
rect 11426 12688 11482 12724
rect 11794 16632 11850 16688
rect 12200 17434 12256 17436
rect 12280 17434 12336 17436
rect 12360 17434 12416 17436
rect 12440 17434 12496 17436
rect 12200 17382 12246 17434
rect 12246 17382 12256 17434
rect 12280 17382 12310 17434
rect 12310 17382 12322 17434
rect 12322 17382 12336 17434
rect 12360 17382 12374 17434
rect 12374 17382 12386 17434
rect 12386 17382 12416 17434
rect 12440 17382 12450 17434
rect 12450 17382 12496 17434
rect 12200 17380 12256 17382
rect 12280 17380 12336 17382
rect 12360 17380 12416 17382
rect 12440 17380 12496 17382
rect 12714 16904 12770 16960
rect 12714 16652 12770 16688
rect 12714 16632 12716 16652
rect 12716 16632 12768 16652
rect 12768 16632 12770 16652
rect 12200 16346 12256 16348
rect 12280 16346 12336 16348
rect 12360 16346 12416 16348
rect 12440 16346 12496 16348
rect 12200 16294 12246 16346
rect 12246 16294 12256 16346
rect 12280 16294 12310 16346
rect 12310 16294 12322 16346
rect 12322 16294 12336 16346
rect 12360 16294 12374 16346
rect 12374 16294 12386 16346
rect 12386 16294 12416 16346
rect 12440 16294 12450 16346
rect 12450 16294 12496 16346
rect 12200 16292 12256 16294
rect 12280 16292 12336 16294
rect 12360 16292 12416 16294
rect 12440 16292 12496 16294
rect 11794 15136 11850 15192
rect 11794 14900 11796 14920
rect 11796 14900 11848 14920
rect 11848 14900 11850 14920
rect 11794 14864 11850 14900
rect 12200 15258 12256 15260
rect 12280 15258 12336 15260
rect 12360 15258 12416 15260
rect 12440 15258 12496 15260
rect 12200 15206 12246 15258
rect 12246 15206 12256 15258
rect 12280 15206 12310 15258
rect 12310 15206 12322 15258
rect 12322 15206 12336 15258
rect 12360 15206 12374 15258
rect 12374 15206 12386 15258
rect 12386 15206 12416 15258
rect 12440 15206 12450 15258
rect 12450 15206 12496 15258
rect 12200 15204 12256 15206
rect 12280 15204 12336 15206
rect 12360 15204 12416 15206
rect 12440 15204 12496 15206
rect 12200 14170 12256 14172
rect 12280 14170 12336 14172
rect 12360 14170 12416 14172
rect 12440 14170 12496 14172
rect 12200 14118 12246 14170
rect 12246 14118 12256 14170
rect 12280 14118 12310 14170
rect 12310 14118 12322 14170
rect 12322 14118 12336 14170
rect 12360 14118 12374 14170
rect 12374 14118 12386 14170
rect 12386 14118 12416 14170
rect 12440 14118 12450 14170
rect 12450 14118 12496 14170
rect 12200 14116 12256 14118
rect 12280 14116 12336 14118
rect 12360 14116 12416 14118
rect 12440 14116 12496 14118
rect 12200 13082 12256 13084
rect 12280 13082 12336 13084
rect 12360 13082 12416 13084
rect 12440 13082 12496 13084
rect 12200 13030 12246 13082
rect 12246 13030 12256 13082
rect 12280 13030 12310 13082
rect 12310 13030 12322 13082
rect 12322 13030 12336 13082
rect 12360 13030 12374 13082
rect 12374 13030 12386 13082
rect 12386 13030 12416 13082
rect 12440 13030 12450 13082
rect 12450 13030 12496 13082
rect 12200 13028 12256 13030
rect 12280 13028 12336 13030
rect 12360 13028 12416 13030
rect 12440 13028 12496 13030
rect 12806 15308 12808 15328
rect 12808 15308 12860 15328
rect 12860 15308 12862 15328
rect 12806 15272 12862 15308
rect 13450 17040 13506 17096
rect 13358 16768 13414 16824
rect 12714 12824 12770 12880
rect 12200 11994 12256 11996
rect 12280 11994 12336 11996
rect 12360 11994 12416 11996
rect 12440 11994 12496 11996
rect 12200 11942 12246 11994
rect 12246 11942 12256 11994
rect 12280 11942 12310 11994
rect 12310 11942 12322 11994
rect 12322 11942 12336 11994
rect 12360 11942 12374 11994
rect 12374 11942 12386 11994
rect 12386 11942 12416 11994
rect 12440 11942 12450 11994
rect 12450 11942 12496 11994
rect 12200 11940 12256 11942
rect 12280 11940 12336 11942
rect 12360 11940 12416 11942
rect 12440 11940 12496 11942
rect 10326 10362 10382 10364
rect 10406 10362 10462 10364
rect 10486 10362 10542 10364
rect 10566 10362 10622 10364
rect 10326 10310 10372 10362
rect 10372 10310 10382 10362
rect 10406 10310 10436 10362
rect 10436 10310 10448 10362
rect 10448 10310 10462 10362
rect 10486 10310 10500 10362
rect 10500 10310 10512 10362
rect 10512 10310 10542 10362
rect 10566 10310 10576 10362
rect 10576 10310 10622 10362
rect 10326 10308 10382 10310
rect 10406 10308 10462 10310
rect 10486 10308 10542 10310
rect 10566 10308 10622 10310
rect 10326 9274 10382 9276
rect 10406 9274 10462 9276
rect 10486 9274 10542 9276
rect 10566 9274 10622 9276
rect 10326 9222 10372 9274
rect 10372 9222 10382 9274
rect 10406 9222 10436 9274
rect 10436 9222 10448 9274
rect 10448 9222 10462 9274
rect 10486 9222 10500 9274
rect 10500 9222 10512 9274
rect 10512 9222 10542 9274
rect 10566 9222 10576 9274
rect 10576 9222 10622 9274
rect 10326 9220 10382 9222
rect 10406 9220 10462 9222
rect 10486 9220 10542 9222
rect 10566 9220 10622 9222
rect 10326 8186 10382 8188
rect 10406 8186 10462 8188
rect 10486 8186 10542 8188
rect 10566 8186 10622 8188
rect 10326 8134 10372 8186
rect 10372 8134 10382 8186
rect 10406 8134 10436 8186
rect 10436 8134 10448 8186
rect 10448 8134 10462 8186
rect 10486 8134 10500 8186
rect 10500 8134 10512 8186
rect 10512 8134 10542 8186
rect 10566 8134 10576 8186
rect 10576 8134 10622 8186
rect 10326 8132 10382 8134
rect 10406 8132 10462 8134
rect 10486 8132 10542 8134
rect 10566 8132 10622 8134
rect 10326 7098 10382 7100
rect 10406 7098 10462 7100
rect 10486 7098 10542 7100
rect 10566 7098 10622 7100
rect 10326 7046 10372 7098
rect 10372 7046 10382 7098
rect 10406 7046 10436 7098
rect 10436 7046 10448 7098
rect 10448 7046 10462 7098
rect 10486 7046 10500 7098
rect 10500 7046 10512 7098
rect 10512 7046 10542 7098
rect 10566 7046 10576 7098
rect 10576 7046 10622 7098
rect 10326 7044 10382 7046
rect 10406 7044 10462 7046
rect 10486 7044 10542 7046
rect 10566 7044 10622 7046
rect 10326 6010 10382 6012
rect 10406 6010 10462 6012
rect 10486 6010 10542 6012
rect 10566 6010 10622 6012
rect 10326 5958 10372 6010
rect 10372 5958 10382 6010
rect 10406 5958 10436 6010
rect 10436 5958 10448 6010
rect 10448 5958 10462 6010
rect 10486 5958 10500 6010
rect 10500 5958 10512 6010
rect 10512 5958 10542 6010
rect 10566 5958 10576 6010
rect 10576 5958 10622 6010
rect 10326 5956 10382 5958
rect 10406 5956 10462 5958
rect 10486 5956 10542 5958
rect 10566 5956 10622 5958
rect 12200 10906 12256 10908
rect 12280 10906 12336 10908
rect 12360 10906 12416 10908
rect 12440 10906 12496 10908
rect 12200 10854 12246 10906
rect 12246 10854 12256 10906
rect 12280 10854 12310 10906
rect 12310 10854 12322 10906
rect 12322 10854 12336 10906
rect 12360 10854 12374 10906
rect 12374 10854 12386 10906
rect 12386 10854 12416 10906
rect 12440 10854 12450 10906
rect 12450 10854 12496 10906
rect 12200 10852 12256 10854
rect 12280 10852 12336 10854
rect 12360 10852 12416 10854
rect 12440 10852 12496 10854
rect 12200 9818 12256 9820
rect 12280 9818 12336 9820
rect 12360 9818 12416 9820
rect 12440 9818 12496 9820
rect 12200 9766 12246 9818
rect 12246 9766 12256 9818
rect 12280 9766 12310 9818
rect 12310 9766 12322 9818
rect 12322 9766 12336 9818
rect 12360 9766 12374 9818
rect 12374 9766 12386 9818
rect 12386 9766 12416 9818
rect 12440 9766 12450 9818
rect 12450 9766 12496 9818
rect 12200 9764 12256 9766
rect 12280 9764 12336 9766
rect 12360 9764 12416 9766
rect 12440 9764 12496 9766
rect 12714 9016 12770 9072
rect 12200 8730 12256 8732
rect 12280 8730 12336 8732
rect 12360 8730 12416 8732
rect 12440 8730 12496 8732
rect 12200 8678 12246 8730
rect 12246 8678 12256 8730
rect 12280 8678 12310 8730
rect 12310 8678 12322 8730
rect 12322 8678 12336 8730
rect 12360 8678 12374 8730
rect 12374 8678 12386 8730
rect 12386 8678 12416 8730
rect 12440 8678 12450 8730
rect 12450 8678 12496 8730
rect 12200 8676 12256 8678
rect 12280 8676 12336 8678
rect 12360 8676 12416 8678
rect 12440 8676 12496 8678
rect 13174 14320 13230 14376
rect 13450 16652 13506 16688
rect 13450 16632 13452 16652
rect 13452 16632 13504 16652
rect 13504 16632 13506 16652
rect 13174 11892 13230 11928
rect 13174 11872 13176 11892
rect 13176 11872 13228 11892
rect 13228 11872 13230 11892
rect 13818 15408 13874 15464
rect 14370 17076 14372 17096
rect 14372 17076 14424 17096
rect 14424 17076 14426 17096
rect 14370 17040 14426 17076
rect 14074 16890 14130 16892
rect 14154 16890 14210 16892
rect 14234 16890 14290 16892
rect 14314 16890 14370 16892
rect 14074 16838 14120 16890
rect 14120 16838 14130 16890
rect 14154 16838 14184 16890
rect 14184 16838 14196 16890
rect 14196 16838 14210 16890
rect 14234 16838 14248 16890
rect 14248 16838 14260 16890
rect 14260 16838 14290 16890
rect 14314 16838 14324 16890
rect 14324 16838 14370 16890
rect 14074 16836 14130 16838
rect 14154 16836 14210 16838
rect 14234 16836 14290 16838
rect 14314 16836 14370 16838
rect 14074 15802 14130 15804
rect 14154 15802 14210 15804
rect 14234 15802 14290 15804
rect 14314 15802 14370 15804
rect 14074 15750 14120 15802
rect 14120 15750 14130 15802
rect 14154 15750 14184 15802
rect 14184 15750 14196 15802
rect 14196 15750 14210 15802
rect 14234 15750 14248 15802
rect 14248 15750 14260 15802
rect 14260 15750 14290 15802
rect 14314 15750 14324 15802
rect 14324 15750 14370 15802
rect 14074 15748 14130 15750
rect 14154 15748 14210 15750
rect 14234 15748 14290 15750
rect 14314 15748 14370 15750
rect 13542 14864 13598 14920
rect 13726 15000 13782 15056
rect 13174 8880 13230 8936
rect 11702 7792 11758 7848
rect 10966 6332 10968 6352
rect 10968 6332 11020 6352
rect 11020 6332 11022 6352
rect 10966 6296 11022 6332
rect 11426 6704 11482 6760
rect 10322 5516 10324 5536
rect 10324 5516 10376 5536
rect 10376 5516 10378 5536
rect 10322 5480 10378 5516
rect 9862 4004 9918 4040
rect 9862 3984 9864 4004
rect 9864 3984 9916 4004
rect 9916 3984 9918 4004
rect 10046 4120 10102 4176
rect 10326 4922 10382 4924
rect 10406 4922 10462 4924
rect 10486 4922 10542 4924
rect 10566 4922 10622 4924
rect 10326 4870 10372 4922
rect 10372 4870 10382 4922
rect 10406 4870 10436 4922
rect 10436 4870 10448 4922
rect 10448 4870 10462 4922
rect 10486 4870 10500 4922
rect 10500 4870 10512 4922
rect 10512 4870 10542 4922
rect 10566 4870 10576 4922
rect 10576 4870 10622 4922
rect 10326 4868 10382 4870
rect 10406 4868 10462 4870
rect 10486 4868 10542 4870
rect 10566 4868 10622 4870
rect 10506 4528 10562 4584
rect 10326 3834 10382 3836
rect 10406 3834 10462 3836
rect 10486 3834 10542 3836
rect 10566 3834 10622 3836
rect 10326 3782 10372 3834
rect 10372 3782 10382 3834
rect 10406 3782 10436 3834
rect 10436 3782 10448 3834
rect 10448 3782 10462 3834
rect 10486 3782 10500 3834
rect 10500 3782 10512 3834
rect 10512 3782 10542 3834
rect 10566 3782 10576 3834
rect 10576 3782 10622 3834
rect 10326 3780 10382 3782
rect 10406 3780 10462 3782
rect 10486 3780 10542 3782
rect 10566 3780 10622 3782
rect 10230 3440 10286 3496
rect 9954 3168 10010 3224
rect 10322 3032 10378 3088
rect 9862 2760 9918 2816
rect 10326 2746 10382 2748
rect 10406 2746 10462 2748
rect 10486 2746 10542 2748
rect 10566 2746 10622 2748
rect 10326 2694 10372 2746
rect 10372 2694 10382 2746
rect 10406 2694 10436 2746
rect 10436 2694 10448 2746
rect 10448 2694 10462 2746
rect 10486 2694 10500 2746
rect 10500 2694 10512 2746
rect 10512 2694 10542 2746
rect 10566 2694 10576 2746
rect 10576 2694 10622 2746
rect 10326 2692 10382 2694
rect 10406 2692 10462 2694
rect 10486 2692 10542 2694
rect 10566 2692 10622 2694
rect 12200 7642 12256 7644
rect 12280 7642 12336 7644
rect 12360 7642 12416 7644
rect 12440 7642 12496 7644
rect 12200 7590 12246 7642
rect 12246 7590 12256 7642
rect 12280 7590 12310 7642
rect 12310 7590 12322 7642
rect 12322 7590 12336 7642
rect 12360 7590 12374 7642
rect 12374 7590 12386 7642
rect 12386 7590 12416 7642
rect 12440 7590 12450 7642
rect 12450 7590 12496 7642
rect 12200 7588 12256 7590
rect 12280 7588 12336 7590
rect 12360 7588 12416 7590
rect 12440 7588 12496 7590
rect 11150 4392 11206 4448
rect 11242 4256 11298 4312
rect 11242 3712 11298 3768
rect 11334 3188 11390 3224
rect 11334 3168 11336 3188
rect 11336 3168 11388 3188
rect 11388 3168 11390 3188
rect 12200 6554 12256 6556
rect 12280 6554 12336 6556
rect 12360 6554 12416 6556
rect 12440 6554 12496 6556
rect 12200 6502 12246 6554
rect 12246 6502 12256 6554
rect 12280 6502 12310 6554
rect 12310 6502 12322 6554
rect 12322 6502 12336 6554
rect 12360 6502 12374 6554
rect 12374 6502 12386 6554
rect 12386 6502 12416 6554
rect 12440 6502 12450 6554
rect 12450 6502 12496 6554
rect 12200 6500 12256 6502
rect 12280 6500 12336 6502
rect 12360 6500 12416 6502
rect 12440 6500 12496 6502
rect 12346 6316 12402 6352
rect 12346 6296 12348 6316
rect 12348 6296 12400 6316
rect 12400 6296 12402 6316
rect 12714 5752 12770 5808
rect 12200 5466 12256 5468
rect 12280 5466 12336 5468
rect 12360 5466 12416 5468
rect 12440 5466 12496 5468
rect 12200 5414 12246 5466
rect 12246 5414 12256 5466
rect 12280 5414 12310 5466
rect 12310 5414 12322 5466
rect 12322 5414 12336 5466
rect 12360 5414 12374 5466
rect 12374 5414 12386 5466
rect 12386 5414 12416 5466
rect 12440 5414 12450 5466
rect 12450 5414 12496 5466
rect 12200 5412 12256 5414
rect 12280 5412 12336 5414
rect 12360 5412 12416 5414
rect 12440 5412 12496 5414
rect 12070 5208 12126 5264
rect 12254 5244 12256 5264
rect 12256 5244 12308 5264
rect 12308 5244 12310 5264
rect 12254 5208 12310 5244
rect 11978 4936 12034 4992
rect 12070 4528 12126 4584
rect 12200 4378 12256 4380
rect 12280 4378 12336 4380
rect 12360 4378 12416 4380
rect 12440 4378 12496 4380
rect 12200 4326 12246 4378
rect 12246 4326 12256 4378
rect 12280 4326 12310 4378
rect 12310 4326 12322 4378
rect 12322 4326 12336 4378
rect 12360 4326 12374 4378
rect 12374 4326 12386 4378
rect 12386 4326 12416 4378
rect 12440 4326 12450 4378
rect 12450 4326 12496 4378
rect 12200 4324 12256 4326
rect 12280 4324 12336 4326
rect 12360 4324 12416 4326
rect 12440 4324 12496 4326
rect 12346 4020 12348 4040
rect 12348 4020 12400 4040
rect 12400 4020 12402 4040
rect 12346 3984 12402 4020
rect 12200 3290 12256 3292
rect 12280 3290 12336 3292
rect 12360 3290 12416 3292
rect 12440 3290 12496 3292
rect 12200 3238 12246 3290
rect 12246 3238 12256 3290
rect 12280 3238 12310 3290
rect 12310 3238 12322 3290
rect 12322 3238 12336 3290
rect 12360 3238 12374 3290
rect 12374 3238 12386 3290
rect 12386 3238 12416 3290
rect 12440 3238 12450 3290
rect 12450 3238 12496 3290
rect 12200 3236 12256 3238
rect 12280 3236 12336 3238
rect 12360 3236 12416 3238
rect 12440 3236 12496 3238
rect 13818 14728 13874 14784
rect 13818 13948 13820 13968
rect 13820 13948 13872 13968
rect 13872 13948 13874 13968
rect 13818 13912 13874 13948
rect 13726 12044 13728 12064
rect 13728 12044 13780 12064
rect 13780 12044 13782 12064
rect 13726 12008 13782 12044
rect 13818 11892 13874 11928
rect 13818 11872 13820 11892
rect 13820 11872 13872 11892
rect 13872 11872 13874 11892
rect 14646 16652 14702 16688
rect 14646 16632 14648 16652
rect 14648 16632 14700 16652
rect 14700 16632 14702 16652
rect 14074 14714 14130 14716
rect 14154 14714 14210 14716
rect 14234 14714 14290 14716
rect 14314 14714 14370 14716
rect 14074 14662 14120 14714
rect 14120 14662 14130 14714
rect 14154 14662 14184 14714
rect 14184 14662 14196 14714
rect 14196 14662 14210 14714
rect 14234 14662 14248 14714
rect 14248 14662 14260 14714
rect 14260 14662 14290 14714
rect 14314 14662 14324 14714
rect 14324 14662 14370 14714
rect 14074 14660 14130 14662
rect 14154 14660 14210 14662
rect 14234 14660 14290 14662
rect 14314 14660 14370 14662
rect 14278 14456 14334 14512
rect 14278 14220 14280 14240
rect 14280 14220 14332 14240
rect 14332 14220 14334 14240
rect 14278 14184 14334 14220
rect 14074 13626 14130 13628
rect 14154 13626 14210 13628
rect 14234 13626 14290 13628
rect 14314 13626 14370 13628
rect 14074 13574 14120 13626
rect 14120 13574 14130 13626
rect 14154 13574 14184 13626
rect 14184 13574 14196 13626
rect 14196 13574 14210 13626
rect 14234 13574 14248 13626
rect 14248 13574 14260 13626
rect 14260 13574 14290 13626
rect 14314 13574 14324 13626
rect 14324 13574 14370 13626
rect 14074 13572 14130 13574
rect 14154 13572 14210 13574
rect 14234 13572 14290 13574
rect 14314 13572 14370 13574
rect 14094 13232 14150 13288
rect 14074 12538 14130 12540
rect 14154 12538 14210 12540
rect 14234 12538 14290 12540
rect 14314 12538 14370 12540
rect 14074 12486 14120 12538
rect 14120 12486 14130 12538
rect 14154 12486 14184 12538
rect 14184 12486 14196 12538
rect 14196 12486 14210 12538
rect 14234 12486 14248 12538
rect 14248 12486 14260 12538
rect 14260 12486 14290 12538
rect 14314 12486 14324 12538
rect 14324 12486 14370 12538
rect 14074 12484 14130 12486
rect 14154 12484 14210 12486
rect 14234 12484 14290 12486
rect 14314 12484 14370 12486
rect 14370 12280 14426 12336
rect 14554 15308 14556 15328
rect 14556 15308 14608 15328
rect 14608 15308 14610 15328
rect 14554 15272 14610 15308
rect 15658 17856 15714 17912
rect 14738 12980 14794 13016
rect 14738 12960 14740 12980
rect 14740 12960 14792 12980
rect 14792 12960 14794 12980
rect 14074 11450 14130 11452
rect 14154 11450 14210 11452
rect 14234 11450 14290 11452
rect 14314 11450 14370 11452
rect 14074 11398 14120 11450
rect 14120 11398 14130 11450
rect 14154 11398 14184 11450
rect 14184 11398 14196 11450
rect 14196 11398 14210 11450
rect 14234 11398 14248 11450
rect 14248 11398 14260 11450
rect 14260 11398 14290 11450
rect 14314 11398 14324 11450
rect 14324 11398 14370 11450
rect 14074 11396 14130 11398
rect 14154 11396 14210 11398
rect 14234 11396 14290 11398
rect 14314 11396 14370 11398
rect 14074 10362 14130 10364
rect 14154 10362 14210 10364
rect 14234 10362 14290 10364
rect 14314 10362 14370 10364
rect 14074 10310 14120 10362
rect 14120 10310 14130 10362
rect 14154 10310 14184 10362
rect 14184 10310 14196 10362
rect 14196 10310 14210 10362
rect 14234 10310 14248 10362
rect 14248 10310 14260 10362
rect 14260 10310 14290 10362
rect 14314 10310 14324 10362
rect 14324 10310 14370 10362
rect 14074 10308 14130 10310
rect 14154 10308 14210 10310
rect 14234 10308 14290 10310
rect 14314 10308 14370 10310
rect 14554 11076 14610 11112
rect 14554 11056 14556 11076
rect 14556 11056 14608 11076
rect 14608 11056 14610 11076
rect 14074 9274 14130 9276
rect 14154 9274 14210 9276
rect 14234 9274 14290 9276
rect 14314 9274 14370 9276
rect 14074 9222 14120 9274
rect 14120 9222 14130 9274
rect 14154 9222 14184 9274
rect 14184 9222 14196 9274
rect 14196 9222 14210 9274
rect 14234 9222 14248 9274
rect 14248 9222 14260 9274
rect 14260 9222 14290 9274
rect 14314 9222 14324 9274
rect 14324 9222 14370 9274
rect 14074 9220 14130 9222
rect 14154 9220 14210 9222
rect 14234 9220 14290 9222
rect 14314 9220 14370 9222
rect 11978 3032 12034 3088
rect 12200 2202 12256 2204
rect 12280 2202 12336 2204
rect 12360 2202 12416 2204
rect 12440 2202 12496 2204
rect 12200 2150 12246 2202
rect 12246 2150 12256 2202
rect 12280 2150 12310 2202
rect 12310 2150 12322 2202
rect 12322 2150 12336 2202
rect 12360 2150 12374 2202
rect 12374 2150 12386 2202
rect 12386 2150 12416 2202
rect 12440 2150 12450 2202
rect 12450 2150 12496 2202
rect 12200 2148 12256 2150
rect 12280 2148 12336 2150
rect 12360 2148 12416 2150
rect 12440 2148 12496 2150
rect 14074 8186 14130 8188
rect 14154 8186 14210 8188
rect 14234 8186 14290 8188
rect 14314 8186 14370 8188
rect 14074 8134 14120 8186
rect 14120 8134 14130 8186
rect 14154 8134 14184 8186
rect 14184 8134 14196 8186
rect 14196 8134 14210 8186
rect 14234 8134 14248 8186
rect 14248 8134 14260 8186
rect 14260 8134 14290 8186
rect 14314 8134 14324 8186
rect 14324 8134 14370 8186
rect 14074 8132 14130 8134
rect 14154 8132 14210 8134
rect 14234 8132 14290 8134
rect 14314 8132 14370 8134
rect 15106 13096 15162 13152
rect 14074 7098 14130 7100
rect 14154 7098 14210 7100
rect 14234 7098 14290 7100
rect 14314 7098 14370 7100
rect 14074 7046 14120 7098
rect 14120 7046 14130 7098
rect 14154 7046 14184 7098
rect 14184 7046 14196 7098
rect 14196 7046 14210 7098
rect 14234 7046 14248 7098
rect 14248 7046 14260 7098
rect 14260 7046 14290 7098
rect 14314 7046 14324 7098
rect 14324 7046 14370 7098
rect 14074 7044 14130 7046
rect 14154 7044 14210 7046
rect 14234 7044 14290 7046
rect 14314 7044 14370 7046
rect 13726 6180 13782 6216
rect 13726 6160 13728 6180
rect 13728 6160 13780 6180
rect 13780 6160 13782 6180
rect 13726 3848 13782 3904
rect 14094 6160 14150 6216
rect 14074 6010 14130 6012
rect 14154 6010 14210 6012
rect 14234 6010 14290 6012
rect 14314 6010 14370 6012
rect 14074 5958 14120 6010
rect 14120 5958 14130 6010
rect 14154 5958 14184 6010
rect 14184 5958 14196 6010
rect 14196 5958 14210 6010
rect 14234 5958 14248 6010
rect 14248 5958 14260 6010
rect 14260 5958 14290 6010
rect 14314 5958 14324 6010
rect 14324 5958 14370 6010
rect 14074 5956 14130 5958
rect 14154 5956 14210 5958
rect 14234 5956 14290 5958
rect 14314 5956 14370 5958
rect 15014 10004 15016 10024
rect 15016 10004 15068 10024
rect 15068 10004 15070 10024
rect 15014 9968 15070 10004
rect 15014 9696 15070 9752
rect 15566 13912 15622 13968
rect 15566 9968 15622 10024
rect 15750 12416 15806 12472
rect 14646 5752 14702 5808
rect 14094 5072 14150 5128
rect 14074 4922 14130 4924
rect 14154 4922 14210 4924
rect 14234 4922 14290 4924
rect 14314 4922 14370 4924
rect 14074 4870 14120 4922
rect 14120 4870 14130 4922
rect 14154 4870 14184 4922
rect 14184 4870 14196 4922
rect 14196 4870 14210 4922
rect 14234 4870 14248 4922
rect 14248 4870 14260 4922
rect 14260 4870 14290 4922
rect 14314 4870 14324 4922
rect 14324 4870 14370 4922
rect 14074 4868 14130 4870
rect 14154 4868 14210 4870
rect 14234 4868 14290 4870
rect 14314 4868 14370 4870
rect 14462 4428 14464 4448
rect 14464 4428 14516 4448
rect 14516 4428 14518 4448
rect 14462 4392 14518 4428
rect 14074 3834 14130 3836
rect 14154 3834 14210 3836
rect 14234 3834 14290 3836
rect 14314 3834 14370 3836
rect 14074 3782 14120 3834
rect 14120 3782 14130 3834
rect 14154 3782 14184 3834
rect 14184 3782 14196 3834
rect 14196 3782 14210 3834
rect 14234 3782 14248 3834
rect 14248 3782 14260 3834
rect 14260 3782 14290 3834
rect 14314 3782 14324 3834
rect 14324 3782 14370 3834
rect 14074 3780 14130 3782
rect 14154 3780 14210 3782
rect 14234 3780 14290 3782
rect 14314 3780 14370 3782
rect 14370 3440 14426 3496
rect 13818 2916 13874 2952
rect 13818 2896 13820 2916
rect 13820 2896 13872 2916
rect 13872 2896 13874 2916
rect 14094 3052 14150 3088
rect 14094 3032 14096 3052
rect 14096 3032 14148 3052
rect 14148 3032 14150 3052
rect 14074 2746 14130 2748
rect 14154 2746 14210 2748
rect 14234 2746 14290 2748
rect 14314 2746 14370 2748
rect 14074 2694 14120 2746
rect 14120 2694 14130 2746
rect 14154 2694 14184 2746
rect 14184 2694 14196 2746
rect 14196 2694 14210 2746
rect 14234 2694 14248 2746
rect 14248 2694 14260 2746
rect 14260 2694 14290 2746
rect 14314 2694 14324 2746
rect 14324 2694 14370 2746
rect 14074 2692 14130 2694
rect 14154 2692 14210 2694
rect 14234 2692 14290 2694
rect 14314 2692 14370 2694
rect 14370 2488 14426 2544
rect 14922 5888 14978 5944
rect 15106 5480 15162 5536
rect 15014 5344 15070 5400
rect 14830 3984 14886 4040
rect 14646 2080 14702 2136
rect 15290 5208 15346 5264
rect 15566 6060 15568 6080
rect 15568 6060 15620 6080
rect 15620 6060 15622 6080
rect 15566 6024 15622 6060
rect 15566 5652 15568 5672
rect 15568 5652 15620 5672
rect 15620 5652 15622 5672
rect 15566 5616 15622 5652
rect 15382 4120 15438 4176
rect 16394 12416 16450 12472
<< metal3 >>
rect 0 19546 800 19576
rect 0 19486 1410 19546
rect 0 19456 800 19486
rect 1350 19138 1410 19486
rect 2773 19138 2839 19141
rect 1350 19136 2839 19138
rect 1350 19080 2778 19136
rect 2834 19080 2839 19136
rect 1350 19078 2839 19080
rect 2773 19075 2839 19078
rect 0 18594 800 18624
rect 1301 18594 1367 18597
rect 0 18592 1367 18594
rect 0 18536 1306 18592
rect 1362 18536 1367 18592
rect 0 18534 1367 18536
rect 0 18504 800 18534
rect 1301 18531 1367 18534
rect 15653 17914 15719 17917
rect 16400 17914 17200 17944
rect 15653 17912 17200 17914
rect 15653 17856 15658 17912
rect 15714 17856 17200 17912
rect 15653 17854 17200 17856
rect 15653 17851 15719 17854
rect 16400 17824 17200 17854
rect 0 17642 800 17672
rect 2313 17642 2379 17645
rect 0 17640 2379 17642
rect 0 17584 2318 17640
rect 2374 17584 2379 17640
rect 0 17582 2379 17584
rect 0 17552 800 17582
rect 2313 17579 2379 17582
rect 4694 17440 5010 17441
rect 4694 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5010 17440
rect 4694 17375 5010 17376
rect 8442 17440 8758 17441
rect 8442 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8758 17440
rect 8442 17375 8758 17376
rect 12190 17440 12506 17441
rect 12190 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12506 17440
rect 12190 17375 12506 17376
rect 4705 17234 4771 17237
rect 8937 17234 9003 17237
rect 4705 17232 9003 17234
rect 4705 17176 4710 17232
rect 4766 17176 8942 17232
rect 8998 17176 9003 17232
rect 4705 17174 9003 17176
rect 4705 17171 4771 17174
rect 8937 17171 9003 17174
rect 10041 17234 10107 17237
rect 10726 17234 10732 17236
rect 10041 17232 10732 17234
rect 10041 17176 10046 17232
rect 10102 17176 10732 17232
rect 10041 17174 10732 17176
rect 10041 17171 10107 17174
rect 10726 17172 10732 17174
rect 10796 17234 10802 17236
rect 10796 17174 13922 17234
rect 10796 17172 10802 17174
rect 5441 17098 5507 17101
rect 11145 17098 11211 17101
rect 13445 17098 13511 17101
rect 13862 17100 13922 17174
rect 5441 17096 10794 17098
rect 5441 17040 5446 17096
rect 5502 17040 10794 17096
rect 5441 17038 10794 17040
rect 5441 17035 5507 17038
rect 2820 16896 3136 16897
rect 2820 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3136 16896
rect 2820 16831 3136 16832
rect 6568 16896 6884 16897
rect 6568 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6884 16896
rect 6568 16831 6884 16832
rect 10316 16896 10632 16897
rect 10316 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10632 16896
rect 10316 16831 10632 16832
rect 9305 16826 9371 16829
rect 9438 16826 9444 16828
rect 9305 16824 9444 16826
rect 9305 16768 9310 16824
rect 9366 16768 9444 16824
rect 9305 16766 9444 16768
rect 9305 16763 9371 16766
rect 9438 16764 9444 16766
rect 9508 16764 9514 16828
rect 10734 16826 10794 17038
rect 11145 17096 13511 17098
rect 11145 17040 11150 17096
rect 11206 17040 13450 17096
rect 13506 17040 13511 17096
rect 11145 17038 13511 17040
rect 11145 17035 11211 17038
rect 13445 17035 13511 17038
rect 13854 17036 13860 17100
rect 13924 17098 13930 17100
rect 14365 17098 14431 17101
rect 13924 17096 14431 17098
rect 13924 17040 14370 17096
rect 14426 17040 14431 17096
rect 13924 17038 14431 17040
rect 13924 17036 13930 17038
rect 14365 17035 14431 17038
rect 10910 16900 10916 16964
rect 10980 16962 10986 16964
rect 12709 16962 12775 16965
rect 10980 16960 12775 16962
rect 10980 16904 12714 16960
rect 12770 16904 12775 16960
rect 10980 16902 12775 16904
rect 10980 16900 10986 16902
rect 12709 16899 12775 16902
rect 14064 16896 14380 16897
rect 14064 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14380 16896
rect 14064 16831 14380 16832
rect 13353 16826 13419 16829
rect 10734 16824 13419 16826
rect 10734 16768 13358 16824
rect 13414 16768 13419 16824
rect 10734 16766 13419 16768
rect 13353 16763 13419 16766
rect 0 16690 800 16720
rect 1945 16690 2011 16693
rect 0 16688 2011 16690
rect 0 16632 1950 16688
rect 2006 16632 2011 16688
rect 0 16630 2011 16632
rect 0 16600 800 16630
rect 1945 16627 2011 16630
rect 7097 16690 7163 16693
rect 7557 16690 7623 16693
rect 11145 16690 11211 16693
rect 7097 16688 7623 16690
rect 7097 16632 7102 16688
rect 7158 16632 7562 16688
rect 7618 16632 7623 16688
rect 7097 16630 7623 16632
rect 7097 16627 7163 16630
rect 7557 16627 7623 16630
rect 7790 16688 11211 16690
rect 7790 16632 11150 16688
rect 11206 16632 11211 16688
rect 7790 16630 11211 16632
rect 7790 16557 7850 16630
rect 11145 16627 11211 16630
rect 11789 16692 11855 16693
rect 11789 16688 11836 16692
rect 11900 16690 11906 16692
rect 11789 16632 11794 16688
rect 11789 16628 11836 16632
rect 11900 16630 11946 16690
rect 11900 16628 11906 16630
rect 12566 16628 12572 16692
rect 12636 16690 12642 16692
rect 12709 16690 12775 16693
rect 13445 16692 13511 16693
rect 13445 16690 13492 16692
rect 12636 16688 12775 16690
rect 12636 16632 12714 16688
rect 12770 16632 12775 16688
rect 12636 16630 12775 16632
rect 13400 16688 13492 16690
rect 13400 16632 13450 16688
rect 13400 16630 13492 16632
rect 12636 16628 12642 16630
rect 11789 16627 11855 16628
rect 12709 16627 12775 16630
rect 13445 16628 13492 16630
rect 13556 16628 13562 16692
rect 14641 16690 14707 16693
rect 14774 16690 14780 16692
rect 14641 16688 14780 16690
rect 14641 16632 14646 16688
rect 14702 16632 14780 16688
rect 14641 16630 14780 16632
rect 13445 16627 13511 16628
rect 14641 16627 14707 16630
rect 14774 16628 14780 16630
rect 14844 16628 14850 16692
rect 4521 16554 4587 16557
rect 4521 16552 5274 16554
rect 4521 16496 4526 16552
rect 4582 16496 5274 16552
rect 4521 16494 5274 16496
rect 4521 16491 4587 16494
rect 2681 16418 2747 16421
rect 3141 16418 3207 16421
rect 2681 16416 3207 16418
rect 2681 16360 2686 16416
rect 2742 16360 3146 16416
rect 3202 16360 3207 16416
rect 2681 16358 3207 16360
rect 5214 16418 5274 16494
rect 7741 16552 7850 16557
rect 9121 16554 9187 16557
rect 9622 16554 9628 16556
rect 7741 16496 7746 16552
rect 7802 16496 7850 16552
rect 7741 16494 7850 16496
rect 7974 16494 8954 16554
rect 7741 16491 7807 16494
rect 7974 16418 8034 16494
rect 5214 16358 8034 16418
rect 8894 16418 8954 16494
rect 9121 16552 9628 16554
rect 9121 16496 9126 16552
rect 9182 16496 9628 16552
rect 9121 16494 9628 16496
rect 9121 16491 9187 16494
rect 9622 16492 9628 16494
rect 9692 16492 9698 16556
rect 10685 16418 10751 16421
rect 8894 16416 10751 16418
rect 8894 16360 10690 16416
rect 10746 16360 10751 16416
rect 8894 16358 10751 16360
rect 2681 16355 2747 16358
rect 3141 16355 3207 16358
rect 10685 16355 10751 16358
rect 4694 16352 5010 16353
rect 4694 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5010 16352
rect 4694 16287 5010 16288
rect 8442 16352 8758 16353
rect 8442 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8758 16352
rect 8442 16287 8758 16288
rect 12190 16352 12506 16353
rect 12190 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12506 16352
rect 12190 16287 12506 16288
rect 2313 16146 2379 16149
rect 11145 16146 11211 16149
rect 2313 16144 11211 16146
rect 2313 16088 2318 16144
rect 2374 16088 11150 16144
rect 11206 16088 11211 16144
rect 2313 16086 11211 16088
rect 2313 16083 2379 16086
rect 11145 16083 11211 16086
rect 4061 16010 4127 16013
rect 6085 16010 6151 16013
rect 8886 16010 8892 16012
rect 4061 16008 8892 16010
rect 4061 15952 4066 16008
rect 4122 15952 6090 16008
rect 6146 15952 8892 16008
rect 4061 15950 8892 15952
rect 4061 15947 4127 15950
rect 6085 15947 6151 15950
rect 8886 15948 8892 15950
rect 8956 15948 8962 16012
rect 9949 16010 10015 16013
rect 10174 16010 10180 16012
rect 9949 16008 10180 16010
rect 9949 15952 9954 16008
rect 10010 15952 10180 16008
rect 9949 15950 10180 15952
rect 9949 15947 10015 15950
rect 10174 15948 10180 15950
rect 10244 16010 10250 16012
rect 10685 16010 10751 16013
rect 10244 16008 10751 16010
rect 10244 15952 10690 16008
rect 10746 15952 10751 16008
rect 10244 15950 10751 15952
rect 10244 15948 10250 15950
rect 10685 15947 10751 15950
rect 7649 15874 7715 15877
rect 7782 15874 7788 15876
rect 7649 15872 7788 15874
rect 7649 15816 7654 15872
rect 7710 15816 7788 15872
rect 7649 15814 7788 15816
rect 7649 15811 7715 15814
rect 7782 15812 7788 15814
rect 7852 15812 7858 15876
rect 2820 15808 3136 15809
rect 0 15738 800 15768
rect 2820 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3136 15808
rect 2820 15743 3136 15744
rect 6568 15808 6884 15809
rect 6568 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6884 15808
rect 6568 15743 6884 15744
rect 10316 15808 10632 15809
rect 10316 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10632 15808
rect 10316 15743 10632 15744
rect 14064 15808 14380 15809
rect 14064 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14380 15808
rect 14064 15743 14380 15744
rect 1485 15738 1551 15741
rect 4613 15738 4679 15741
rect 0 15736 1551 15738
rect 0 15680 1490 15736
rect 1546 15680 1551 15736
rect 0 15678 1551 15680
rect 0 15648 800 15678
rect 1485 15675 1551 15678
rect 4110 15736 4679 15738
rect 4110 15680 4618 15736
rect 4674 15680 4679 15736
rect 4110 15678 4679 15680
rect 3417 15602 3483 15605
rect 4110 15602 4170 15678
rect 4613 15675 4679 15678
rect 9438 15676 9444 15740
rect 9508 15738 9514 15740
rect 9857 15738 9923 15741
rect 9508 15736 9923 15738
rect 9508 15680 9862 15736
rect 9918 15680 9923 15736
rect 9508 15678 9923 15680
rect 9508 15676 9514 15678
rect 9857 15675 9923 15678
rect 3417 15600 4170 15602
rect 3417 15544 3422 15600
rect 3478 15544 4170 15600
rect 3417 15542 4170 15544
rect 4337 15602 4403 15605
rect 4337 15600 14106 15602
rect 4337 15544 4342 15600
rect 4398 15544 14106 15600
rect 4337 15542 14106 15544
rect 3417 15539 3483 15542
rect 4337 15539 4403 15542
rect 2037 15466 2103 15469
rect 13813 15466 13879 15469
rect 2037 15464 13879 15466
rect 2037 15408 2042 15464
rect 2098 15408 13818 15464
rect 13874 15408 13879 15464
rect 2037 15406 13879 15408
rect 2037 15403 2103 15406
rect 13813 15403 13879 15406
rect 1894 15268 1900 15332
rect 1964 15330 1970 15332
rect 2129 15330 2195 15333
rect 1964 15328 2195 15330
rect 1964 15272 2134 15328
rect 2190 15272 2195 15328
rect 1964 15270 2195 15272
rect 1964 15268 1970 15270
rect 2129 15267 2195 15270
rect 2405 15330 2471 15333
rect 3601 15330 3667 15333
rect 3877 15330 3943 15333
rect 12801 15330 12867 15333
rect 2405 15328 3943 15330
rect 2405 15272 2410 15328
rect 2466 15272 3606 15328
rect 3662 15272 3882 15328
rect 3938 15272 3943 15328
rect 2405 15270 3943 15272
rect 2405 15267 2471 15270
rect 3601 15267 3667 15270
rect 3877 15267 3943 15270
rect 12758 15328 12867 15330
rect 12758 15272 12806 15328
rect 12862 15272 12867 15328
rect 12758 15267 12867 15272
rect 14046 15330 14106 15542
rect 14549 15332 14615 15333
rect 14549 15330 14596 15332
rect 14046 15328 14596 15330
rect 14046 15272 14554 15328
rect 14046 15270 14596 15272
rect 14549 15268 14596 15270
rect 14660 15268 14666 15332
rect 14549 15267 14615 15268
rect 4694 15264 5010 15265
rect 4694 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5010 15264
rect 4694 15199 5010 15200
rect 8442 15264 8758 15265
rect 8442 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8758 15264
rect 8442 15199 8758 15200
rect 12190 15264 12506 15265
rect 12190 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12506 15264
rect 12190 15199 12506 15200
rect 6177 15194 6243 15197
rect 8201 15194 8267 15197
rect 6177 15192 8267 15194
rect 6177 15136 6182 15192
rect 6238 15136 8206 15192
rect 8262 15136 8267 15192
rect 6177 15134 8267 15136
rect 6177 15131 6243 15134
rect 8201 15131 8267 15134
rect 10777 15194 10843 15197
rect 11145 15194 11211 15197
rect 11789 15194 11855 15197
rect 10777 15192 11855 15194
rect 10777 15136 10782 15192
rect 10838 15136 11150 15192
rect 11206 15136 11794 15192
rect 11850 15136 11855 15192
rect 10777 15134 11855 15136
rect 10777 15131 10843 15134
rect 11145 15131 11211 15134
rect 11789 15131 11855 15134
rect 1945 15058 2011 15061
rect 5625 15058 5691 15061
rect 1945 15056 5691 15058
rect 1945 15000 1950 15056
rect 2006 15000 5630 15056
rect 5686 15000 5691 15056
rect 1945 14998 5691 15000
rect 1945 14995 2011 14998
rect 5625 14995 5691 14998
rect 6913 15058 6979 15061
rect 8845 15058 8911 15061
rect 6913 15056 8911 15058
rect 6913 15000 6918 15056
rect 6974 15000 8850 15056
rect 8906 15000 8911 15056
rect 6913 14998 8911 15000
rect 6913 14995 6979 14998
rect 8845 14995 8911 14998
rect 10961 15058 11027 15061
rect 12758 15058 12818 15267
rect 12934 15058 12940 15060
rect 10961 15056 12940 15058
rect 10961 15000 10966 15056
rect 11022 15000 12940 15056
rect 10961 14998 12940 15000
rect 10961 14995 11027 14998
rect 12934 14996 12940 14998
rect 13004 14996 13010 15060
rect 13721 15056 13787 15061
rect 13721 15000 13726 15056
rect 13782 15000 13787 15056
rect 13721 14995 13787 15000
rect 3049 14922 3115 14925
rect 3509 14922 3575 14925
rect 11789 14922 11855 14925
rect 3049 14920 11855 14922
rect 3049 14864 3054 14920
rect 3110 14864 3514 14920
rect 3570 14864 11794 14920
rect 11850 14864 11855 14920
rect 3049 14862 11855 14864
rect 3049 14859 3115 14862
rect 3509 14859 3575 14862
rect 11789 14859 11855 14862
rect 13537 14922 13603 14925
rect 13724 14922 13784 14995
rect 13537 14920 13784 14922
rect 13537 14864 13542 14920
rect 13598 14864 13784 14920
rect 13537 14862 13784 14864
rect 13537 14859 13603 14862
rect 0 14786 800 14816
rect 1485 14786 1551 14789
rect 0 14784 1551 14786
rect 0 14728 1490 14784
rect 1546 14728 1551 14784
rect 0 14726 1551 14728
rect 0 14696 800 14726
rect 1485 14723 1551 14726
rect 7782 14724 7788 14788
rect 7852 14786 7858 14788
rect 8569 14786 8635 14789
rect 7852 14784 8635 14786
rect 7852 14728 8574 14784
rect 8630 14728 8635 14784
rect 7852 14726 8635 14728
rect 7852 14724 7858 14726
rect 8569 14723 8635 14726
rect 10777 14786 10843 14789
rect 13670 14786 13676 14788
rect 10777 14784 13676 14786
rect 10777 14728 10782 14784
rect 10838 14728 13676 14784
rect 10777 14726 13676 14728
rect 10777 14723 10843 14726
rect 13670 14724 13676 14726
rect 13740 14786 13746 14788
rect 13813 14786 13879 14789
rect 13740 14784 13879 14786
rect 13740 14728 13818 14784
rect 13874 14728 13879 14784
rect 13740 14726 13879 14728
rect 13740 14724 13746 14726
rect 13813 14723 13879 14726
rect 2820 14720 3136 14721
rect 2820 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3136 14720
rect 2820 14655 3136 14656
rect 6568 14720 6884 14721
rect 6568 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6884 14720
rect 6568 14655 6884 14656
rect 10316 14720 10632 14721
rect 10316 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10632 14720
rect 10316 14655 10632 14656
rect 14064 14720 14380 14721
rect 14064 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14380 14720
rect 14064 14655 14380 14656
rect 7741 14650 7807 14653
rect 8569 14650 8635 14653
rect 9673 14650 9739 14653
rect 7741 14648 8635 14650
rect 7741 14592 7746 14648
rect 7802 14592 8574 14648
rect 8630 14592 8635 14648
rect 7741 14590 8635 14592
rect 7741 14587 7807 14590
rect 8569 14587 8635 14590
rect 8710 14648 9739 14650
rect 8710 14592 9678 14648
rect 9734 14592 9739 14648
rect 8710 14590 9739 14592
rect 4245 14514 4311 14517
rect 8710 14514 8770 14590
rect 9673 14587 9739 14590
rect 4245 14512 8770 14514
rect 4245 14456 4250 14512
rect 4306 14456 8770 14512
rect 4245 14454 8770 14456
rect 4245 14451 4311 14454
rect 8886 14452 8892 14516
rect 8956 14514 8962 14516
rect 14273 14514 14339 14517
rect 8956 14512 14339 14514
rect 8956 14456 14278 14512
rect 14334 14456 14339 14512
rect 8956 14454 14339 14456
rect 8956 14452 8962 14454
rect 14273 14451 14339 14454
rect 1894 14316 1900 14380
rect 1964 14378 1970 14380
rect 7189 14378 7255 14381
rect 9857 14378 9923 14381
rect 13169 14378 13235 14381
rect 1964 14376 7255 14378
rect 1964 14320 7194 14376
rect 7250 14320 7255 14376
rect 1964 14318 7255 14320
rect 1964 14316 1970 14318
rect 7189 14315 7255 14318
rect 8158 14376 9923 14378
rect 8158 14320 9862 14376
rect 9918 14320 9923 14376
rect 8158 14318 9923 14320
rect 5257 14242 5323 14245
rect 8158 14242 8218 14318
rect 9857 14315 9923 14318
rect 9998 14376 13235 14378
rect 9998 14320 13174 14376
rect 13230 14320 13235 14376
rect 9998 14318 13235 14320
rect 9998 14245 10058 14318
rect 13169 14315 13235 14318
rect 9949 14244 10058 14245
rect 9949 14242 9996 14244
rect 5257 14240 8218 14242
rect 5257 14184 5262 14240
rect 5318 14184 8218 14240
rect 5257 14182 8218 14184
rect 9904 14240 9996 14242
rect 9904 14184 9954 14240
rect 9904 14182 9996 14184
rect 5257 14179 5323 14182
rect 9949 14180 9996 14182
rect 10060 14180 10066 14244
rect 14273 14242 14339 14245
rect 15142 14242 15148 14244
rect 14273 14240 15148 14242
rect 14273 14184 14278 14240
rect 14334 14184 15148 14240
rect 14273 14182 15148 14184
rect 9949 14179 10015 14180
rect 14273 14179 14339 14182
rect 15142 14180 15148 14182
rect 15212 14180 15218 14244
rect 4694 14176 5010 14177
rect 4694 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5010 14176
rect 4694 14111 5010 14112
rect 8442 14176 8758 14177
rect 8442 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8758 14176
rect 8442 14111 8758 14112
rect 12190 14176 12506 14177
rect 12190 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12506 14176
rect 12190 14111 12506 14112
rect 3417 14106 3483 14109
rect 10961 14108 11027 14109
rect 3417 14104 4538 14106
rect 3417 14048 3422 14104
rect 3478 14048 4538 14104
rect 3417 14046 4538 14048
rect 3417 14043 3483 14046
rect 1945 13970 2011 13973
rect 4245 13970 4311 13973
rect 1945 13968 4311 13970
rect 1945 13912 1950 13968
rect 2006 13912 4250 13968
rect 4306 13912 4311 13968
rect 1945 13910 4311 13912
rect 4478 13970 4538 14046
rect 10910 14044 10916 14108
rect 10980 14106 11027 14108
rect 10980 14104 11072 14106
rect 11022 14048 11072 14104
rect 10980 14046 11072 14048
rect 10980 14044 11027 14046
rect 10961 14043 11027 14044
rect 7189 13970 7255 13973
rect 13813 13970 13879 13973
rect 4478 13910 6562 13970
rect 1945 13907 2011 13910
rect 4245 13907 4311 13910
rect 0 13834 800 13864
rect 1485 13834 1551 13837
rect 0 13832 1551 13834
rect 0 13776 1490 13832
rect 1546 13776 1551 13832
rect 0 13774 1551 13776
rect 0 13744 800 13774
rect 1485 13771 1551 13774
rect 3366 13772 3372 13836
rect 3436 13834 3442 13836
rect 4153 13834 4219 13837
rect 3436 13832 4219 13834
rect 3436 13776 4158 13832
rect 4214 13776 4219 13832
rect 3436 13774 4219 13776
rect 6502 13834 6562 13910
rect 7189 13968 13879 13970
rect 7189 13912 7194 13968
rect 7250 13912 13818 13968
rect 13874 13912 13879 13968
rect 7189 13910 13879 13912
rect 7189 13907 7255 13910
rect 13813 13907 13879 13910
rect 15561 13970 15627 13973
rect 16400 13970 17200 14000
rect 15561 13968 17200 13970
rect 15561 13912 15566 13968
rect 15622 13912 17200 13968
rect 15561 13910 17200 13912
rect 15561 13907 15627 13910
rect 16400 13880 17200 13910
rect 9397 13834 9463 13837
rect 6502 13832 9463 13834
rect 6502 13776 9402 13832
rect 9458 13776 9463 13832
rect 6502 13774 9463 13776
rect 3436 13772 3442 13774
rect 4153 13771 4219 13774
rect 9397 13771 9463 13774
rect 2820 13632 3136 13633
rect 2820 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3136 13632
rect 2820 13567 3136 13568
rect 6568 13632 6884 13633
rect 6568 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6884 13632
rect 6568 13567 6884 13568
rect 10316 13632 10632 13633
rect 10316 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10632 13632
rect 10316 13567 10632 13568
rect 14064 13632 14380 13633
rect 14064 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14380 13632
rect 14064 13567 14380 13568
rect 2681 13290 2747 13293
rect 14089 13290 14155 13293
rect 2681 13288 14155 13290
rect 2681 13232 2686 13288
rect 2742 13232 14094 13288
rect 14150 13232 14155 13288
rect 2681 13230 14155 13232
rect 2681 13227 2747 13230
rect 14089 13227 14155 13230
rect 14958 13092 14964 13156
rect 15028 13154 15034 13156
rect 15101 13154 15167 13157
rect 15028 13152 15167 13154
rect 15028 13096 15106 13152
rect 15162 13096 15167 13152
rect 15028 13094 15167 13096
rect 15028 13092 15034 13094
rect 15101 13091 15167 13094
rect 4694 13088 5010 13089
rect 4694 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5010 13088
rect 4694 13023 5010 13024
rect 8442 13088 8758 13089
rect 8442 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8758 13088
rect 8442 13023 8758 13024
rect 12190 13088 12506 13089
rect 12190 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12506 13088
rect 12190 13023 12506 13024
rect 10593 13018 10659 13021
rect 14733 13020 14799 13021
rect 10726 13018 10732 13020
rect 10593 13016 10732 13018
rect 10593 12960 10598 13016
rect 10654 12960 10732 13016
rect 10593 12958 10732 12960
rect 10593 12955 10659 12958
rect 10726 12956 10732 12958
rect 10796 12956 10802 13020
rect 14733 13018 14780 13020
rect 14688 13016 14780 13018
rect 14688 12960 14738 13016
rect 14688 12958 14780 12960
rect 14733 12956 14780 12958
rect 14844 12956 14850 13020
rect 14733 12955 14799 12956
rect 0 12882 800 12912
rect 1485 12882 1551 12885
rect 0 12880 1551 12882
rect 0 12824 1490 12880
rect 1546 12824 1551 12880
rect 0 12822 1551 12824
rect 0 12792 800 12822
rect 1485 12819 1551 12822
rect 12709 12882 12775 12885
rect 13118 12882 13124 12884
rect 12709 12880 13124 12882
rect 12709 12824 12714 12880
rect 12770 12824 13124 12880
rect 12709 12822 13124 12824
rect 12709 12819 12775 12822
rect 13118 12820 13124 12822
rect 13188 12820 13194 12884
rect 9438 12746 9444 12748
rect 6318 12686 9444 12746
rect 3233 12610 3299 12613
rect 6318 12610 6378 12686
rect 9438 12684 9444 12686
rect 9508 12684 9514 12748
rect 11421 12746 11487 12749
rect 12014 12746 12020 12748
rect 11421 12744 12020 12746
rect 11421 12688 11426 12744
rect 11482 12688 12020 12744
rect 11421 12686 12020 12688
rect 11421 12683 11487 12686
rect 12014 12684 12020 12686
rect 12084 12684 12090 12748
rect 10777 12612 10843 12613
rect 3233 12608 6378 12610
rect 3233 12552 3238 12608
rect 3294 12552 6378 12608
rect 3233 12550 6378 12552
rect 3233 12547 3299 12550
rect 10726 12548 10732 12612
rect 10796 12610 10843 12612
rect 10796 12608 10888 12610
rect 10838 12552 10888 12608
rect 10796 12550 10888 12552
rect 10796 12548 10843 12550
rect 10777 12547 10843 12548
rect 2820 12544 3136 12545
rect 2820 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3136 12544
rect 2820 12479 3136 12480
rect 6568 12544 6884 12545
rect 6568 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6884 12544
rect 6568 12479 6884 12480
rect 10316 12544 10632 12545
rect 10316 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10632 12544
rect 10316 12479 10632 12480
rect 14064 12544 14380 12545
rect 14064 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14380 12544
rect 14064 12479 14380 12480
rect 15745 12474 15811 12477
rect 16389 12474 16455 12477
rect 15745 12472 16455 12474
rect 15745 12416 15750 12472
rect 15806 12416 16394 12472
rect 16450 12416 16455 12472
rect 15745 12414 16455 12416
rect 15745 12411 15811 12414
rect 16389 12411 16455 12414
rect 13670 12276 13676 12340
rect 13740 12338 13746 12340
rect 14365 12338 14431 12341
rect 13740 12336 14431 12338
rect 13740 12280 14370 12336
rect 14426 12280 14431 12336
rect 13740 12278 14431 12280
rect 13740 12276 13746 12278
rect 14365 12275 14431 12278
rect 3877 12204 3943 12205
rect 3877 12202 3924 12204
rect 3832 12200 3924 12202
rect 3832 12144 3882 12200
rect 3832 12142 3924 12144
rect 3877 12140 3924 12142
rect 3988 12140 3994 12204
rect 10174 12140 10180 12204
rect 10244 12202 10250 12204
rect 10244 12142 13738 12202
rect 10244 12140 10250 12142
rect 3877 12139 3943 12140
rect 13678 12069 13738 12142
rect 13678 12068 13787 12069
rect 13670 12004 13676 12068
rect 13740 12066 13787 12068
rect 13740 12064 13832 12066
rect 13782 12008 13832 12064
rect 13740 12006 13832 12008
rect 13740 12004 13787 12006
rect 13721 12003 13787 12004
rect 4694 12000 5010 12001
rect 0 11930 800 11960
rect 4694 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5010 12000
rect 4694 11935 5010 11936
rect 8442 12000 8758 12001
rect 8442 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8758 12000
rect 8442 11935 8758 11936
rect 12190 12000 12506 12001
rect 12190 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12506 12000
rect 12190 11935 12506 11936
rect 1485 11930 1551 11933
rect 0 11928 1551 11930
rect 0 11872 1490 11928
rect 1546 11872 1551 11928
rect 0 11870 1551 11872
rect 0 11840 800 11870
rect 1485 11867 1551 11870
rect 12934 11868 12940 11932
rect 13004 11930 13010 11932
rect 13169 11930 13235 11933
rect 13813 11932 13879 11933
rect 13813 11930 13860 11932
rect 13004 11928 13235 11930
rect 13004 11872 13174 11928
rect 13230 11872 13235 11928
rect 13004 11870 13235 11872
rect 13768 11928 13860 11930
rect 13768 11872 13818 11928
rect 13768 11870 13860 11872
rect 13004 11868 13010 11870
rect 13169 11867 13235 11870
rect 13813 11868 13860 11870
rect 13924 11868 13930 11932
rect 13813 11867 13879 11868
rect 2820 11456 3136 11457
rect 2820 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3136 11456
rect 2820 11391 3136 11392
rect 6568 11456 6884 11457
rect 6568 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6884 11456
rect 6568 11391 6884 11392
rect 10316 11456 10632 11457
rect 10316 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10632 11456
rect 10316 11391 10632 11392
rect 14064 11456 14380 11457
rect 14064 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14380 11456
rect 14064 11391 14380 11392
rect 3233 11386 3299 11389
rect 3366 11386 3372 11388
rect 3233 11384 3372 11386
rect 3233 11328 3238 11384
rect 3294 11328 3372 11384
rect 3233 11326 3372 11328
rect 3233 11323 3299 11326
rect 3366 11324 3372 11326
rect 3436 11324 3442 11388
rect 13854 11052 13860 11116
rect 13924 11114 13930 11116
rect 14549 11114 14615 11117
rect 15142 11114 15148 11116
rect 13924 11112 15148 11114
rect 13924 11056 14554 11112
rect 14610 11056 15148 11112
rect 13924 11054 15148 11056
rect 13924 11052 13930 11054
rect 14549 11051 14615 11054
rect 15142 11052 15148 11054
rect 15212 11052 15218 11116
rect 0 10978 800 11008
rect 1485 10978 1551 10981
rect 0 10976 1551 10978
rect 0 10920 1490 10976
rect 1546 10920 1551 10976
rect 0 10918 1551 10920
rect 0 10888 800 10918
rect 1485 10915 1551 10918
rect 4694 10912 5010 10913
rect 4694 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5010 10912
rect 4694 10847 5010 10848
rect 8442 10912 8758 10913
rect 8442 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8758 10912
rect 8442 10847 8758 10848
rect 12190 10912 12506 10913
rect 12190 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12506 10912
rect 12190 10847 12506 10848
rect 2820 10368 3136 10369
rect 2820 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3136 10368
rect 2820 10303 3136 10304
rect 6568 10368 6884 10369
rect 6568 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6884 10368
rect 6568 10303 6884 10304
rect 10316 10368 10632 10369
rect 10316 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10632 10368
rect 10316 10303 10632 10304
rect 14064 10368 14380 10369
rect 14064 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14380 10368
rect 14064 10303 14380 10304
rect 0 10026 800 10056
rect 1485 10026 1551 10029
rect 0 10024 1551 10026
rect 0 9968 1490 10024
rect 1546 9968 1551 10024
rect 0 9966 1551 9968
rect 0 9936 800 9966
rect 1485 9963 1551 9966
rect 11278 9964 11284 10028
rect 11348 10026 11354 10028
rect 15009 10026 15075 10029
rect 11348 10024 15075 10026
rect 11348 9968 15014 10024
rect 15070 9968 15075 10024
rect 11348 9966 15075 9968
rect 11348 9964 11354 9966
rect 15009 9963 15075 9966
rect 15561 10026 15627 10029
rect 16400 10026 17200 10056
rect 15561 10024 17200 10026
rect 15561 9968 15566 10024
rect 15622 9968 17200 10024
rect 15561 9966 17200 9968
rect 15561 9963 15627 9966
rect 16400 9936 17200 9966
rect 4694 9824 5010 9825
rect 4694 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5010 9824
rect 4694 9759 5010 9760
rect 8442 9824 8758 9825
rect 8442 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8758 9824
rect 8442 9759 8758 9760
rect 12190 9824 12506 9825
rect 12190 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12506 9824
rect 12190 9759 12506 9760
rect 13486 9692 13492 9756
rect 13556 9754 13562 9756
rect 15009 9754 15075 9757
rect 13556 9752 15075 9754
rect 13556 9696 15014 9752
rect 15070 9696 15075 9752
rect 13556 9694 15075 9696
rect 13556 9692 13562 9694
rect 15009 9691 15075 9694
rect 1577 9618 1643 9621
rect 3366 9618 3372 9620
rect 1577 9616 3372 9618
rect 1577 9560 1582 9616
rect 1638 9560 3372 9616
rect 1577 9558 3372 9560
rect 1577 9555 1643 9558
rect 3366 9556 3372 9558
rect 3436 9556 3442 9620
rect 7741 9482 7807 9485
rect 13854 9482 13860 9484
rect 7741 9480 13860 9482
rect 7741 9424 7746 9480
rect 7802 9424 13860 9480
rect 7741 9422 13860 9424
rect 7741 9419 7807 9422
rect 13854 9420 13860 9422
rect 13924 9420 13930 9484
rect 2820 9280 3136 9281
rect 2820 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3136 9280
rect 2820 9215 3136 9216
rect 6568 9280 6884 9281
rect 6568 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6884 9280
rect 6568 9215 6884 9216
rect 10316 9280 10632 9281
rect 10316 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10632 9280
rect 10316 9215 10632 9216
rect 14064 9280 14380 9281
rect 14064 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14380 9280
rect 14064 9215 14380 9216
rect 0 9074 800 9104
rect 1485 9074 1551 9077
rect 0 9072 1551 9074
rect 0 9016 1490 9072
rect 1546 9016 1551 9072
rect 0 9014 1551 9016
rect 0 8984 800 9014
rect 1485 9011 1551 9014
rect 12566 9012 12572 9076
rect 12636 9074 12642 9076
rect 12709 9074 12775 9077
rect 12636 9072 12775 9074
rect 12636 9016 12714 9072
rect 12770 9016 12775 9072
rect 12636 9014 12775 9016
rect 12636 9012 12642 9014
rect 12709 9011 12775 9014
rect 9622 8876 9628 8940
rect 9692 8938 9698 8940
rect 13169 8938 13235 8941
rect 9692 8936 13235 8938
rect 9692 8880 13174 8936
rect 13230 8880 13235 8936
rect 9692 8878 13235 8880
rect 9692 8876 9698 8878
rect 13169 8875 13235 8878
rect 4694 8736 5010 8737
rect 4694 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5010 8736
rect 4694 8671 5010 8672
rect 8442 8736 8758 8737
rect 8442 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8758 8736
rect 8442 8671 8758 8672
rect 12190 8736 12506 8737
rect 12190 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12506 8736
rect 12190 8671 12506 8672
rect 2820 8192 3136 8193
rect 0 8122 800 8152
rect 2820 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3136 8192
rect 2820 8127 3136 8128
rect 6568 8192 6884 8193
rect 6568 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6884 8192
rect 6568 8127 6884 8128
rect 10316 8192 10632 8193
rect 10316 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10632 8192
rect 10316 8127 10632 8128
rect 14064 8192 14380 8193
rect 14064 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14380 8192
rect 14064 8127 14380 8128
rect 1485 8122 1551 8125
rect 0 8120 1551 8122
rect 0 8064 1490 8120
rect 1546 8064 1551 8120
rect 0 8062 1551 8064
rect 0 8032 800 8062
rect 1485 8059 1551 8062
rect 3601 7850 3667 7853
rect 11697 7850 11763 7853
rect 3601 7848 11763 7850
rect 3601 7792 3606 7848
rect 3662 7792 11702 7848
rect 11758 7792 11763 7848
rect 3601 7790 11763 7792
rect 3601 7787 3667 7790
rect 11697 7787 11763 7790
rect 4694 7648 5010 7649
rect 4694 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5010 7648
rect 4694 7583 5010 7584
rect 8442 7648 8758 7649
rect 8442 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8758 7648
rect 8442 7583 8758 7584
rect 12190 7648 12506 7649
rect 12190 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12506 7648
rect 12190 7583 12506 7584
rect 2313 7306 2379 7309
rect 7281 7306 7347 7309
rect 2313 7304 7347 7306
rect 2313 7248 2318 7304
rect 2374 7248 7286 7304
rect 7342 7248 7347 7304
rect 2313 7246 7347 7248
rect 2313 7243 2379 7246
rect 7281 7243 7347 7246
rect 0 7170 800 7200
rect 1485 7170 1551 7173
rect 0 7168 1551 7170
rect 0 7112 1490 7168
rect 1546 7112 1551 7168
rect 0 7110 1551 7112
rect 0 7080 800 7110
rect 1485 7107 1551 7110
rect 2820 7104 3136 7105
rect 2820 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3136 7104
rect 2820 7039 3136 7040
rect 6568 7104 6884 7105
rect 6568 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6884 7104
rect 6568 7039 6884 7040
rect 10316 7104 10632 7105
rect 10316 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10632 7104
rect 10316 7039 10632 7040
rect 14064 7104 14380 7105
rect 14064 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14380 7104
rect 14064 7039 14380 7040
rect 11421 6762 11487 6765
rect 13118 6762 13124 6764
rect 11421 6760 13124 6762
rect 11421 6704 11426 6760
rect 11482 6704 13124 6760
rect 11421 6702 13124 6704
rect 11421 6699 11487 6702
rect 13118 6700 13124 6702
rect 13188 6700 13194 6764
rect 2129 6626 2195 6629
rect 2262 6626 2268 6628
rect 2129 6624 2268 6626
rect 2129 6568 2134 6624
rect 2190 6568 2268 6624
rect 2129 6566 2268 6568
rect 2129 6563 2195 6566
rect 2262 6564 2268 6566
rect 2332 6626 2338 6628
rect 3550 6626 3556 6628
rect 2332 6566 3556 6626
rect 2332 6564 2338 6566
rect 3550 6564 3556 6566
rect 3620 6564 3626 6628
rect 4694 6560 5010 6561
rect 4694 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5010 6560
rect 4694 6495 5010 6496
rect 8442 6560 8758 6561
rect 8442 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8758 6560
rect 8442 6495 8758 6496
rect 12190 6560 12506 6561
rect 12190 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12506 6560
rect 12190 6495 12506 6496
rect 10961 6354 11027 6357
rect 11646 6354 11652 6356
rect 10961 6352 11652 6354
rect 10961 6296 10966 6352
rect 11022 6296 11652 6352
rect 10961 6294 11652 6296
rect 10961 6291 11027 6294
rect 11646 6292 11652 6294
rect 11716 6354 11722 6356
rect 12341 6354 12407 6357
rect 11716 6352 12407 6354
rect 11716 6296 12346 6352
rect 12402 6296 12407 6352
rect 11716 6294 12407 6296
rect 11716 6292 11722 6294
rect 12341 6291 12407 6294
rect 0 6218 800 6248
rect 1485 6218 1551 6221
rect 0 6216 1551 6218
rect 0 6160 1490 6216
rect 1546 6160 1551 6216
rect 0 6158 1551 6160
rect 0 6128 800 6158
rect 1485 6155 1551 6158
rect 2630 6156 2636 6220
rect 2700 6218 2706 6220
rect 2773 6218 2839 6221
rect 3601 6218 3667 6221
rect 2700 6216 3667 6218
rect 2700 6160 2778 6216
rect 2834 6160 3606 6216
rect 3662 6160 3667 6216
rect 2700 6158 3667 6160
rect 2700 6156 2706 6158
rect 2773 6155 2839 6158
rect 3601 6155 3667 6158
rect 6361 6218 6427 6221
rect 9990 6218 9996 6220
rect 6361 6216 9996 6218
rect 6361 6160 6366 6216
rect 6422 6160 9996 6216
rect 6361 6158 9996 6160
rect 6361 6155 6427 6158
rect 9990 6156 9996 6158
rect 10060 6218 10066 6220
rect 13721 6218 13787 6221
rect 10060 6216 13787 6218
rect 10060 6160 13726 6216
rect 13782 6160 13787 6216
rect 10060 6158 13787 6160
rect 10060 6156 10066 6158
rect 13721 6155 13787 6158
rect 13854 6156 13860 6220
rect 13924 6218 13930 6220
rect 14089 6218 14155 6221
rect 13924 6216 14155 6218
rect 13924 6160 14094 6216
rect 14150 6160 14155 6216
rect 13924 6158 14155 6160
rect 13924 6156 13930 6158
rect 14089 6155 14155 6158
rect 15561 6082 15627 6085
rect 16400 6082 17200 6112
rect 15561 6080 17200 6082
rect 15561 6024 15566 6080
rect 15622 6024 17200 6080
rect 15561 6022 17200 6024
rect 15561 6019 15627 6022
rect 2820 6016 3136 6017
rect 2820 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3136 6016
rect 2820 5951 3136 5952
rect 6568 6016 6884 6017
rect 6568 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6884 6016
rect 6568 5951 6884 5952
rect 10316 6016 10632 6017
rect 10316 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10632 6016
rect 10316 5951 10632 5952
rect 14064 6016 14380 6017
rect 14064 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14380 6016
rect 16400 5992 17200 6022
rect 14064 5951 14380 5952
rect 7557 5946 7623 5949
rect 9121 5946 9187 5949
rect 14917 5946 14983 5949
rect 7557 5944 9187 5946
rect 7557 5888 7562 5944
rect 7618 5888 9126 5944
rect 9182 5888 9187 5944
rect 7557 5886 9187 5888
rect 7557 5883 7623 5886
rect 9121 5883 9187 5886
rect 14460 5944 14983 5946
rect 14460 5888 14922 5944
rect 14978 5888 14983 5944
rect 14460 5886 14983 5888
rect 5073 5810 5139 5813
rect 9213 5810 9279 5813
rect 5073 5808 9279 5810
rect 5073 5752 5078 5808
rect 5134 5752 9218 5808
rect 9274 5752 9279 5808
rect 5073 5750 9279 5752
rect 5073 5747 5139 5750
rect 9213 5747 9279 5750
rect 12566 5748 12572 5812
rect 12636 5810 12642 5812
rect 12709 5810 12775 5813
rect 14460 5810 14520 5886
rect 14917 5883 14983 5886
rect 12636 5808 14520 5810
rect 12636 5752 12714 5808
rect 12770 5752 14520 5808
rect 12636 5750 14520 5752
rect 14641 5810 14707 5813
rect 14774 5810 14780 5812
rect 14641 5808 14780 5810
rect 14641 5752 14646 5808
rect 14702 5752 14780 5808
rect 14641 5750 14780 5752
rect 12636 5748 12642 5750
rect 12709 5747 12775 5750
rect 14641 5747 14707 5750
rect 14774 5748 14780 5750
rect 14844 5748 14850 5812
rect 2497 5674 2563 5677
rect 3969 5674 4035 5677
rect 2497 5672 2790 5674
rect 2497 5616 2502 5672
rect 2558 5616 2790 5672
rect 2497 5614 2790 5616
rect 2497 5611 2563 5614
rect 2730 5538 2790 5614
rect 3969 5672 7482 5674
rect 3969 5616 3974 5672
rect 4030 5616 7482 5672
rect 3969 5614 7482 5616
rect 3969 5611 4035 5614
rect 3325 5538 3391 5541
rect 2730 5536 3391 5538
rect 2730 5480 3330 5536
rect 3386 5480 3391 5536
rect 2730 5478 3391 5480
rect 3325 5475 3391 5478
rect 4694 5472 5010 5473
rect 4694 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5010 5472
rect 4694 5407 5010 5408
rect 7422 5402 7482 5614
rect 9990 5612 9996 5676
rect 10060 5674 10066 5676
rect 15561 5674 15627 5677
rect 10060 5672 15627 5674
rect 10060 5616 15566 5672
rect 15622 5616 15627 5672
rect 10060 5614 15627 5616
rect 10060 5612 10066 5614
rect 15561 5611 15627 5614
rect 10174 5476 10180 5540
rect 10244 5538 10250 5540
rect 10317 5538 10383 5541
rect 10244 5536 10383 5538
rect 10244 5480 10322 5536
rect 10378 5480 10383 5536
rect 10244 5478 10383 5480
rect 10244 5476 10250 5478
rect 10317 5475 10383 5478
rect 14590 5476 14596 5540
rect 14660 5538 14666 5540
rect 15101 5538 15167 5541
rect 14660 5536 15167 5538
rect 14660 5480 15106 5536
rect 15162 5480 15167 5536
rect 14660 5478 15167 5480
rect 14660 5476 14666 5478
rect 15101 5475 15167 5478
rect 8442 5472 8758 5473
rect 8442 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8758 5472
rect 8442 5407 8758 5408
rect 12190 5472 12506 5473
rect 12190 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12506 5472
rect 12190 5407 12506 5408
rect 7741 5402 7807 5405
rect 8017 5402 8083 5405
rect 7422 5400 8083 5402
rect 7422 5344 7746 5400
rect 7802 5344 8022 5400
rect 8078 5344 8083 5400
rect 7422 5342 8083 5344
rect 7741 5339 7807 5342
rect 8017 5339 8083 5342
rect 10133 5402 10199 5405
rect 15009 5404 15075 5405
rect 10910 5402 10916 5404
rect 10133 5400 10916 5402
rect 10133 5344 10138 5400
rect 10194 5344 10916 5400
rect 10133 5342 10916 5344
rect 10133 5339 10199 5342
rect 10910 5340 10916 5342
rect 10980 5340 10986 5404
rect 14958 5340 14964 5404
rect 15028 5402 15075 5404
rect 15028 5400 15120 5402
rect 15070 5344 15120 5400
rect 15028 5342 15120 5344
rect 15028 5340 15075 5342
rect 15009 5339 15075 5340
rect 0 5266 800 5296
rect 1485 5266 1551 5269
rect 0 5264 1551 5266
rect 0 5208 1490 5264
rect 1546 5208 1551 5264
rect 0 5206 1551 5208
rect 0 5176 800 5206
rect 1485 5203 1551 5206
rect 2497 5266 2563 5269
rect 12065 5266 12131 5269
rect 2497 5264 12131 5266
rect 2497 5208 2502 5264
rect 2558 5208 12070 5264
rect 12126 5208 12131 5264
rect 2497 5206 12131 5208
rect 2497 5203 2563 5206
rect 12065 5203 12131 5206
rect 12249 5266 12315 5269
rect 15285 5266 15351 5269
rect 12249 5264 15351 5266
rect 12249 5208 12254 5264
rect 12310 5208 15290 5264
rect 15346 5208 15351 5264
rect 12249 5206 15351 5208
rect 12249 5203 12315 5206
rect 15285 5203 15351 5206
rect 2262 5068 2268 5132
rect 2332 5130 2338 5132
rect 3141 5130 3207 5133
rect 14089 5130 14155 5133
rect 2332 5128 14155 5130
rect 2332 5072 3146 5128
rect 3202 5072 14094 5128
rect 14150 5072 14155 5128
rect 2332 5070 14155 5072
rect 2332 5068 2338 5070
rect 3141 5067 3207 5070
rect 14089 5067 14155 5070
rect 3785 4994 3851 4997
rect 6085 4994 6151 4997
rect 3785 4992 6151 4994
rect 3785 4936 3790 4992
rect 3846 4936 6090 4992
rect 6146 4936 6151 4992
rect 3785 4934 6151 4936
rect 3785 4931 3851 4934
rect 6085 4931 6151 4934
rect 11973 4994 12039 4997
rect 12566 4994 12572 4996
rect 11973 4992 12572 4994
rect 11973 4936 11978 4992
rect 12034 4936 12572 4992
rect 11973 4934 12572 4936
rect 11973 4931 12039 4934
rect 12566 4932 12572 4934
rect 12636 4932 12642 4996
rect 2820 4928 3136 4929
rect 2820 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3136 4928
rect 2820 4863 3136 4864
rect 6568 4928 6884 4929
rect 6568 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6884 4928
rect 6568 4863 6884 4864
rect 10316 4928 10632 4929
rect 10316 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10632 4928
rect 10316 4863 10632 4864
rect 14064 4928 14380 4929
rect 14064 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14380 4928
rect 14064 4863 14380 4864
rect 7373 4858 7439 4861
rect 8109 4858 8175 4861
rect 9857 4860 9923 4861
rect 9806 4858 9812 4860
rect 7373 4856 8175 4858
rect 7373 4800 7378 4856
rect 7434 4800 8114 4856
rect 8170 4800 8175 4856
rect 7373 4798 8175 4800
rect 9766 4798 9812 4858
rect 9876 4856 9923 4860
rect 9918 4800 9923 4856
rect 7373 4795 7439 4798
rect 8109 4795 8175 4798
rect 9806 4796 9812 4798
rect 9876 4796 9923 4800
rect 9857 4795 9923 4796
rect 2630 4660 2636 4724
rect 2700 4722 2706 4724
rect 3049 4722 3115 4725
rect 2700 4720 3115 4722
rect 2700 4664 3054 4720
rect 3110 4664 3115 4720
rect 2700 4662 3115 4664
rect 2700 4660 2706 4662
rect 3049 4659 3115 4662
rect 5625 4722 5691 4725
rect 5625 4720 12450 4722
rect 5625 4664 5630 4720
rect 5686 4664 12450 4720
rect 5625 4662 12450 4664
rect 5625 4659 5691 4662
rect 2773 4586 2839 4589
rect 4797 4586 4863 4589
rect 6821 4586 6887 4589
rect 10501 4586 10567 4589
rect 12065 4586 12131 4589
rect 2773 4584 5458 4586
rect 2773 4528 2778 4584
rect 2834 4528 4802 4584
rect 4858 4528 5458 4584
rect 2773 4526 5458 4528
rect 2773 4523 2839 4526
rect 4797 4523 4863 4526
rect 5398 4453 5458 4526
rect 6821 4584 10242 4586
rect 6821 4528 6826 4584
rect 6882 4528 10242 4584
rect 6821 4526 10242 4528
rect 6821 4523 6887 4526
rect 5398 4448 5507 4453
rect 5398 4392 5446 4448
rect 5502 4392 5507 4448
rect 5398 4390 5507 4392
rect 5441 4387 5507 4390
rect 4694 4384 5010 4385
rect 0 4314 800 4344
rect 4694 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5010 4384
rect 4694 4319 5010 4320
rect 8442 4384 8758 4385
rect 8442 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8758 4384
rect 8442 4319 8758 4320
rect 1485 4314 1551 4317
rect 0 4312 1551 4314
rect 0 4256 1490 4312
rect 1546 4256 1551 4312
rect 0 4254 1551 4256
rect 0 4224 800 4254
rect 1485 4251 1551 4254
rect 5574 4252 5580 4316
rect 5644 4314 5650 4316
rect 7281 4314 7347 4317
rect 5644 4312 7347 4314
rect 5644 4256 7286 4312
rect 7342 4256 7347 4312
rect 5644 4254 7347 4256
rect 5644 4252 5650 4254
rect 7281 4251 7347 4254
rect 10041 4178 10107 4181
rect 2730 4176 10107 4178
rect 2730 4120 10046 4176
rect 10102 4120 10107 4176
rect 2730 4118 10107 4120
rect 10182 4178 10242 4526
rect 10501 4584 12131 4586
rect 10501 4528 10506 4584
rect 10562 4528 12070 4584
rect 12126 4528 12131 4584
rect 10501 4526 12131 4528
rect 12390 4586 12450 4662
rect 12390 4526 14290 4586
rect 10501 4523 10567 4526
rect 12065 4523 12131 4526
rect 11145 4452 11211 4453
rect 11094 4450 11100 4452
rect 11054 4390 11100 4450
rect 11164 4448 11211 4452
rect 11206 4392 11211 4448
rect 11094 4388 11100 4390
rect 11164 4388 11211 4392
rect 14230 4450 14290 4526
rect 14457 4450 14523 4453
rect 14590 4450 14596 4452
rect 14230 4448 14596 4450
rect 14230 4392 14462 4448
rect 14518 4392 14596 4448
rect 14230 4390 14596 4392
rect 11145 4387 11211 4388
rect 14457 4387 14523 4390
rect 14590 4388 14596 4390
rect 14660 4388 14666 4452
rect 12190 4384 12506 4385
rect 12190 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12506 4384
rect 12190 4319 12506 4320
rect 11237 4316 11303 4317
rect 11237 4312 11284 4316
rect 11348 4314 11354 4316
rect 11237 4256 11242 4312
rect 11237 4252 11284 4256
rect 11348 4254 11394 4314
rect 11348 4252 11354 4254
rect 11237 4251 11303 4252
rect 15377 4178 15443 4181
rect 10182 4176 15443 4178
rect 10182 4120 15382 4176
rect 15438 4120 15443 4176
rect 10182 4118 15443 4120
rect 1577 4042 1643 4045
rect 2730 4042 2790 4118
rect 10041 4115 10107 4118
rect 15377 4115 15443 4118
rect 1577 4040 2790 4042
rect 1577 3984 1582 4040
rect 1638 3984 2790 4040
rect 1577 3982 2790 3984
rect 5441 4042 5507 4045
rect 9857 4042 9923 4045
rect 9990 4042 9996 4044
rect 5441 4040 7114 4042
rect 5441 3984 5446 4040
rect 5502 3984 7114 4040
rect 5441 3982 7114 3984
rect 1577 3979 1643 3982
rect 5441 3979 5507 3982
rect 7054 3906 7114 3982
rect 9857 4040 9996 4042
rect 9857 3984 9862 4040
rect 9918 3984 9996 4040
rect 9857 3982 9996 3984
rect 9857 3979 9923 3982
rect 9990 3980 9996 3982
rect 10060 3980 10066 4044
rect 10182 3982 10794 4042
rect 10182 3906 10242 3982
rect 7054 3846 10242 3906
rect 10734 3906 10794 3982
rect 12014 3980 12020 4044
rect 12084 4042 12090 4044
rect 12341 4042 12407 4045
rect 14825 4044 14891 4045
rect 12084 4040 12407 4042
rect 12084 3984 12346 4040
rect 12402 3984 12407 4040
rect 12084 3982 12407 3984
rect 12084 3980 12090 3982
rect 12022 3906 12082 3980
rect 12341 3979 12407 3982
rect 14774 3980 14780 4044
rect 14844 4042 14891 4044
rect 14844 4040 14936 4042
rect 14886 3984 14936 4040
rect 14844 3982 14936 3984
rect 14844 3980 14891 3982
rect 14825 3979 14891 3980
rect 13721 3906 13787 3909
rect 10734 3846 12082 3906
rect 12390 3904 13787 3906
rect 12390 3848 13726 3904
rect 13782 3848 13787 3904
rect 12390 3846 13787 3848
rect 2820 3840 3136 3841
rect 2820 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3136 3840
rect 2820 3775 3136 3776
rect 6568 3840 6884 3841
rect 6568 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6884 3840
rect 6568 3775 6884 3776
rect 10316 3840 10632 3841
rect 10316 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10632 3840
rect 10316 3775 10632 3776
rect 9397 3770 9463 3773
rect 7100 3768 9463 3770
rect 7100 3712 9402 3768
rect 9458 3712 9463 3768
rect 7100 3710 9463 3712
rect 7100 3637 7160 3710
rect 9397 3707 9463 3710
rect 11094 3708 11100 3772
rect 11164 3770 11170 3772
rect 11237 3770 11303 3773
rect 11164 3768 11303 3770
rect 11164 3712 11242 3768
rect 11298 3712 11303 3768
rect 11164 3710 11303 3712
rect 11164 3708 11170 3710
rect 11237 3707 11303 3710
rect 1853 3634 1919 3637
rect 4153 3634 4219 3637
rect 1853 3632 4219 3634
rect 1853 3576 1858 3632
rect 1914 3576 4158 3632
rect 4214 3576 4219 3632
rect 1853 3574 4219 3576
rect 1853 3571 1919 3574
rect 4153 3571 4219 3574
rect 4429 3634 4495 3637
rect 5533 3634 5599 3637
rect 7097 3634 7163 3637
rect 4429 3632 7163 3634
rect 4429 3576 4434 3632
rect 4490 3576 5538 3632
rect 5594 3576 7102 3632
rect 7158 3576 7163 3632
rect 4429 3574 7163 3576
rect 4429 3571 4495 3574
rect 5533 3571 5599 3574
rect 7097 3571 7163 3574
rect 7230 3572 7236 3636
rect 7300 3634 7306 3636
rect 12390 3634 12450 3846
rect 13721 3843 13787 3846
rect 14064 3840 14380 3841
rect 14064 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14380 3840
rect 14064 3775 14380 3776
rect 7300 3574 12450 3634
rect 7300 3572 7306 3574
rect 4061 3498 4127 3501
rect 10225 3498 10291 3501
rect 14365 3498 14431 3501
rect 4061 3496 9322 3498
rect 4061 3440 4066 3496
rect 4122 3440 9322 3496
rect 4061 3438 9322 3440
rect 4061 3435 4127 3438
rect 0 3362 800 3392
rect 1577 3362 1643 3365
rect 5533 3364 5599 3365
rect 5533 3362 5580 3364
rect 0 3360 1643 3362
rect 0 3304 1582 3360
rect 1638 3304 1643 3360
rect 0 3302 1643 3304
rect 5488 3360 5580 3362
rect 5488 3304 5538 3360
rect 5488 3302 5580 3304
rect 0 3272 800 3302
rect 1577 3299 1643 3302
rect 5533 3300 5580 3302
rect 5644 3300 5650 3364
rect 6085 3362 6151 3365
rect 7925 3362 7991 3365
rect 6085 3360 7991 3362
rect 6085 3304 6090 3360
rect 6146 3304 7930 3360
rect 7986 3304 7991 3360
rect 6085 3302 7991 3304
rect 5533 3299 5599 3300
rect 6085 3299 6151 3302
rect 7925 3299 7991 3302
rect 4694 3296 5010 3297
rect 4694 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5010 3296
rect 4694 3231 5010 3232
rect 8442 3296 8758 3297
rect 8442 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8758 3296
rect 8442 3231 8758 3232
rect 9262 3090 9322 3438
rect 10225 3496 14431 3498
rect 10225 3440 10230 3496
rect 10286 3440 14370 3496
rect 14426 3440 14431 3496
rect 10225 3438 14431 3440
rect 10225 3435 10291 3438
rect 14365 3435 14431 3438
rect 12190 3296 12506 3297
rect 12190 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12506 3296
rect 12190 3231 12506 3232
rect 9806 3164 9812 3228
rect 9876 3226 9882 3228
rect 9949 3226 10015 3229
rect 9876 3224 10015 3226
rect 9876 3168 9954 3224
rect 10010 3168 10015 3224
rect 9876 3166 10015 3168
rect 9876 3164 9882 3166
rect 9949 3163 10015 3166
rect 10910 3164 10916 3228
rect 10980 3226 10986 3228
rect 11329 3226 11395 3229
rect 10980 3224 11395 3226
rect 10980 3168 11334 3224
rect 11390 3168 11395 3224
rect 10980 3166 11395 3168
rect 10980 3164 10986 3166
rect 11329 3163 11395 3166
rect 10317 3090 10383 3093
rect 11646 3090 11652 3092
rect 9262 3088 11652 3090
rect 9262 3032 10322 3088
rect 10378 3032 11652 3088
rect 9262 3030 11652 3032
rect 10317 3027 10383 3030
rect 11646 3028 11652 3030
rect 11716 3090 11722 3092
rect 11973 3090 12039 3093
rect 14089 3090 14155 3093
rect 11716 3088 12039 3090
rect 11716 3032 11978 3088
rect 12034 3032 12039 3088
rect 11716 3030 12039 3032
rect 11716 3028 11722 3030
rect 11973 3027 12039 3030
rect 12390 3088 14155 3090
rect 12390 3032 14094 3088
rect 14150 3032 14155 3088
rect 12390 3030 14155 3032
rect 3233 2954 3299 2957
rect 7230 2954 7236 2956
rect 3233 2952 7236 2954
rect 3233 2896 3238 2952
rect 3294 2896 7236 2952
rect 3233 2894 7236 2896
rect 3233 2891 3299 2894
rect 7230 2892 7236 2894
rect 7300 2892 7306 2956
rect 7741 2954 7807 2957
rect 12390 2954 12450 3030
rect 14089 3027 14155 3030
rect 7741 2952 12450 2954
rect 7741 2896 7746 2952
rect 7802 2896 12450 2952
rect 7741 2894 12450 2896
rect 13813 2956 13879 2957
rect 13813 2952 13860 2956
rect 13924 2954 13930 2956
rect 13813 2896 13818 2952
rect 7741 2891 7807 2894
rect 13813 2892 13860 2896
rect 13924 2894 13970 2954
rect 13924 2892 13930 2894
rect 13813 2891 13879 2892
rect 7189 2818 7255 2821
rect 9857 2818 9923 2821
rect 10174 2818 10180 2820
rect 7189 2816 10180 2818
rect 7189 2760 7194 2816
rect 7250 2760 9862 2816
rect 9918 2760 10180 2816
rect 7189 2758 10180 2760
rect 7189 2755 7255 2758
rect 9857 2755 9923 2758
rect 10174 2756 10180 2758
rect 10244 2756 10250 2820
rect 2820 2752 3136 2753
rect 2820 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3136 2752
rect 2820 2687 3136 2688
rect 6568 2752 6884 2753
rect 6568 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6884 2752
rect 6568 2687 6884 2688
rect 10316 2752 10632 2753
rect 10316 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10632 2752
rect 10316 2687 10632 2688
rect 14064 2752 14380 2753
rect 14064 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14380 2752
rect 14064 2687 14380 2688
rect 13670 2484 13676 2548
rect 13740 2546 13746 2548
rect 14365 2546 14431 2549
rect 13740 2544 14431 2546
rect 13740 2488 14370 2544
rect 14426 2488 14431 2544
rect 13740 2486 14431 2488
rect 13740 2484 13746 2486
rect 14365 2483 14431 2486
rect 0 2410 800 2440
rect 3601 2410 3667 2413
rect 3918 2410 3924 2412
rect 0 2408 3924 2410
rect 0 2352 3606 2408
rect 3662 2352 3924 2408
rect 0 2350 3924 2352
rect 0 2320 800 2350
rect 3601 2347 3667 2350
rect 3918 2348 3924 2350
rect 3988 2348 3994 2412
rect 4694 2208 5010 2209
rect 4694 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5010 2208
rect 4694 2143 5010 2144
rect 8442 2208 8758 2209
rect 8442 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8758 2208
rect 8442 2143 8758 2144
rect 12190 2208 12506 2209
rect 12190 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12506 2208
rect 12190 2143 12506 2144
rect 14641 2138 14707 2141
rect 16400 2138 17200 2168
rect 14641 2136 17200 2138
rect 14641 2080 14646 2136
rect 14702 2080 17200 2136
rect 14641 2078 17200 2080
rect 14641 2075 14707 2078
rect 16400 2048 17200 2078
rect 0 1458 800 1488
rect 2497 1458 2563 1461
rect 0 1456 2563 1458
rect 0 1400 2502 1456
rect 2558 1400 2563 1456
rect 0 1398 2563 1400
rect 0 1368 800 1398
rect 2497 1395 2563 1398
rect 0 506 800 536
rect 1894 506 1900 508
rect 0 446 1900 506
rect 0 416 800 446
rect 1894 444 1900 446
rect 1964 444 1970 508
<< via3 >>
rect 4700 17436 4764 17440
rect 4700 17380 4704 17436
rect 4704 17380 4760 17436
rect 4760 17380 4764 17436
rect 4700 17376 4764 17380
rect 4780 17436 4844 17440
rect 4780 17380 4784 17436
rect 4784 17380 4840 17436
rect 4840 17380 4844 17436
rect 4780 17376 4844 17380
rect 4860 17436 4924 17440
rect 4860 17380 4864 17436
rect 4864 17380 4920 17436
rect 4920 17380 4924 17436
rect 4860 17376 4924 17380
rect 4940 17436 5004 17440
rect 4940 17380 4944 17436
rect 4944 17380 5000 17436
rect 5000 17380 5004 17436
rect 4940 17376 5004 17380
rect 8448 17436 8512 17440
rect 8448 17380 8452 17436
rect 8452 17380 8508 17436
rect 8508 17380 8512 17436
rect 8448 17376 8512 17380
rect 8528 17436 8592 17440
rect 8528 17380 8532 17436
rect 8532 17380 8588 17436
rect 8588 17380 8592 17436
rect 8528 17376 8592 17380
rect 8608 17436 8672 17440
rect 8608 17380 8612 17436
rect 8612 17380 8668 17436
rect 8668 17380 8672 17436
rect 8608 17376 8672 17380
rect 8688 17436 8752 17440
rect 8688 17380 8692 17436
rect 8692 17380 8748 17436
rect 8748 17380 8752 17436
rect 8688 17376 8752 17380
rect 12196 17436 12260 17440
rect 12196 17380 12200 17436
rect 12200 17380 12256 17436
rect 12256 17380 12260 17436
rect 12196 17376 12260 17380
rect 12276 17436 12340 17440
rect 12276 17380 12280 17436
rect 12280 17380 12336 17436
rect 12336 17380 12340 17436
rect 12276 17376 12340 17380
rect 12356 17436 12420 17440
rect 12356 17380 12360 17436
rect 12360 17380 12416 17436
rect 12416 17380 12420 17436
rect 12356 17376 12420 17380
rect 12436 17436 12500 17440
rect 12436 17380 12440 17436
rect 12440 17380 12496 17436
rect 12496 17380 12500 17436
rect 12436 17376 12500 17380
rect 10732 17172 10796 17236
rect 2826 16892 2890 16896
rect 2826 16836 2830 16892
rect 2830 16836 2886 16892
rect 2886 16836 2890 16892
rect 2826 16832 2890 16836
rect 2906 16892 2970 16896
rect 2906 16836 2910 16892
rect 2910 16836 2966 16892
rect 2966 16836 2970 16892
rect 2906 16832 2970 16836
rect 2986 16892 3050 16896
rect 2986 16836 2990 16892
rect 2990 16836 3046 16892
rect 3046 16836 3050 16892
rect 2986 16832 3050 16836
rect 3066 16892 3130 16896
rect 3066 16836 3070 16892
rect 3070 16836 3126 16892
rect 3126 16836 3130 16892
rect 3066 16832 3130 16836
rect 6574 16892 6638 16896
rect 6574 16836 6578 16892
rect 6578 16836 6634 16892
rect 6634 16836 6638 16892
rect 6574 16832 6638 16836
rect 6654 16892 6718 16896
rect 6654 16836 6658 16892
rect 6658 16836 6714 16892
rect 6714 16836 6718 16892
rect 6654 16832 6718 16836
rect 6734 16892 6798 16896
rect 6734 16836 6738 16892
rect 6738 16836 6794 16892
rect 6794 16836 6798 16892
rect 6734 16832 6798 16836
rect 6814 16892 6878 16896
rect 6814 16836 6818 16892
rect 6818 16836 6874 16892
rect 6874 16836 6878 16892
rect 6814 16832 6878 16836
rect 10322 16892 10386 16896
rect 10322 16836 10326 16892
rect 10326 16836 10382 16892
rect 10382 16836 10386 16892
rect 10322 16832 10386 16836
rect 10402 16892 10466 16896
rect 10402 16836 10406 16892
rect 10406 16836 10462 16892
rect 10462 16836 10466 16892
rect 10402 16832 10466 16836
rect 10482 16892 10546 16896
rect 10482 16836 10486 16892
rect 10486 16836 10542 16892
rect 10542 16836 10546 16892
rect 10482 16832 10546 16836
rect 10562 16892 10626 16896
rect 10562 16836 10566 16892
rect 10566 16836 10622 16892
rect 10622 16836 10626 16892
rect 10562 16832 10626 16836
rect 9444 16764 9508 16828
rect 13860 17036 13924 17100
rect 10916 16900 10980 16964
rect 14070 16892 14134 16896
rect 14070 16836 14074 16892
rect 14074 16836 14130 16892
rect 14130 16836 14134 16892
rect 14070 16832 14134 16836
rect 14150 16892 14214 16896
rect 14150 16836 14154 16892
rect 14154 16836 14210 16892
rect 14210 16836 14214 16892
rect 14150 16832 14214 16836
rect 14230 16892 14294 16896
rect 14230 16836 14234 16892
rect 14234 16836 14290 16892
rect 14290 16836 14294 16892
rect 14230 16832 14294 16836
rect 14310 16892 14374 16896
rect 14310 16836 14314 16892
rect 14314 16836 14370 16892
rect 14370 16836 14374 16892
rect 14310 16832 14374 16836
rect 11836 16688 11900 16692
rect 11836 16632 11850 16688
rect 11850 16632 11900 16688
rect 11836 16628 11900 16632
rect 12572 16628 12636 16692
rect 13492 16688 13556 16692
rect 13492 16632 13506 16688
rect 13506 16632 13556 16688
rect 13492 16628 13556 16632
rect 14780 16628 14844 16692
rect 9628 16492 9692 16556
rect 4700 16348 4764 16352
rect 4700 16292 4704 16348
rect 4704 16292 4760 16348
rect 4760 16292 4764 16348
rect 4700 16288 4764 16292
rect 4780 16348 4844 16352
rect 4780 16292 4784 16348
rect 4784 16292 4840 16348
rect 4840 16292 4844 16348
rect 4780 16288 4844 16292
rect 4860 16348 4924 16352
rect 4860 16292 4864 16348
rect 4864 16292 4920 16348
rect 4920 16292 4924 16348
rect 4860 16288 4924 16292
rect 4940 16348 5004 16352
rect 4940 16292 4944 16348
rect 4944 16292 5000 16348
rect 5000 16292 5004 16348
rect 4940 16288 5004 16292
rect 8448 16348 8512 16352
rect 8448 16292 8452 16348
rect 8452 16292 8508 16348
rect 8508 16292 8512 16348
rect 8448 16288 8512 16292
rect 8528 16348 8592 16352
rect 8528 16292 8532 16348
rect 8532 16292 8588 16348
rect 8588 16292 8592 16348
rect 8528 16288 8592 16292
rect 8608 16348 8672 16352
rect 8608 16292 8612 16348
rect 8612 16292 8668 16348
rect 8668 16292 8672 16348
rect 8608 16288 8672 16292
rect 8688 16348 8752 16352
rect 8688 16292 8692 16348
rect 8692 16292 8748 16348
rect 8748 16292 8752 16348
rect 8688 16288 8752 16292
rect 12196 16348 12260 16352
rect 12196 16292 12200 16348
rect 12200 16292 12256 16348
rect 12256 16292 12260 16348
rect 12196 16288 12260 16292
rect 12276 16348 12340 16352
rect 12276 16292 12280 16348
rect 12280 16292 12336 16348
rect 12336 16292 12340 16348
rect 12276 16288 12340 16292
rect 12356 16348 12420 16352
rect 12356 16292 12360 16348
rect 12360 16292 12416 16348
rect 12416 16292 12420 16348
rect 12356 16288 12420 16292
rect 12436 16348 12500 16352
rect 12436 16292 12440 16348
rect 12440 16292 12496 16348
rect 12496 16292 12500 16348
rect 12436 16288 12500 16292
rect 8892 15948 8956 16012
rect 10180 15948 10244 16012
rect 7788 15812 7852 15876
rect 2826 15804 2890 15808
rect 2826 15748 2830 15804
rect 2830 15748 2886 15804
rect 2886 15748 2890 15804
rect 2826 15744 2890 15748
rect 2906 15804 2970 15808
rect 2906 15748 2910 15804
rect 2910 15748 2966 15804
rect 2966 15748 2970 15804
rect 2906 15744 2970 15748
rect 2986 15804 3050 15808
rect 2986 15748 2990 15804
rect 2990 15748 3046 15804
rect 3046 15748 3050 15804
rect 2986 15744 3050 15748
rect 3066 15804 3130 15808
rect 3066 15748 3070 15804
rect 3070 15748 3126 15804
rect 3126 15748 3130 15804
rect 3066 15744 3130 15748
rect 6574 15804 6638 15808
rect 6574 15748 6578 15804
rect 6578 15748 6634 15804
rect 6634 15748 6638 15804
rect 6574 15744 6638 15748
rect 6654 15804 6718 15808
rect 6654 15748 6658 15804
rect 6658 15748 6714 15804
rect 6714 15748 6718 15804
rect 6654 15744 6718 15748
rect 6734 15804 6798 15808
rect 6734 15748 6738 15804
rect 6738 15748 6794 15804
rect 6794 15748 6798 15804
rect 6734 15744 6798 15748
rect 6814 15804 6878 15808
rect 6814 15748 6818 15804
rect 6818 15748 6874 15804
rect 6874 15748 6878 15804
rect 6814 15744 6878 15748
rect 10322 15804 10386 15808
rect 10322 15748 10326 15804
rect 10326 15748 10382 15804
rect 10382 15748 10386 15804
rect 10322 15744 10386 15748
rect 10402 15804 10466 15808
rect 10402 15748 10406 15804
rect 10406 15748 10462 15804
rect 10462 15748 10466 15804
rect 10402 15744 10466 15748
rect 10482 15804 10546 15808
rect 10482 15748 10486 15804
rect 10486 15748 10542 15804
rect 10542 15748 10546 15804
rect 10482 15744 10546 15748
rect 10562 15804 10626 15808
rect 10562 15748 10566 15804
rect 10566 15748 10622 15804
rect 10622 15748 10626 15804
rect 10562 15744 10626 15748
rect 14070 15804 14134 15808
rect 14070 15748 14074 15804
rect 14074 15748 14130 15804
rect 14130 15748 14134 15804
rect 14070 15744 14134 15748
rect 14150 15804 14214 15808
rect 14150 15748 14154 15804
rect 14154 15748 14210 15804
rect 14210 15748 14214 15804
rect 14150 15744 14214 15748
rect 14230 15804 14294 15808
rect 14230 15748 14234 15804
rect 14234 15748 14290 15804
rect 14290 15748 14294 15804
rect 14230 15744 14294 15748
rect 14310 15804 14374 15808
rect 14310 15748 14314 15804
rect 14314 15748 14370 15804
rect 14370 15748 14374 15804
rect 14310 15744 14374 15748
rect 9444 15676 9508 15740
rect 1900 15268 1964 15332
rect 14596 15328 14660 15332
rect 14596 15272 14610 15328
rect 14610 15272 14660 15328
rect 14596 15268 14660 15272
rect 4700 15260 4764 15264
rect 4700 15204 4704 15260
rect 4704 15204 4760 15260
rect 4760 15204 4764 15260
rect 4700 15200 4764 15204
rect 4780 15260 4844 15264
rect 4780 15204 4784 15260
rect 4784 15204 4840 15260
rect 4840 15204 4844 15260
rect 4780 15200 4844 15204
rect 4860 15260 4924 15264
rect 4860 15204 4864 15260
rect 4864 15204 4920 15260
rect 4920 15204 4924 15260
rect 4860 15200 4924 15204
rect 4940 15260 5004 15264
rect 4940 15204 4944 15260
rect 4944 15204 5000 15260
rect 5000 15204 5004 15260
rect 4940 15200 5004 15204
rect 8448 15260 8512 15264
rect 8448 15204 8452 15260
rect 8452 15204 8508 15260
rect 8508 15204 8512 15260
rect 8448 15200 8512 15204
rect 8528 15260 8592 15264
rect 8528 15204 8532 15260
rect 8532 15204 8588 15260
rect 8588 15204 8592 15260
rect 8528 15200 8592 15204
rect 8608 15260 8672 15264
rect 8608 15204 8612 15260
rect 8612 15204 8668 15260
rect 8668 15204 8672 15260
rect 8608 15200 8672 15204
rect 8688 15260 8752 15264
rect 8688 15204 8692 15260
rect 8692 15204 8748 15260
rect 8748 15204 8752 15260
rect 8688 15200 8752 15204
rect 12196 15260 12260 15264
rect 12196 15204 12200 15260
rect 12200 15204 12256 15260
rect 12256 15204 12260 15260
rect 12196 15200 12260 15204
rect 12276 15260 12340 15264
rect 12276 15204 12280 15260
rect 12280 15204 12336 15260
rect 12336 15204 12340 15260
rect 12276 15200 12340 15204
rect 12356 15260 12420 15264
rect 12356 15204 12360 15260
rect 12360 15204 12416 15260
rect 12416 15204 12420 15260
rect 12356 15200 12420 15204
rect 12436 15260 12500 15264
rect 12436 15204 12440 15260
rect 12440 15204 12496 15260
rect 12496 15204 12500 15260
rect 12436 15200 12500 15204
rect 12940 14996 13004 15060
rect 7788 14724 7852 14788
rect 13676 14724 13740 14788
rect 2826 14716 2890 14720
rect 2826 14660 2830 14716
rect 2830 14660 2886 14716
rect 2886 14660 2890 14716
rect 2826 14656 2890 14660
rect 2906 14716 2970 14720
rect 2906 14660 2910 14716
rect 2910 14660 2966 14716
rect 2966 14660 2970 14716
rect 2906 14656 2970 14660
rect 2986 14716 3050 14720
rect 2986 14660 2990 14716
rect 2990 14660 3046 14716
rect 3046 14660 3050 14716
rect 2986 14656 3050 14660
rect 3066 14716 3130 14720
rect 3066 14660 3070 14716
rect 3070 14660 3126 14716
rect 3126 14660 3130 14716
rect 3066 14656 3130 14660
rect 6574 14716 6638 14720
rect 6574 14660 6578 14716
rect 6578 14660 6634 14716
rect 6634 14660 6638 14716
rect 6574 14656 6638 14660
rect 6654 14716 6718 14720
rect 6654 14660 6658 14716
rect 6658 14660 6714 14716
rect 6714 14660 6718 14716
rect 6654 14656 6718 14660
rect 6734 14716 6798 14720
rect 6734 14660 6738 14716
rect 6738 14660 6794 14716
rect 6794 14660 6798 14716
rect 6734 14656 6798 14660
rect 6814 14716 6878 14720
rect 6814 14660 6818 14716
rect 6818 14660 6874 14716
rect 6874 14660 6878 14716
rect 6814 14656 6878 14660
rect 10322 14716 10386 14720
rect 10322 14660 10326 14716
rect 10326 14660 10382 14716
rect 10382 14660 10386 14716
rect 10322 14656 10386 14660
rect 10402 14716 10466 14720
rect 10402 14660 10406 14716
rect 10406 14660 10462 14716
rect 10462 14660 10466 14716
rect 10402 14656 10466 14660
rect 10482 14716 10546 14720
rect 10482 14660 10486 14716
rect 10486 14660 10542 14716
rect 10542 14660 10546 14716
rect 10482 14656 10546 14660
rect 10562 14716 10626 14720
rect 10562 14660 10566 14716
rect 10566 14660 10622 14716
rect 10622 14660 10626 14716
rect 10562 14656 10626 14660
rect 14070 14716 14134 14720
rect 14070 14660 14074 14716
rect 14074 14660 14130 14716
rect 14130 14660 14134 14716
rect 14070 14656 14134 14660
rect 14150 14716 14214 14720
rect 14150 14660 14154 14716
rect 14154 14660 14210 14716
rect 14210 14660 14214 14716
rect 14150 14656 14214 14660
rect 14230 14716 14294 14720
rect 14230 14660 14234 14716
rect 14234 14660 14290 14716
rect 14290 14660 14294 14716
rect 14230 14656 14294 14660
rect 14310 14716 14374 14720
rect 14310 14660 14314 14716
rect 14314 14660 14370 14716
rect 14370 14660 14374 14716
rect 14310 14656 14374 14660
rect 8892 14452 8956 14516
rect 1900 14316 1964 14380
rect 9996 14240 10060 14244
rect 9996 14184 10010 14240
rect 10010 14184 10060 14240
rect 9996 14180 10060 14184
rect 15148 14180 15212 14244
rect 4700 14172 4764 14176
rect 4700 14116 4704 14172
rect 4704 14116 4760 14172
rect 4760 14116 4764 14172
rect 4700 14112 4764 14116
rect 4780 14172 4844 14176
rect 4780 14116 4784 14172
rect 4784 14116 4840 14172
rect 4840 14116 4844 14172
rect 4780 14112 4844 14116
rect 4860 14172 4924 14176
rect 4860 14116 4864 14172
rect 4864 14116 4920 14172
rect 4920 14116 4924 14172
rect 4860 14112 4924 14116
rect 4940 14172 5004 14176
rect 4940 14116 4944 14172
rect 4944 14116 5000 14172
rect 5000 14116 5004 14172
rect 4940 14112 5004 14116
rect 8448 14172 8512 14176
rect 8448 14116 8452 14172
rect 8452 14116 8508 14172
rect 8508 14116 8512 14172
rect 8448 14112 8512 14116
rect 8528 14172 8592 14176
rect 8528 14116 8532 14172
rect 8532 14116 8588 14172
rect 8588 14116 8592 14172
rect 8528 14112 8592 14116
rect 8608 14172 8672 14176
rect 8608 14116 8612 14172
rect 8612 14116 8668 14172
rect 8668 14116 8672 14172
rect 8608 14112 8672 14116
rect 8688 14172 8752 14176
rect 8688 14116 8692 14172
rect 8692 14116 8748 14172
rect 8748 14116 8752 14172
rect 8688 14112 8752 14116
rect 12196 14172 12260 14176
rect 12196 14116 12200 14172
rect 12200 14116 12256 14172
rect 12256 14116 12260 14172
rect 12196 14112 12260 14116
rect 12276 14172 12340 14176
rect 12276 14116 12280 14172
rect 12280 14116 12336 14172
rect 12336 14116 12340 14172
rect 12276 14112 12340 14116
rect 12356 14172 12420 14176
rect 12356 14116 12360 14172
rect 12360 14116 12416 14172
rect 12416 14116 12420 14172
rect 12356 14112 12420 14116
rect 12436 14172 12500 14176
rect 12436 14116 12440 14172
rect 12440 14116 12496 14172
rect 12496 14116 12500 14172
rect 12436 14112 12500 14116
rect 10916 14104 10980 14108
rect 10916 14048 10966 14104
rect 10966 14048 10980 14104
rect 10916 14044 10980 14048
rect 3372 13772 3436 13836
rect 2826 13628 2890 13632
rect 2826 13572 2830 13628
rect 2830 13572 2886 13628
rect 2886 13572 2890 13628
rect 2826 13568 2890 13572
rect 2906 13628 2970 13632
rect 2906 13572 2910 13628
rect 2910 13572 2966 13628
rect 2966 13572 2970 13628
rect 2906 13568 2970 13572
rect 2986 13628 3050 13632
rect 2986 13572 2990 13628
rect 2990 13572 3046 13628
rect 3046 13572 3050 13628
rect 2986 13568 3050 13572
rect 3066 13628 3130 13632
rect 3066 13572 3070 13628
rect 3070 13572 3126 13628
rect 3126 13572 3130 13628
rect 3066 13568 3130 13572
rect 6574 13628 6638 13632
rect 6574 13572 6578 13628
rect 6578 13572 6634 13628
rect 6634 13572 6638 13628
rect 6574 13568 6638 13572
rect 6654 13628 6718 13632
rect 6654 13572 6658 13628
rect 6658 13572 6714 13628
rect 6714 13572 6718 13628
rect 6654 13568 6718 13572
rect 6734 13628 6798 13632
rect 6734 13572 6738 13628
rect 6738 13572 6794 13628
rect 6794 13572 6798 13628
rect 6734 13568 6798 13572
rect 6814 13628 6878 13632
rect 6814 13572 6818 13628
rect 6818 13572 6874 13628
rect 6874 13572 6878 13628
rect 6814 13568 6878 13572
rect 10322 13628 10386 13632
rect 10322 13572 10326 13628
rect 10326 13572 10382 13628
rect 10382 13572 10386 13628
rect 10322 13568 10386 13572
rect 10402 13628 10466 13632
rect 10402 13572 10406 13628
rect 10406 13572 10462 13628
rect 10462 13572 10466 13628
rect 10402 13568 10466 13572
rect 10482 13628 10546 13632
rect 10482 13572 10486 13628
rect 10486 13572 10542 13628
rect 10542 13572 10546 13628
rect 10482 13568 10546 13572
rect 10562 13628 10626 13632
rect 10562 13572 10566 13628
rect 10566 13572 10622 13628
rect 10622 13572 10626 13628
rect 10562 13568 10626 13572
rect 14070 13628 14134 13632
rect 14070 13572 14074 13628
rect 14074 13572 14130 13628
rect 14130 13572 14134 13628
rect 14070 13568 14134 13572
rect 14150 13628 14214 13632
rect 14150 13572 14154 13628
rect 14154 13572 14210 13628
rect 14210 13572 14214 13628
rect 14150 13568 14214 13572
rect 14230 13628 14294 13632
rect 14230 13572 14234 13628
rect 14234 13572 14290 13628
rect 14290 13572 14294 13628
rect 14230 13568 14294 13572
rect 14310 13628 14374 13632
rect 14310 13572 14314 13628
rect 14314 13572 14370 13628
rect 14370 13572 14374 13628
rect 14310 13568 14374 13572
rect 14964 13092 15028 13156
rect 4700 13084 4764 13088
rect 4700 13028 4704 13084
rect 4704 13028 4760 13084
rect 4760 13028 4764 13084
rect 4700 13024 4764 13028
rect 4780 13084 4844 13088
rect 4780 13028 4784 13084
rect 4784 13028 4840 13084
rect 4840 13028 4844 13084
rect 4780 13024 4844 13028
rect 4860 13084 4924 13088
rect 4860 13028 4864 13084
rect 4864 13028 4920 13084
rect 4920 13028 4924 13084
rect 4860 13024 4924 13028
rect 4940 13084 5004 13088
rect 4940 13028 4944 13084
rect 4944 13028 5000 13084
rect 5000 13028 5004 13084
rect 4940 13024 5004 13028
rect 8448 13084 8512 13088
rect 8448 13028 8452 13084
rect 8452 13028 8508 13084
rect 8508 13028 8512 13084
rect 8448 13024 8512 13028
rect 8528 13084 8592 13088
rect 8528 13028 8532 13084
rect 8532 13028 8588 13084
rect 8588 13028 8592 13084
rect 8528 13024 8592 13028
rect 8608 13084 8672 13088
rect 8608 13028 8612 13084
rect 8612 13028 8668 13084
rect 8668 13028 8672 13084
rect 8608 13024 8672 13028
rect 8688 13084 8752 13088
rect 8688 13028 8692 13084
rect 8692 13028 8748 13084
rect 8748 13028 8752 13084
rect 8688 13024 8752 13028
rect 12196 13084 12260 13088
rect 12196 13028 12200 13084
rect 12200 13028 12256 13084
rect 12256 13028 12260 13084
rect 12196 13024 12260 13028
rect 12276 13084 12340 13088
rect 12276 13028 12280 13084
rect 12280 13028 12336 13084
rect 12336 13028 12340 13084
rect 12276 13024 12340 13028
rect 12356 13084 12420 13088
rect 12356 13028 12360 13084
rect 12360 13028 12416 13084
rect 12416 13028 12420 13084
rect 12356 13024 12420 13028
rect 12436 13084 12500 13088
rect 12436 13028 12440 13084
rect 12440 13028 12496 13084
rect 12496 13028 12500 13084
rect 12436 13024 12500 13028
rect 10732 12956 10796 13020
rect 14780 13016 14844 13020
rect 14780 12960 14794 13016
rect 14794 12960 14844 13016
rect 14780 12956 14844 12960
rect 13124 12820 13188 12884
rect 9444 12684 9508 12748
rect 12020 12684 12084 12748
rect 10732 12608 10796 12612
rect 10732 12552 10782 12608
rect 10782 12552 10796 12608
rect 10732 12548 10796 12552
rect 2826 12540 2890 12544
rect 2826 12484 2830 12540
rect 2830 12484 2886 12540
rect 2886 12484 2890 12540
rect 2826 12480 2890 12484
rect 2906 12540 2970 12544
rect 2906 12484 2910 12540
rect 2910 12484 2966 12540
rect 2966 12484 2970 12540
rect 2906 12480 2970 12484
rect 2986 12540 3050 12544
rect 2986 12484 2990 12540
rect 2990 12484 3046 12540
rect 3046 12484 3050 12540
rect 2986 12480 3050 12484
rect 3066 12540 3130 12544
rect 3066 12484 3070 12540
rect 3070 12484 3126 12540
rect 3126 12484 3130 12540
rect 3066 12480 3130 12484
rect 6574 12540 6638 12544
rect 6574 12484 6578 12540
rect 6578 12484 6634 12540
rect 6634 12484 6638 12540
rect 6574 12480 6638 12484
rect 6654 12540 6718 12544
rect 6654 12484 6658 12540
rect 6658 12484 6714 12540
rect 6714 12484 6718 12540
rect 6654 12480 6718 12484
rect 6734 12540 6798 12544
rect 6734 12484 6738 12540
rect 6738 12484 6794 12540
rect 6794 12484 6798 12540
rect 6734 12480 6798 12484
rect 6814 12540 6878 12544
rect 6814 12484 6818 12540
rect 6818 12484 6874 12540
rect 6874 12484 6878 12540
rect 6814 12480 6878 12484
rect 10322 12540 10386 12544
rect 10322 12484 10326 12540
rect 10326 12484 10382 12540
rect 10382 12484 10386 12540
rect 10322 12480 10386 12484
rect 10402 12540 10466 12544
rect 10402 12484 10406 12540
rect 10406 12484 10462 12540
rect 10462 12484 10466 12540
rect 10402 12480 10466 12484
rect 10482 12540 10546 12544
rect 10482 12484 10486 12540
rect 10486 12484 10542 12540
rect 10542 12484 10546 12540
rect 10482 12480 10546 12484
rect 10562 12540 10626 12544
rect 10562 12484 10566 12540
rect 10566 12484 10622 12540
rect 10622 12484 10626 12540
rect 10562 12480 10626 12484
rect 14070 12540 14134 12544
rect 14070 12484 14074 12540
rect 14074 12484 14130 12540
rect 14130 12484 14134 12540
rect 14070 12480 14134 12484
rect 14150 12540 14214 12544
rect 14150 12484 14154 12540
rect 14154 12484 14210 12540
rect 14210 12484 14214 12540
rect 14150 12480 14214 12484
rect 14230 12540 14294 12544
rect 14230 12484 14234 12540
rect 14234 12484 14290 12540
rect 14290 12484 14294 12540
rect 14230 12480 14294 12484
rect 14310 12540 14374 12544
rect 14310 12484 14314 12540
rect 14314 12484 14370 12540
rect 14370 12484 14374 12540
rect 14310 12480 14374 12484
rect 13676 12276 13740 12340
rect 3924 12200 3988 12204
rect 3924 12144 3938 12200
rect 3938 12144 3988 12200
rect 3924 12140 3988 12144
rect 10180 12140 10244 12204
rect 13676 12064 13740 12068
rect 13676 12008 13726 12064
rect 13726 12008 13740 12064
rect 13676 12004 13740 12008
rect 4700 11996 4764 12000
rect 4700 11940 4704 11996
rect 4704 11940 4760 11996
rect 4760 11940 4764 11996
rect 4700 11936 4764 11940
rect 4780 11996 4844 12000
rect 4780 11940 4784 11996
rect 4784 11940 4840 11996
rect 4840 11940 4844 11996
rect 4780 11936 4844 11940
rect 4860 11996 4924 12000
rect 4860 11940 4864 11996
rect 4864 11940 4920 11996
rect 4920 11940 4924 11996
rect 4860 11936 4924 11940
rect 4940 11996 5004 12000
rect 4940 11940 4944 11996
rect 4944 11940 5000 11996
rect 5000 11940 5004 11996
rect 4940 11936 5004 11940
rect 8448 11996 8512 12000
rect 8448 11940 8452 11996
rect 8452 11940 8508 11996
rect 8508 11940 8512 11996
rect 8448 11936 8512 11940
rect 8528 11996 8592 12000
rect 8528 11940 8532 11996
rect 8532 11940 8588 11996
rect 8588 11940 8592 11996
rect 8528 11936 8592 11940
rect 8608 11996 8672 12000
rect 8608 11940 8612 11996
rect 8612 11940 8668 11996
rect 8668 11940 8672 11996
rect 8608 11936 8672 11940
rect 8688 11996 8752 12000
rect 8688 11940 8692 11996
rect 8692 11940 8748 11996
rect 8748 11940 8752 11996
rect 8688 11936 8752 11940
rect 12196 11996 12260 12000
rect 12196 11940 12200 11996
rect 12200 11940 12256 11996
rect 12256 11940 12260 11996
rect 12196 11936 12260 11940
rect 12276 11996 12340 12000
rect 12276 11940 12280 11996
rect 12280 11940 12336 11996
rect 12336 11940 12340 11996
rect 12276 11936 12340 11940
rect 12356 11996 12420 12000
rect 12356 11940 12360 11996
rect 12360 11940 12416 11996
rect 12416 11940 12420 11996
rect 12356 11936 12420 11940
rect 12436 11996 12500 12000
rect 12436 11940 12440 11996
rect 12440 11940 12496 11996
rect 12496 11940 12500 11996
rect 12436 11936 12500 11940
rect 12940 11868 13004 11932
rect 13860 11928 13924 11932
rect 13860 11872 13874 11928
rect 13874 11872 13924 11928
rect 13860 11868 13924 11872
rect 2826 11452 2890 11456
rect 2826 11396 2830 11452
rect 2830 11396 2886 11452
rect 2886 11396 2890 11452
rect 2826 11392 2890 11396
rect 2906 11452 2970 11456
rect 2906 11396 2910 11452
rect 2910 11396 2966 11452
rect 2966 11396 2970 11452
rect 2906 11392 2970 11396
rect 2986 11452 3050 11456
rect 2986 11396 2990 11452
rect 2990 11396 3046 11452
rect 3046 11396 3050 11452
rect 2986 11392 3050 11396
rect 3066 11452 3130 11456
rect 3066 11396 3070 11452
rect 3070 11396 3126 11452
rect 3126 11396 3130 11452
rect 3066 11392 3130 11396
rect 6574 11452 6638 11456
rect 6574 11396 6578 11452
rect 6578 11396 6634 11452
rect 6634 11396 6638 11452
rect 6574 11392 6638 11396
rect 6654 11452 6718 11456
rect 6654 11396 6658 11452
rect 6658 11396 6714 11452
rect 6714 11396 6718 11452
rect 6654 11392 6718 11396
rect 6734 11452 6798 11456
rect 6734 11396 6738 11452
rect 6738 11396 6794 11452
rect 6794 11396 6798 11452
rect 6734 11392 6798 11396
rect 6814 11452 6878 11456
rect 6814 11396 6818 11452
rect 6818 11396 6874 11452
rect 6874 11396 6878 11452
rect 6814 11392 6878 11396
rect 10322 11452 10386 11456
rect 10322 11396 10326 11452
rect 10326 11396 10382 11452
rect 10382 11396 10386 11452
rect 10322 11392 10386 11396
rect 10402 11452 10466 11456
rect 10402 11396 10406 11452
rect 10406 11396 10462 11452
rect 10462 11396 10466 11452
rect 10402 11392 10466 11396
rect 10482 11452 10546 11456
rect 10482 11396 10486 11452
rect 10486 11396 10542 11452
rect 10542 11396 10546 11452
rect 10482 11392 10546 11396
rect 10562 11452 10626 11456
rect 10562 11396 10566 11452
rect 10566 11396 10622 11452
rect 10622 11396 10626 11452
rect 10562 11392 10626 11396
rect 14070 11452 14134 11456
rect 14070 11396 14074 11452
rect 14074 11396 14130 11452
rect 14130 11396 14134 11452
rect 14070 11392 14134 11396
rect 14150 11452 14214 11456
rect 14150 11396 14154 11452
rect 14154 11396 14210 11452
rect 14210 11396 14214 11452
rect 14150 11392 14214 11396
rect 14230 11452 14294 11456
rect 14230 11396 14234 11452
rect 14234 11396 14290 11452
rect 14290 11396 14294 11452
rect 14230 11392 14294 11396
rect 14310 11452 14374 11456
rect 14310 11396 14314 11452
rect 14314 11396 14370 11452
rect 14370 11396 14374 11452
rect 14310 11392 14374 11396
rect 3372 11324 3436 11388
rect 13860 11052 13924 11116
rect 15148 11052 15212 11116
rect 4700 10908 4764 10912
rect 4700 10852 4704 10908
rect 4704 10852 4760 10908
rect 4760 10852 4764 10908
rect 4700 10848 4764 10852
rect 4780 10908 4844 10912
rect 4780 10852 4784 10908
rect 4784 10852 4840 10908
rect 4840 10852 4844 10908
rect 4780 10848 4844 10852
rect 4860 10908 4924 10912
rect 4860 10852 4864 10908
rect 4864 10852 4920 10908
rect 4920 10852 4924 10908
rect 4860 10848 4924 10852
rect 4940 10908 5004 10912
rect 4940 10852 4944 10908
rect 4944 10852 5000 10908
rect 5000 10852 5004 10908
rect 4940 10848 5004 10852
rect 8448 10908 8512 10912
rect 8448 10852 8452 10908
rect 8452 10852 8508 10908
rect 8508 10852 8512 10908
rect 8448 10848 8512 10852
rect 8528 10908 8592 10912
rect 8528 10852 8532 10908
rect 8532 10852 8588 10908
rect 8588 10852 8592 10908
rect 8528 10848 8592 10852
rect 8608 10908 8672 10912
rect 8608 10852 8612 10908
rect 8612 10852 8668 10908
rect 8668 10852 8672 10908
rect 8608 10848 8672 10852
rect 8688 10908 8752 10912
rect 8688 10852 8692 10908
rect 8692 10852 8748 10908
rect 8748 10852 8752 10908
rect 8688 10848 8752 10852
rect 12196 10908 12260 10912
rect 12196 10852 12200 10908
rect 12200 10852 12256 10908
rect 12256 10852 12260 10908
rect 12196 10848 12260 10852
rect 12276 10908 12340 10912
rect 12276 10852 12280 10908
rect 12280 10852 12336 10908
rect 12336 10852 12340 10908
rect 12276 10848 12340 10852
rect 12356 10908 12420 10912
rect 12356 10852 12360 10908
rect 12360 10852 12416 10908
rect 12416 10852 12420 10908
rect 12356 10848 12420 10852
rect 12436 10908 12500 10912
rect 12436 10852 12440 10908
rect 12440 10852 12496 10908
rect 12496 10852 12500 10908
rect 12436 10848 12500 10852
rect 2826 10364 2890 10368
rect 2826 10308 2830 10364
rect 2830 10308 2886 10364
rect 2886 10308 2890 10364
rect 2826 10304 2890 10308
rect 2906 10364 2970 10368
rect 2906 10308 2910 10364
rect 2910 10308 2966 10364
rect 2966 10308 2970 10364
rect 2906 10304 2970 10308
rect 2986 10364 3050 10368
rect 2986 10308 2990 10364
rect 2990 10308 3046 10364
rect 3046 10308 3050 10364
rect 2986 10304 3050 10308
rect 3066 10364 3130 10368
rect 3066 10308 3070 10364
rect 3070 10308 3126 10364
rect 3126 10308 3130 10364
rect 3066 10304 3130 10308
rect 6574 10364 6638 10368
rect 6574 10308 6578 10364
rect 6578 10308 6634 10364
rect 6634 10308 6638 10364
rect 6574 10304 6638 10308
rect 6654 10364 6718 10368
rect 6654 10308 6658 10364
rect 6658 10308 6714 10364
rect 6714 10308 6718 10364
rect 6654 10304 6718 10308
rect 6734 10364 6798 10368
rect 6734 10308 6738 10364
rect 6738 10308 6794 10364
rect 6794 10308 6798 10364
rect 6734 10304 6798 10308
rect 6814 10364 6878 10368
rect 6814 10308 6818 10364
rect 6818 10308 6874 10364
rect 6874 10308 6878 10364
rect 6814 10304 6878 10308
rect 10322 10364 10386 10368
rect 10322 10308 10326 10364
rect 10326 10308 10382 10364
rect 10382 10308 10386 10364
rect 10322 10304 10386 10308
rect 10402 10364 10466 10368
rect 10402 10308 10406 10364
rect 10406 10308 10462 10364
rect 10462 10308 10466 10364
rect 10402 10304 10466 10308
rect 10482 10364 10546 10368
rect 10482 10308 10486 10364
rect 10486 10308 10542 10364
rect 10542 10308 10546 10364
rect 10482 10304 10546 10308
rect 10562 10364 10626 10368
rect 10562 10308 10566 10364
rect 10566 10308 10622 10364
rect 10622 10308 10626 10364
rect 10562 10304 10626 10308
rect 14070 10364 14134 10368
rect 14070 10308 14074 10364
rect 14074 10308 14130 10364
rect 14130 10308 14134 10364
rect 14070 10304 14134 10308
rect 14150 10364 14214 10368
rect 14150 10308 14154 10364
rect 14154 10308 14210 10364
rect 14210 10308 14214 10364
rect 14150 10304 14214 10308
rect 14230 10364 14294 10368
rect 14230 10308 14234 10364
rect 14234 10308 14290 10364
rect 14290 10308 14294 10364
rect 14230 10304 14294 10308
rect 14310 10364 14374 10368
rect 14310 10308 14314 10364
rect 14314 10308 14370 10364
rect 14370 10308 14374 10364
rect 14310 10304 14374 10308
rect 11284 9964 11348 10028
rect 4700 9820 4764 9824
rect 4700 9764 4704 9820
rect 4704 9764 4760 9820
rect 4760 9764 4764 9820
rect 4700 9760 4764 9764
rect 4780 9820 4844 9824
rect 4780 9764 4784 9820
rect 4784 9764 4840 9820
rect 4840 9764 4844 9820
rect 4780 9760 4844 9764
rect 4860 9820 4924 9824
rect 4860 9764 4864 9820
rect 4864 9764 4920 9820
rect 4920 9764 4924 9820
rect 4860 9760 4924 9764
rect 4940 9820 5004 9824
rect 4940 9764 4944 9820
rect 4944 9764 5000 9820
rect 5000 9764 5004 9820
rect 4940 9760 5004 9764
rect 8448 9820 8512 9824
rect 8448 9764 8452 9820
rect 8452 9764 8508 9820
rect 8508 9764 8512 9820
rect 8448 9760 8512 9764
rect 8528 9820 8592 9824
rect 8528 9764 8532 9820
rect 8532 9764 8588 9820
rect 8588 9764 8592 9820
rect 8528 9760 8592 9764
rect 8608 9820 8672 9824
rect 8608 9764 8612 9820
rect 8612 9764 8668 9820
rect 8668 9764 8672 9820
rect 8608 9760 8672 9764
rect 8688 9820 8752 9824
rect 8688 9764 8692 9820
rect 8692 9764 8748 9820
rect 8748 9764 8752 9820
rect 8688 9760 8752 9764
rect 12196 9820 12260 9824
rect 12196 9764 12200 9820
rect 12200 9764 12256 9820
rect 12256 9764 12260 9820
rect 12196 9760 12260 9764
rect 12276 9820 12340 9824
rect 12276 9764 12280 9820
rect 12280 9764 12336 9820
rect 12336 9764 12340 9820
rect 12276 9760 12340 9764
rect 12356 9820 12420 9824
rect 12356 9764 12360 9820
rect 12360 9764 12416 9820
rect 12416 9764 12420 9820
rect 12356 9760 12420 9764
rect 12436 9820 12500 9824
rect 12436 9764 12440 9820
rect 12440 9764 12496 9820
rect 12496 9764 12500 9820
rect 12436 9760 12500 9764
rect 13492 9692 13556 9756
rect 3372 9556 3436 9620
rect 13860 9420 13924 9484
rect 2826 9276 2890 9280
rect 2826 9220 2830 9276
rect 2830 9220 2886 9276
rect 2886 9220 2890 9276
rect 2826 9216 2890 9220
rect 2906 9276 2970 9280
rect 2906 9220 2910 9276
rect 2910 9220 2966 9276
rect 2966 9220 2970 9276
rect 2906 9216 2970 9220
rect 2986 9276 3050 9280
rect 2986 9220 2990 9276
rect 2990 9220 3046 9276
rect 3046 9220 3050 9276
rect 2986 9216 3050 9220
rect 3066 9276 3130 9280
rect 3066 9220 3070 9276
rect 3070 9220 3126 9276
rect 3126 9220 3130 9276
rect 3066 9216 3130 9220
rect 6574 9276 6638 9280
rect 6574 9220 6578 9276
rect 6578 9220 6634 9276
rect 6634 9220 6638 9276
rect 6574 9216 6638 9220
rect 6654 9276 6718 9280
rect 6654 9220 6658 9276
rect 6658 9220 6714 9276
rect 6714 9220 6718 9276
rect 6654 9216 6718 9220
rect 6734 9276 6798 9280
rect 6734 9220 6738 9276
rect 6738 9220 6794 9276
rect 6794 9220 6798 9276
rect 6734 9216 6798 9220
rect 6814 9276 6878 9280
rect 6814 9220 6818 9276
rect 6818 9220 6874 9276
rect 6874 9220 6878 9276
rect 6814 9216 6878 9220
rect 10322 9276 10386 9280
rect 10322 9220 10326 9276
rect 10326 9220 10382 9276
rect 10382 9220 10386 9276
rect 10322 9216 10386 9220
rect 10402 9276 10466 9280
rect 10402 9220 10406 9276
rect 10406 9220 10462 9276
rect 10462 9220 10466 9276
rect 10402 9216 10466 9220
rect 10482 9276 10546 9280
rect 10482 9220 10486 9276
rect 10486 9220 10542 9276
rect 10542 9220 10546 9276
rect 10482 9216 10546 9220
rect 10562 9276 10626 9280
rect 10562 9220 10566 9276
rect 10566 9220 10622 9276
rect 10622 9220 10626 9276
rect 10562 9216 10626 9220
rect 14070 9276 14134 9280
rect 14070 9220 14074 9276
rect 14074 9220 14130 9276
rect 14130 9220 14134 9276
rect 14070 9216 14134 9220
rect 14150 9276 14214 9280
rect 14150 9220 14154 9276
rect 14154 9220 14210 9276
rect 14210 9220 14214 9276
rect 14150 9216 14214 9220
rect 14230 9276 14294 9280
rect 14230 9220 14234 9276
rect 14234 9220 14290 9276
rect 14290 9220 14294 9276
rect 14230 9216 14294 9220
rect 14310 9276 14374 9280
rect 14310 9220 14314 9276
rect 14314 9220 14370 9276
rect 14370 9220 14374 9276
rect 14310 9216 14374 9220
rect 12572 9012 12636 9076
rect 9628 8876 9692 8940
rect 4700 8732 4764 8736
rect 4700 8676 4704 8732
rect 4704 8676 4760 8732
rect 4760 8676 4764 8732
rect 4700 8672 4764 8676
rect 4780 8732 4844 8736
rect 4780 8676 4784 8732
rect 4784 8676 4840 8732
rect 4840 8676 4844 8732
rect 4780 8672 4844 8676
rect 4860 8732 4924 8736
rect 4860 8676 4864 8732
rect 4864 8676 4920 8732
rect 4920 8676 4924 8732
rect 4860 8672 4924 8676
rect 4940 8732 5004 8736
rect 4940 8676 4944 8732
rect 4944 8676 5000 8732
rect 5000 8676 5004 8732
rect 4940 8672 5004 8676
rect 8448 8732 8512 8736
rect 8448 8676 8452 8732
rect 8452 8676 8508 8732
rect 8508 8676 8512 8732
rect 8448 8672 8512 8676
rect 8528 8732 8592 8736
rect 8528 8676 8532 8732
rect 8532 8676 8588 8732
rect 8588 8676 8592 8732
rect 8528 8672 8592 8676
rect 8608 8732 8672 8736
rect 8608 8676 8612 8732
rect 8612 8676 8668 8732
rect 8668 8676 8672 8732
rect 8608 8672 8672 8676
rect 8688 8732 8752 8736
rect 8688 8676 8692 8732
rect 8692 8676 8748 8732
rect 8748 8676 8752 8732
rect 8688 8672 8752 8676
rect 12196 8732 12260 8736
rect 12196 8676 12200 8732
rect 12200 8676 12256 8732
rect 12256 8676 12260 8732
rect 12196 8672 12260 8676
rect 12276 8732 12340 8736
rect 12276 8676 12280 8732
rect 12280 8676 12336 8732
rect 12336 8676 12340 8732
rect 12276 8672 12340 8676
rect 12356 8732 12420 8736
rect 12356 8676 12360 8732
rect 12360 8676 12416 8732
rect 12416 8676 12420 8732
rect 12356 8672 12420 8676
rect 12436 8732 12500 8736
rect 12436 8676 12440 8732
rect 12440 8676 12496 8732
rect 12496 8676 12500 8732
rect 12436 8672 12500 8676
rect 2826 8188 2890 8192
rect 2826 8132 2830 8188
rect 2830 8132 2886 8188
rect 2886 8132 2890 8188
rect 2826 8128 2890 8132
rect 2906 8188 2970 8192
rect 2906 8132 2910 8188
rect 2910 8132 2966 8188
rect 2966 8132 2970 8188
rect 2906 8128 2970 8132
rect 2986 8188 3050 8192
rect 2986 8132 2990 8188
rect 2990 8132 3046 8188
rect 3046 8132 3050 8188
rect 2986 8128 3050 8132
rect 3066 8188 3130 8192
rect 3066 8132 3070 8188
rect 3070 8132 3126 8188
rect 3126 8132 3130 8188
rect 3066 8128 3130 8132
rect 6574 8188 6638 8192
rect 6574 8132 6578 8188
rect 6578 8132 6634 8188
rect 6634 8132 6638 8188
rect 6574 8128 6638 8132
rect 6654 8188 6718 8192
rect 6654 8132 6658 8188
rect 6658 8132 6714 8188
rect 6714 8132 6718 8188
rect 6654 8128 6718 8132
rect 6734 8188 6798 8192
rect 6734 8132 6738 8188
rect 6738 8132 6794 8188
rect 6794 8132 6798 8188
rect 6734 8128 6798 8132
rect 6814 8188 6878 8192
rect 6814 8132 6818 8188
rect 6818 8132 6874 8188
rect 6874 8132 6878 8188
rect 6814 8128 6878 8132
rect 10322 8188 10386 8192
rect 10322 8132 10326 8188
rect 10326 8132 10382 8188
rect 10382 8132 10386 8188
rect 10322 8128 10386 8132
rect 10402 8188 10466 8192
rect 10402 8132 10406 8188
rect 10406 8132 10462 8188
rect 10462 8132 10466 8188
rect 10402 8128 10466 8132
rect 10482 8188 10546 8192
rect 10482 8132 10486 8188
rect 10486 8132 10542 8188
rect 10542 8132 10546 8188
rect 10482 8128 10546 8132
rect 10562 8188 10626 8192
rect 10562 8132 10566 8188
rect 10566 8132 10622 8188
rect 10622 8132 10626 8188
rect 10562 8128 10626 8132
rect 14070 8188 14134 8192
rect 14070 8132 14074 8188
rect 14074 8132 14130 8188
rect 14130 8132 14134 8188
rect 14070 8128 14134 8132
rect 14150 8188 14214 8192
rect 14150 8132 14154 8188
rect 14154 8132 14210 8188
rect 14210 8132 14214 8188
rect 14150 8128 14214 8132
rect 14230 8188 14294 8192
rect 14230 8132 14234 8188
rect 14234 8132 14290 8188
rect 14290 8132 14294 8188
rect 14230 8128 14294 8132
rect 14310 8188 14374 8192
rect 14310 8132 14314 8188
rect 14314 8132 14370 8188
rect 14370 8132 14374 8188
rect 14310 8128 14374 8132
rect 4700 7644 4764 7648
rect 4700 7588 4704 7644
rect 4704 7588 4760 7644
rect 4760 7588 4764 7644
rect 4700 7584 4764 7588
rect 4780 7644 4844 7648
rect 4780 7588 4784 7644
rect 4784 7588 4840 7644
rect 4840 7588 4844 7644
rect 4780 7584 4844 7588
rect 4860 7644 4924 7648
rect 4860 7588 4864 7644
rect 4864 7588 4920 7644
rect 4920 7588 4924 7644
rect 4860 7584 4924 7588
rect 4940 7644 5004 7648
rect 4940 7588 4944 7644
rect 4944 7588 5000 7644
rect 5000 7588 5004 7644
rect 4940 7584 5004 7588
rect 8448 7644 8512 7648
rect 8448 7588 8452 7644
rect 8452 7588 8508 7644
rect 8508 7588 8512 7644
rect 8448 7584 8512 7588
rect 8528 7644 8592 7648
rect 8528 7588 8532 7644
rect 8532 7588 8588 7644
rect 8588 7588 8592 7644
rect 8528 7584 8592 7588
rect 8608 7644 8672 7648
rect 8608 7588 8612 7644
rect 8612 7588 8668 7644
rect 8668 7588 8672 7644
rect 8608 7584 8672 7588
rect 8688 7644 8752 7648
rect 8688 7588 8692 7644
rect 8692 7588 8748 7644
rect 8748 7588 8752 7644
rect 8688 7584 8752 7588
rect 12196 7644 12260 7648
rect 12196 7588 12200 7644
rect 12200 7588 12256 7644
rect 12256 7588 12260 7644
rect 12196 7584 12260 7588
rect 12276 7644 12340 7648
rect 12276 7588 12280 7644
rect 12280 7588 12336 7644
rect 12336 7588 12340 7644
rect 12276 7584 12340 7588
rect 12356 7644 12420 7648
rect 12356 7588 12360 7644
rect 12360 7588 12416 7644
rect 12416 7588 12420 7644
rect 12356 7584 12420 7588
rect 12436 7644 12500 7648
rect 12436 7588 12440 7644
rect 12440 7588 12496 7644
rect 12496 7588 12500 7644
rect 12436 7584 12500 7588
rect 2826 7100 2890 7104
rect 2826 7044 2830 7100
rect 2830 7044 2886 7100
rect 2886 7044 2890 7100
rect 2826 7040 2890 7044
rect 2906 7100 2970 7104
rect 2906 7044 2910 7100
rect 2910 7044 2966 7100
rect 2966 7044 2970 7100
rect 2906 7040 2970 7044
rect 2986 7100 3050 7104
rect 2986 7044 2990 7100
rect 2990 7044 3046 7100
rect 3046 7044 3050 7100
rect 2986 7040 3050 7044
rect 3066 7100 3130 7104
rect 3066 7044 3070 7100
rect 3070 7044 3126 7100
rect 3126 7044 3130 7100
rect 3066 7040 3130 7044
rect 6574 7100 6638 7104
rect 6574 7044 6578 7100
rect 6578 7044 6634 7100
rect 6634 7044 6638 7100
rect 6574 7040 6638 7044
rect 6654 7100 6718 7104
rect 6654 7044 6658 7100
rect 6658 7044 6714 7100
rect 6714 7044 6718 7100
rect 6654 7040 6718 7044
rect 6734 7100 6798 7104
rect 6734 7044 6738 7100
rect 6738 7044 6794 7100
rect 6794 7044 6798 7100
rect 6734 7040 6798 7044
rect 6814 7100 6878 7104
rect 6814 7044 6818 7100
rect 6818 7044 6874 7100
rect 6874 7044 6878 7100
rect 6814 7040 6878 7044
rect 10322 7100 10386 7104
rect 10322 7044 10326 7100
rect 10326 7044 10382 7100
rect 10382 7044 10386 7100
rect 10322 7040 10386 7044
rect 10402 7100 10466 7104
rect 10402 7044 10406 7100
rect 10406 7044 10462 7100
rect 10462 7044 10466 7100
rect 10402 7040 10466 7044
rect 10482 7100 10546 7104
rect 10482 7044 10486 7100
rect 10486 7044 10542 7100
rect 10542 7044 10546 7100
rect 10482 7040 10546 7044
rect 10562 7100 10626 7104
rect 10562 7044 10566 7100
rect 10566 7044 10622 7100
rect 10622 7044 10626 7100
rect 10562 7040 10626 7044
rect 14070 7100 14134 7104
rect 14070 7044 14074 7100
rect 14074 7044 14130 7100
rect 14130 7044 14134 7100
rect 14070 7040 14134 7044
rect 14150 7100 14214 7104
rect 14150 7044 14154 7100
rect 14154 7044 14210 7100
rect 14210 7044 14214 7100
rect 14150 7040 14214 7044
rect 14230 7100 14294 7104
rect 14230 7044 14234 7100
rect 14234 7044 14290 7100
rect 14290 7044 14294 7100
rect 14230 7040 14294 7044
rect 14310 7100 14374 7104
rect 14310 7044 14314 7100
rect 14314 7044 14370 7100
rect 14370 7044 14374 7100
rect 14310 7040 14374 7044
rect 13124 6700 13188 6764
rect 2268 6564 2332 6628
rect 3556 6564 3620 6628
rect 4700 6556 4764 6560
rect 4700 6500 4704 6556
rect 4704 6500 4760 6556
rect 4760 6500 4764 6556
rect 4700 6496 4764 6500
rect 4780 6556 4844 6560
rect 4780 6500 4784 6556
rect 4784 6500 4840 6556
rect 4840 6500 4844 6556
rect 4780 6496 4844 6500
rect 4860 6556 4924 6560
rect 4860 6500 4864 6556
rect 4864 6500 4920 6556
rect 4920 6500 4924 6556
rect 4860 6496 4924 6500
rect 4940 6556 5004 6560
rect 4940 6500 4944 6556
rect 4944 6500 5000 6556
rect 5000 6500 5004 6556
rect 4940 6496 5004 6500
rect 8448 6556 8512 6560
rect 8448 6500 8452 6556
rect 8452 6500 8508 6556
rect 8508 6500 8512 6556
rect 8448 6496 8512 6500
rect 8528 6556 8592 6560
rect 8528 6500 8532 6556
rect 8532 6500 8588 6556
rect 8588 6500 8592 6556
rect 8528 6496 8592 6500
rect 8608 6556 8672 6560
rect 8608 6500 8612 6556
rect 8612 6500 8668 6556
rect 8668 6500 8672 6556
rect 8608 6496 8672 6500
rect 8688 6556 8752 6560
rect 8688 6500 8692 6556
rect 8692 6500 8748 6556
rect 8748 6500 8752 6556
rect 8688 6496 8752 6500
rect 12196 6556 12260 6560
rect 12196 6500 12200 6556
rect 12200 6500 12256 6556
rect 12256 6500 12260 6556
rect 12196 6496 12260 6500
rect 12276 6556 12340 6560
rect 12276 6500 12280 6556
rect 12280 6500 12336 6556
rect 12336 6500 12340 6556
rect 12276 6496 12340 6500
rect 12356 6556 12420 6560
rect 12356 6500 12360 6556
rect 12360 6500 12416 6556
rect 12416 6500 12420 6556
rect 12356 6496 12420 6500
rect 12436 6556 12500 6560
rect 12436 6500 12440 6556
rect 12440 6500 12496 6556
rect 12496 6500 12500 6556
rect 12436 6496 12500 6500
rect 11652 6292 11716 6356
rect 2636 6156 2700 6220
rect 9996 6156 10060 6220
rect 13860 6156 13924 6220
rect 2826 6012 2890 6016
rect 2826 5956 2830 6012
rect 2830 5956 2886 6012
rect 2886 5956 2890 6012
rect 2826 5952 2890 5956
rect 2906 6012 2970 6016
rect 2906 5956 2910 6012
rect 2910 5956 2966 6012
rect 2966 5956 2970 6012
rect 2906 5952 2970 5956
rect 2986 6012 3050 6016
rect 2986 5956 2990 6012
rect 2990 5956 3046 6012
rect 3046 5956 3050 6012
rect 2986 5952 3050 5956
rect 3066 6012 3130 6016
rect 3066 5956 3070 6012
rect 3070 5956 3126 6012
rect 3126 5956 3130 6012
rect 3066 5952 3130 5956
rect 6574 6012 6638 6016
rect 6574 5956 6578 6012
rect 6578 5956 6634 6012
rect 6634 5956 6638 6012
rect 6574 5952 6638 5956
rect 6654 6012 6718 6016
rect 6654 5956 6658 6012
rect 6658 5956 6714 6012
rect 6714 5956 6718 6012
rect 6654 5952 6718 5956
rect 6734 6012 6798 6016
rect 6734 5956 6738 6012
rect 6738 5956 6794 6012
rect 6794 5956 6798 6012
rect 6734 5952 6798 5956
rect 6814 6012 6878 6016
rect 6814 5956 6818 6012
rect 6818 5956 6874 6012
rect 6874 5956 6878 6012
rect 6814 5952 6878 5956
rect 10322 6012 10386 6016
rect 10322 5956 10326 6012
rect 10326 5956 10382 6012
rect 10382 5956 10386 6012
rect 10322 5952 10386 5956
rect 10402 6012 10466 6016
rect 10402 5956 10406 6012
rect 10406 5956 10462 6012
rect 10462 5956 10466 6012
rect 10402 5952 10466 5956
rect 10482 6012 10546 6016
rect 10482 5956 10486 6012
rect 10486 5956 10542 6012
rect 10542 5956 10546 6012
rect 10482 5952 10546 5956
rect 10562 6012 10626 6016
rect 10562 5956 10566 6012
rect 10566 5956 10622 6012
rect 10622 5956 10626 6012
rect 10562 5952 10626 5956
rect 14070 6012 14134 6016
rect 14070 5956 14074 6012
rect 14074 5956 14130 6012
rect 14130 5956 14134 6012
rect 14070 5952 14134 5956
rect 14150 6012 14214 6016
rect 14150 5956 14154 6012
rect 14154 5956 14210 6012
rect 14210 5956 14214 6012
rect 14150 5952 14214 5956
rect 14230 6012 14294 6016
rect 14230 5956 14234 6012
rect 14234 5956 14290 6012
rect 14290 5956 14294 6012
rect 14230 5952 14294 5956
rect 14310 6012 14374 6016
rect 14310 5956 14314 6012
rect 14314 5956 14370 6012
rect 14370 5956 14374 6012
rect 14310 5952 14374 5956
rect 12572 5748 12636 5812
rect 14780 5748 14844 5812
rect 4700 5468 4764 5472
rect 4700 5412 4704 5468
rect 4704 5412 4760 5468
rect 4760 5412 4764 5468
rect 4700 5408 4764 5412
rect 4780 5468 4844 5472
rect 4780 5412 4784 5468
rect 4784 5412 4840 5468
rect 4840 5412 4844 5468
rect 4780 5408 4844 5412
rect 4860 5468 4924 5472
rect 4860 5412 4864 5468
rect 4864 5412 4920 5468
rect 4920 5412 4924 5468
rect 4860 5408 4924 5412
rect 4940 5468 5004 5472
rect 4940 5412 4944 5468
rect 4944 5412 5000 5468
rect 5000 5412 5004 5468
rect 4940 5408 5004 5412
rect 9996 5612 10060 5676
rect 10180 5476 10244 5540
rect 14596 5476 14660 5540
rect 8448 5468 8512 5472
rect 8448 5412 8452 5468
rect 8452 5412 8508 5468
rect 8508 5412 8512 5468
rect 8448 5408 8512 5412
rect 8528 5468 8592 5472
rect 8528 5412 8532 5468
rect 8532 5412 8588 5468
rect 8588 5412 8592 5468
rect 8528 5408 8592 5412
rect 8608 5468 8672 5472
rect 8608 5412 8612 5468
rect 8612 5412 8668 5468
rect 8668 5412 8672 5468
rect 8608 5408 8672 5412
rect 8688 5468 8752 5472
rect 8688 5412 8692 5468
rect 8692 5412 8748 5468
rect 8748 5412 8752 5468
rect 8688 5408 8752 5412
rect 12196 5468 12260 5472
rect 12196 5412 12200 5468
rect 12200 5412 12256 5468
rect 12256 5412 12260 5468
rect 12196 5408 12260 5412
rect 12276 5468 12340 5472
rect 12276 5412 12280 5468
rect 12280 5412 12336 5468
rect 12336 5412 12340 5468
rect 12276 5408 12340 5412
rect 12356 5468 12420 5472
rect 12356 5412 12360 5468
rect 12360 5412 12416 5468
rect 12416 5412 12420 5468
rect 12356 5408 12420 5412
rect 12436 5468 12500 5472
rect 12436 5412 12440 5468
rect 12440 5412 12496 5468
rect 12496 5412 12500 5468
rect 12436 5408 12500 5412
rect 10916 5340 10980 5404
rect 14964 5400 15028 5404
rect 14964 5344 15014 5400
rect 15014 5344 15028 5400
rect 14964 5340 15028 5344
rect 2268 5068 2332 5132
rect 12572 4932 12636 4996
rect 2826 4924 2890 4928
rect 2826 4868 2830 4924
rect 2830 4868 2886 4924
rect 2886 4868 2890 4924
rect 2826 4864 2890 4868
rect 2906 4924 2970 4928
rect 2906 4868 2910 4924
rect 2910 4868 2966 4924
rect 2966 4868 2970 4924
rect 2906 4864 2970 4868
rect 2986 4924 3050 4928
rect 2986 4868 2990 4924
rect 2990 4868 3046 4924
rect 3046 4868 3050 4924
rect 2986 4864 3050 4868
rect 3066 4924 3130 4928
rect 3066 4868 3070 4924
rect 3070 4868 3126 4924
rect 3126 4868 3130 4924
rect 3066 4864 3130 4868
rect 6574 4924 6638 4928
rect 6574 4868 6578 4924
rect 6578 4868 6634 4924
rect 6634 4868 6638 4924
rect 6574 4864 6638 4868
rect 6654 4924 6718 4928
rect 6654 4868 6658 4924
rect 6658 4868 6714 4924
rect 6714 4868 6718 4924
rect 6654 4864 6718 4868
rect 6734 4924 6798 4928
rect 6734 4868 6738 4924
rect 6738 4868 6794 4924
rect 6794 4868 6798 4924
rect 6734 4864 6798 4868
rect 6814 4924 6878 4928
rect 6814 4868 6818 4924
rect 6818 4868 6874 4924
rect 6874 4868 6878 4924
rect 6814 4864 6878 4868
rect 10322 4924 10386 4928
rect 10322 4868 10326 4924
rect 10326 4868 10382 4924
rect 10382 4868 10386 4924
rect 10322 4864 10386 4868
rect 10402 4924 10466 4928
rect 10402 4868 10406 4924
rect 10406 4868 10462 4924
rect 10462 4868 10466 4924
rect 10402 4864 10466 4868
rect 10482 4924 10546 4928
rect 10482 4868 10486 4924
rect 10486 4868 10542 4924
rect 10542 4868 10546 4924
rect 10482 4864 10546 4868
rect 10562 4924 10626 4928
rect 10562 4868 10566 4924
rect 10566 4868 10622 4924
rect 10622 4868 10626 4924
rect 10562 4864 10626 4868
rect 14070 4924 14134 4928
rect 14070 4868 14074 4924
rect 14074 4868 14130 4924
rect 14130 4868 14134 4924
rect 14070 4864 14134 4868
rect 14150 4924 14214 4928
rect 14150 4868 14154 4924
rect 14154 4868 14210 4924
rect 14210 4868 14214 4924
rect 14150 4864 14214 4868
rect 14230 4924 14294 4928
rect 14230 4868 14234 4924
rect 14234 4868 14290 4924
rect 14290 4868 14294 4924
rect 14230 4864 14294 4868
rect 14310 4924 14374 4928
rect 14310 4868 14314 4924
rect 14314 4868 14370 4924
rect 14370 4868 14374 4924
rect 14310 4864 14374 4868
rect 9812 4856 9876 4860
rect 9812 4800 9862 4856
rect 9862 4800 9876 4856
rect 9812 4796 9876 4800
rect 2636 4660 2700 4724
rect 4700 4380 4764 4384
rect 4700 4324 4704 4380
rect 4704 4324 4760 4380
rect 4760 4324 4764 4380
rect 4700 4320 4764 4324
rect 4780 4380 4844 4384
rect 4780 4324 4784 4380
rect 4784 4324 4840 4380
rect 4840 4324 4844 4380
rect 4780 4320 4844 4324
rect 4860 4380 4924 4384
rect 4860 4324 4864 4380
rect 4864 4324 4920 4380
rect 4920 4324 4924 4380
rect 4860 4320 4924 4324
rect 4940 4380 5004 4384
rect 4940 4324 4944 4380
rect 4944 4324 5000 4380
rect 5000 4324 5004 4380
rect 4940 4320 5004 4324
rect 8448 4380 8512 4384
rect 8448 4324 8452 4380
rect 8452 4324 8508 4380
rect 8508 4324 8512 4380
rect 8448 4320 8512 4324
rect 8528 4380 8592 4384
rect 8528 4324 8532 4380
rect 8532 4324 8588 4380
rect 8588 4324 8592 4380
rect 8528 4320 8592 4324
rect 8608 4380 8672 4384
rect 8608 4324 8612 4380
rect 8612 4324 8668 4380
rect 8668 4324 8672 4380
rect 8608 4320 8672 4324
rect 8688 4380 8752 4384
rect 8688 4324 8692 4380
rect 8692 4324 8748 4380
rect 8748 4324 8752 4380
rect 8688 4320 8752 4324
rect 5580 4252 5644 4316
rect 11100 4448 11164 4452
rect 11100 4392 11150 4448
rect 11150 4392 11164 4448
rect 11100 4388 11164 4392
rect 14596 4388 14660 4452
rect 12196 4380 12260 4384
rect 12196 4324 12200 4380
rect 12200 4324 12256 4380
rect 12256 4324 12260 4380
rect 12196 4320 12260 4324
rect 12276 4380 12340 4384
rect 12276 4324 12280 4380
rect 12280 4324 12336 4380
rect 12336 4324 12340 4380
rect 12276 4320 12340 4324
rect 12356 4380 12420 4384
rect 12356 4324 12360 4380
rect 12360 4324 12416 4380
rect 12416 4324 12420 4380
rect 12356 4320 12420 4324
rect 12436 4380 12500 4384
rect 12436 4324 12440 4380
rect 12440 4324 12496 4380
rect 12496 4324 12500 4380
rect 12436 4320 12500 4324
rect 11284 4312 11348 4316
rect 11284 4256 11298 4312
rect 11298 4256 11348 4312
rect 11284 4252 11348 4256
rect 9996 3980 10060 4044
rect 12020 3980 12084 4044
rect 14780 4040 14844 4044
rect 14780 3984 14830 4040
rect 14830 3984 14844 4040
rect 14780 3980 14844 3984
rect 2826 3836 2890 3840
rect 2826 3780 2830 3836
rect 2830 3780 2886 3836
rect 2886 3780 2890 3836
rect 2826 3776 2890 3780
rect 2906 3836 2970 3840
rect 2906 3780 2910 3836
rect 2910 3780 2966 3836
rect 2966 3780 2970 3836
rect 2906 3776 2970 3780
rect 2986 3836 3050 3840
rect 2986 3780 2990 3836
rect 2990 3780 3046 3836
rect 3046 3780 3050 3836
rect 2986 3776 3050 3780
rect 3066 3836 3130 3840
rect 3066 3780 3070 3836
rect 3070 3780 3126 3836
rect 3126 3780 3130 3836
rect 3066 3776 3130 3780
rect 6574 3836 6638 3840
rect 6574 3780 6578 3836
rect 6578 3780 6634 3836
rect 6634 3780 6638 3836
rect 6574 3776 6638 3780
rect 6654 3836 6718 3840
rect 6654 3780 6658 3836
rect 6658 3780 6714 3836
rect 6714 3780 6718 3836
rect 6654 3776 6718 3780
rect 6734 3836 6798 3840
rect 6734 3780 6738 3836
rect 6738 3780 6794 3836
rect 6794 3780 6798 3836
rect 6734 3776 6798 3780
rect 6814 3836 6878 3840
rect 6814 3780 6818 3836
rect 6818 3780 6874 3836
rect 6874 3780 6878 3836
rect 6814 3776 6878 3780
rect 10322 3836 10386 3840
rect 10322 3780 10326 3836
rect 10326 3780 10382 3836
rect 10382 3780 10386 3836
rect 10322 3776 10386 3780
rect 10402 3836 10466 3840
rect 10402 3780 10406 3836
rect 10406 3780 10462 3836
rect 10462 3780 10466 3836
rect 10402 3776 10466 3780
rect 10482 3836 10546 3840
rect 10482 3780 10486 3836
rect 10486 3780 10542 3836
rect 10542 3780 10546 3836
rect 10482 3776 10546 3780
rect 10562 3836 10626 3840
rect 10562 3780 10566 3836
rect 10566 3780 10622 3836
rect 10622 3780 10626 3836
rect 10562 3776 10626 3780
rect 11100 3708 11164 3772
rect 7236 3572 7300 3636
rect 14070 3836 14134 3840
rect 14070 3780 14074 3836
rect 14074 3780 14130 3836
rect 14130 3780 14134 3836
rect 14070 3776 14134 3780
rect 14150 3836 14214 3840
rect 14150 3780 14154 3836
rect 14154 3780 14210 3836
rect 14210 3780 14214 3836
rect 14150 3776 14214 3780
rect 14230 3836 14294 3840
rect 14230 3780 14234 3836
rect 14234 3780 14290 3836
rect 14290 3780 14294 3836
rect 14230 3776 14294 3780
rect 14310 3836 14374 3840
rect 14310 3780 14314 3836
rect 14314 3780 14370 3836
rect 14370 3780 14374 3836
rect 14310 3776 14374 3780
rect 5580 3360 5644 3364
rect 5580 3304 5594 3360
rect 5594 3304 5644 3360
rect 5580 3300 5644 3304
rect 4700 3292 4764 3296
rect 4700 3236 4704 3292
rect 4704 3236 4760 3292
rect 4760 3236 4764 3292
rect 4700 3232 4764 3236
rect 4780 3292 4844 3296
rect 4780 3236 4784 3292
rect 4784 3236 4840 3292
rect 4840 3236 4844 3292
rect 4780 3232 4844 3236
rect 4860 3292 4924 3296
rect 4860 3236 4864 3292
rect 4864 3236 4920 3292
rect 4920 3236 4924 3292
rect 4860 3232 4924 3236
rect 4940 3292 5004 3296
rect 4940 3236 4944 3292
rect 4944 3236 5000 3292
rect 5000 3236 5004 3292
rect 4940 3232 5004 3236
rect 8448 3292 8512 3296
rect 8448 3236 8452 3292
rect 8452 3236 8508 3292
rect 8508 3236 8512 3292
rect 8448 3232 8512 3236
rect 8528 3292 8592 3296
rect 8528 3236 8532 3292
rect 8532 3236 8588 3292
rect 8588 3236 8592 3292
rect 8528 3232 8592 3236
rect 8608 3292 8672 3296
rect 8608 3236 8612 3292
rect 8612 3236 8668 3292
rect 8668 3236 8672 3292
rect 8608 3232 8672 3236
rect 8688 3292 8752 3296
rect 8688 3236 8692 3292
rect 8692 3236 8748 3292
rect 8748 3236 8752 3292
rect 8688 3232 8752 3236
rect 12196 3292 12260 3296
rect 12196 3236 12200 3292
rect 12200 3236 12256 3292
rect 12256 3236 12260 3292
rect 12196 3232 12260 3236
rect 12276 3292 12340 3296
rect 12276 3236 12280 3292
rect 12280 3236 12336 3292
rect 12336 3236 12340 3292
rect 12276 3232 12340 3236
rect 12356 3292 12420 3296
rect 12356 3236 12360 3292
rect 12360 3236 12416 3292
rect 12416 3236 12420 3292
rect 12356 3232 12420 3236
rect 12436 3292 12500 3296
rect 12436 3236 12440 3292
rect 12440 3236 12496 3292
rect 12496 3236 12500 3292
rect 12436 3232 12500 3236
rect 9812 3164 9876 3228
rect 10916 3164 10980 3228
rect 11652 3028 11716 3092
rect 7236 2892 7300 2956
rect 13860 2952 13924 2956
rect 13860 2896 13874 2952
rect 13874 2896 13924 2952
rect 13860 2892 13924 2896
rect 10180 2756 10244 2820
rect 2826 2748 2890 2752
rect 2826 2692 2830 2748
rect 2830 2692 2886 2748
rect 2886 2692 2890 2748
rect 2826 2688 2890 2692
rect 2906 2748 2970 2752
rect 2906 2692 2910 2748
rect 2910 2692 2966 2748
rect 2966 2692 2970 2748
rect 2906 2688 2970 2692
rect 2986 2748 3050 2752
rect 2986 2692 2990 2748
rect 2990 2692 3046 2748
rect 3046 2692 3050 2748
rect 2986 2688 3050 2692
rect 3066 2748 3130 2752
rect 3066 2692 3070 2748
rect 3070 2692 3126 2748
rect 3126 2692 3130 2748
rect 3066 2688 3130 2692
rect 6574 2748 6638 2752
rect 6574 2692 6578 2748
rect 6578 2692 6634 2748
rect 6634 2692 6638 2748
rect 6574 2688 6638 2692
rect 6654 2748 6718 2752
rect 6654 2692 6658 2748
rect 6658 2692 6714 2748
rect 6714 2692 6718 2748
rect 6654 2688 6718 2692
rect 6734 2748 6798 2752
rect 6734 2692 6738 2748
rect 6738 2692 6794 2748
rect 6794 2692 6798 2748
rect 6734 2688 6798 2692
rect 6814 2748 6878 2752
rect 6814 2692 6818 2748
rect 6818 2692 6874 2748
rect 6874 2692 6878 2748
rect 6814 2688 6878 2692
rect 10322 2748 10386 2752
rect 10322 2692 10326 2748
rect 10326 2692 10382 2748
rect 10382 2692 10386 2748
rect 10322 2688 10386 2692
rect 10402 2748 10466 2752
rect 10402 2692 10406 2748
rect 10406 2692 10462 2748
rect 10462 2692 10466 2748
rect 10402 2688 10466 2692
rect 10482 2748 10546 2752
rect 10482 2692 10486 2748
rect 10486 2692 10542 2748
rect 10542 2692 10546 2748
rect 10482 2688 10546 2692
rect 10562 2748 10626 2752
rect 10562 2692 10566 2748
rect 10566 2692 10622 2748
rect 10622 2692 10626 2748
rect 10562 2688 10626 2692
rect 14070 2748 14134 2752
rect 14070 2692 14074 2748
rect 14074 2692 14130 2748
rect 14130 2692 14134 2748
rect 14070 2688 14134 2692
rect 14150 2748 14214 2752
rect 14150 2692 14154 2748
rect 14154 2692 14210 2748
rect 14210 2692 14214 2748
rect 14150 2688 14214 2692
rect 14230 2748 14294 2752
rect 14230 2692 14234 2748
rect 14234 2692 14290 2748
rect 14290 2692 14294 2748
rect 14230 2688 14294 2692
rect 14310 2748 14374 2752
rect 14310 2692 14314 2748
rect 14314 2692 14370 2748
rect 14370 2692 14374 2748
rect 14310 2688 14374 2692
rect 13676 2484 13740 2548
rect 3924 2348 3988 2412
rect 4700 2204 4764 2208
rect 4700 2148 4704 2204
rect 4704 2148 4760 2204
rect 4760 2148 4764 2204
rect 4700 2144 4764 2148
rect 4780 2204 4844 2208
rect 4780 2148 4784 2204
rect 4784 2148 4840 2204
rect 4840 2148 4844 2204
rect 4780 2144 4844 2148
rect 4860 2204 4924 2208
rect 4860 2148 4864 2204
rect 4864 2148 4920 2204
rect 4920 2148 4924 2204
rect 4860 2144 4924 2148
rect 4940 2204 5004 2208
rect 4940 2148 4944 2204
rect 4944 2148 5000 2204
rect 5000 2148 5004 2204
rect 4940 2144 5004 2148
rect 8448 2204 8512 2208
rect 8448 2148 8452 2204
rect 8452 2148 8508 2204
rect 8508 2148 8512 2204
rect 8448 2144 8512 2148
rect 8528 2204 8592 2208
rect 8528 2148 8532 2204
rect 8532 2148 8588 2204
rect 8588 2148 8592 2204
rect 8528 2144 8592 2148
rect 8608 2204 8672 2208
rect 8608 2148 8612 2204
rect 8612 2148 8668 2204
rect 8668 2148 8672 2204
rect 8608 2144 8672 2148
rect 8688 2204 8752 2208
rect 8688 2148 8692 2204
rect 8692 2148 8748 2204
rect 8748 2148 8752 2204
rect 8688 2144 8752 2148
rect 12196 2204 12260 2208
rect 12196 2148 12200 2204
rect 12200 2148 12256 2204
rect 12256 2148 12260 2204
rect 12196 2144 12260 2148
rect 12276 2204 12340 2208
rect 12276 2148 12280 2204
rect 12280 2148 12336 2204
rect 12336 2148 12340 2204
rect 12276 2144 12340 2148
rect 12356 2204 12420 2208
rect 12356 2148 12360 2204
rect 12360 2148 12416 2204
rect 12416 2148 12420 2204
rect 12356 2144 12420 2148
rect 12436 2204 12500 2208
rect 12436 2148 12440 2204
rect 12440 2148 12496 2204
rect 12496 2148 12500 2204
rect 12436 2144 12500 2148
rect 1900 444 1964 508
<< metal4 >>
rect 2818 16896 3138 17456
rect 2818 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3138 16896
rect 2818 15808 3138 16832
rect 2818 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3138 15808
rect 1899 15332 1965 15333
rect 1899 15268 1900 15332
rect 1964 15268 1965 15332
rect 1899 15267 1965 15268
rect 1902 14381 1962 15267
rect 2818 14720 3138 15744
rect 2818 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3138 14720
rect 1899 14380 1965 14381
rect 1899 14316 1900 14380
rect 1964 14316 1965 14380
rect 1899 14315 1965 14316
rect 1902 509 1962 14315
rect 2818 13632 3138 14656
rect 4692 17440 5012 17456
rect 4692 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5012 17440
rect 4692 16352 5012 17376
rect 4692 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5012 16352
rect 4692 15264 5012 16288
rect 4692 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5012 15264
rect 4692 14176 5012 15200
rect 4692 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5012 14176
rect 3371 13836 3437 13837
rect 3371 13772 3372 13836
rect 3436 13772 3437 13836
rect 3371 13771 3437 13772
rect 2818 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3138 13632
rect 2818 12544 3138 13568
rect 2818 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3138 12544
rect 2818 11456 3138 12480
rect 3374 12450 3434 13771
rect 4692 13088 5012 14112
rect 4692 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5012 13088
rect 3374 12390 3618 12450
rect 2818 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3138 11456
rect 2818 10368 3138 11392
rect 3371 11388 3437 11389
rect 3371 11324 3372 11388
rect 3436 11324 3437 11388
rect 3371 11323 3437 11324
rect 2818 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3138 10368
rect 2818 9280 3138 10304
rect 3374 9621 3434 11323
rect 3371 9620 3437 9621
rect 3371 9556 3372 9620
rect 3436 9556 3437 9620
rect 3371 9555 3437 9556
rect 2818 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3138 9280
rect 2818 8192 3138 9216
rect 2818 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3138 8192
rect 2818 7104 3138 8128
rect 2818 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3138 7104
rect 2267 6628 2333 6629
rect 2267 6564 2268 6628
rect 2332 6564 2333 6628
rect 2267 6563 2333 6564
rect 2270 5133 2330 6563
rect 2635 6220 2701 6221
rect 2635 6156 2636 6220
rect 2700 6156 2701 6220
rect 2635 6155 2701 6156
rect 2267 5132 2333 5133
rect 2267 5068 2268 5132
rect 2332 5068 2333 5132
rect 2267 5067 2333 5068
rect 2638 4725 2698 6155
rect 2818 6016 3138 7040
rect 3558 6629 3618 12390
rect 3923 12204 3989 12205
rect 3923 12140 3924 12204
rect 3988 12140 3989 12204
rect 3923 12139 3989 12140
rect 3555 6628 3621 6629
rect 3555 6564 3556 6628
rect 3620 6564 3621 6628
rect 3555 6563 3621 6564
rect 2818 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3138 6016
rect 2818 4928 3138 5952
rect 2818 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3138 4928
rect 2635 4724 2701 4725
rect 2635 4660 2636 4724
rect 2700 4660 2701 4724
rect 2635 4659 2701 4660
rect 2818 3840 3138 4864
rect 2818 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3138 3840
rect 2818 2752 3138 3776
rect 2818 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3138 2752
rect 2818 2128 3138 2688
rect 3926 2413 3986 12139
rect 4692 12000 5012 13024
rect 4692 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5012 12000
rect 4692 10912 5012 11936
rect 4692 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5012 10912
rect 4692 9824 5012 10848
rect 4692 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5012 9824
rect 4692 8736 5012 9760
rect 4692 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5012 8736
rect 4692 7648 5012 8672
rect 4692 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5012 7648
rect 4692 6560 5012 7584
rect 4692 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5012 6560
rect 4692 5472 5012 6496
rect 4692 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5012 5472
rect 4692 4384 5012 5408
rect 4692 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5012 4384
rect 4692 3296 5012 4320
rect 6566 16896 6886 17456
rect 6566 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6886 16896
rect 6566 15808 6886 16832
rect 8440 17440 8760 17456
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 16352 8760 17376
rect 10314 16896 10634 17456
rect 12188 17440 12508 17456
rect 12188 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12508 17440
rect 10731 17236 10797 17237
rect 10731 17172 10732 17236
rect 10796 17172 10797 17236
rect 10731 17171 10797 17172
rect 10314 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10634 16896
rect 9443 16828 9509 16829
rect 9443 16764 9444 16828
rect 9508 16764 9509 16828
rect 9443 16763 9509 16764
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 7787 15876 7853 15877
rect 7787 15812 7788 15876
rect 7852 15812 7853 15876
rect 7787 15811 7853 15812
rect 6566 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6886 15808
rect 6566 14720 6886 15744
rect 7790 14789 7850 15811
rect 8440 15264 8760 16288
rect 8891 16012 8957 16013
rect 8891 15948 8892 16012
rect 8956 15948 8957 16012
rect 8891 15947 8957 15948
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 7787 14788 7853 14789
rect 7787 14724 7788 14788
rect 7852 14724 7853 14788
rect 7787 14723 7853 14724
rect 6566 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6886 14720
rect 6566 13632 6886 14656
rect 6566 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6886 13632
rect 6566 12544 6886 13568
rect 6566 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6886 12544
rect 6566 11456 6886 12480
rect 6566 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6886 11456
rect 6566 10368 6886 11392
rect 6566 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6886 10368
rect 6566 9280 6886 10304
rect 6566 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6886 9280
rect 6566 8192 6886 9216
rect 6566 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6886 8192
rect 6566 7104 6886 8128
rect 6566 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6886 7104
rect 6566 6016 6886 7040
rect 6566 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6886 6016
rect 6566 4928 6886 5952
rect 6566 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6886 4928
rect 5579 4316 5645 4317
rect 5579 4252 5580 4316
rect 5644 4252 5645 4316
rect 5579 4251 5645 4252
rect 5582 3365 5642 4251
rect 6566 3840 6886 4864
rect 6566 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6886 3840
rect 5579 3364 5645 3365
rect 5579 3300 5580 3364
rect 5644 3300 5645 3364
rect 5579 3299 5645 3300
rect 4692 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5012 3296
rect 3923 2412 3989 2413
rect 3923 2348 3924 2412
rect 3988 2348 3989 2412
rect 3923 2347 3989 2348
rect 4692 2208 5012 3232
rect 4692 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5012 2208
rect 4692 2128 5012 2144
rect 6566 2752 6886 3776
rect 8440 14176 8760 15200
rect 8894 14517 8954 15947
rect 9446 15741 9506 16763
rect 9627 16556 9693 16557
rect 9627 16492 9628 16556
rect 9692 16492 9693 16556
rect 9627 16491 9693 16492
rect 9443 15740 9509 15741
rect 9443 15676 9444 15740
rect 9508 15676 9509 15740
rect 9443 15675 9509 15676
rect 8891 14516 8957 14517
rect 8891 14452 8892 14516
rect 8956 14452 8957 14516
rect 8891 14451 8957 14452
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 13088 8760 14112
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 12000 8760 13024
rect 9446 12749 9506 15675
rect 9443 12748 9509 12749
rect 9443 12684 9444 12748
rect 9508 12684 9509 12748
rect 9443 12683 9509 12684
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 10912 8760 11936
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 9824 8760 10848
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 8736 8760 9760
rect 9630 8941 9690 16491
rect 10179 16012 10245 16013
rect 10179 15948 10180 16012
rect 10244 15948 10245 16012
rect 10179 15947 10245 15948
rect 9995 14244 10061 14245
rect 9995 14180 9996 14244
rect 10060 14180 10061 14244
rect 9995 14179 10061 14180
rect 9627 8940 9693 8941
rect 9627 8876 9628 8940
rect 9692 8876 9693 8940
rect 9627 8875 9693 8876
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 7648 8760 8672
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 6560 8760 7584
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 5472 8760 6496
rect 9998 6221 10058 14179
rect 10182 12205 10242 15947
rect 10314 15808 10634 16832
rect 10314 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10634 15808
rect 10314 14720 10634 15744
rect 10314 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10634 14720
rect 10314 13632 10634 14656
rect 10314 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10634 13632
rect 10314 12544 10634 13568
rect 10734 13021 10794 17171
rect 10915 16964 10981 16965
rect 10915 16900 10916 16964
rect 10980 16900 10981 16964
rect 10915 16899 10981 16900
rect 10918 14109 10978 16899
rect 11835 16692 11901 16693
rect 11835 16628 11836 16692
rect 11900 16628 11901 16692
rect 11835 16627 11901 16628
rect 10915 14108 10981 14109
rect 10915 14044 10916 14108
rect 10980 14044 10981 14108
rect 10915 14043 10981 14044
rect 10731 13020 10797 13021
rect 10731 12956 10732 13020
rect 10796 12956 10797 13020
rect 10731 12955 10797 12956
rect 10734 12613 10794 12955
rect 10731 12612 10797 12613
rect 10731 12548 10732 12612
rect 10796 12548 10797 12612
rect 10731 12547 10797 12548
rect 10314 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10634 12544
rect 10179 12204 10245 12205
rect 10179 12140 10180 12204
rect 10244 12140 10245 12204
rect 10179 12139 10245 12140
rect 10314 11456 10634 12480
rect 11838 12450 11898 16627
rect 12188 16352 12508 17376
rect 13859 17100 13925 17101
rect 13859 17036 13860 17100
rect 13924 17036 13925 17100
rect 13859 17035 13925 17036
rect 12571 16692 12637 16693
rect 12571 16628 12572 16692
rect 12636 16628 12637 16692
rect 12571 16627 12637 16628
rect 13491 16692 13557 16693
rect 13491 16628 13492 16692
rect 13556 16628 13557 16692
rect 13491 16627 13557 16628
rect 12188 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12508 16352
rect 12188 15264 12508 16288
rect 12188 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12508 15264
rect 12188 14176 12508 15200
rect 12188 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12508 14176
rect 12188 13088 12508 14112
rect 12188 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12508 13088
rect 12019 12748 12085 12749
rect 12019 12684 12020 12748
rect 12084 12684 12085 12748
rect 12019 12683 12085 12684
rect 10314 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10634 11456
rect 10314 10368 10634 11392
rect 10314 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10634 10368
rect 10314 9280 10634 10304
rect 11654 12390 11898 12450
rect 11283 10028 11349 10029
rect 11283 9964 11284 10028
rect 11348 9964 11349 10028
rect 11283 9963 11349 9964
rect 10314 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10634 9280
rect 10314 8192 10634 9216
rect 10314 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10634 8192
rect 10314 7104 10634 8128
rect 10314 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10634 7104
rect 9995 6220 10061 6221
rect 9995 6156 9996 6220
rect 10060 6156 10061 6220
rect 9995 6155 10061 6156
rect 10314 6016 10634 7040
rect 10314 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10634 6016
rect 9995 5676 10061 5677
rect 9995 5612 9996 5676
rect 10060 5612 10061 5676
rect 9995 5611 10061 5612
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 4384 8760 5408
rect 9811 4860 9877 4861
rect 9811 4796 9812 4860
rect 9876 4796 9877 4860
rect 9811 4795 9877 4796
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 7235 3636 7301 3637
rect 7235 3572 7236 3636
rect 7300 3572 7301 3636
rect 7235 3571 7301 3572
rect 7238 2957 7298 3571
rect 8440 3296 8760 4320
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 7235 2956 7301 2957
rect 7235 2892 7236 2956
rect 7300 2892 7301 2956
rect 7235 2891 7301 2892
rect 6566 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6886 2752
rect 6566 2128 6886 2688
rect 8440 2208 8760 3232
rect 9814 3229 9874 4795
rect 9998 4045 10058 5611
rect 10179 5540 10245 5541
rect 10179 5476 10180 5540
rect 10244 5476 10245 5540
rect 10179 5475 10245 5476
rect 9995 4044 10061 4045
rect 9995 3980 9996 4044
rect 10060 3980 10061 4044
rect 9995 3979 10061 3980
rect 9811 3228 9877 3229
rect 9811 3164 9812 3228
rect 9876 3164 9877 3228
rect 9811 3163 9877 3164
rect 10182 2821 10242 5475
rect 10314 4928 10634 5952
rect 10915 5404 10981 5405
rect 10915 5340 10916 5404
rect 10980 5340 10981 5404
rect 10915 5339 10981 5340
rect 10314 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10634 4928
rect 10314 3840 10634 4864
rect 10314 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10634 3840
rect 10179 2820 10245 2821
rect 10179 2756 10180 2820
rect 10244 2756 10245 2820
rect 10179 2755 10245 2756
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2128 8760 2144
rect 10314 2752 10634 3776
rect 10918 3229 10978 5339
rect 11099 4452 11165 4453
rect 11099 4388 11100 4452
rect 11164 4388 11165 4452
rect 11099 4387 11165 4388
rect 11102 3773 11162 4387
rect 11286 4317 11346 9963
rect 11654 6357 11714 12390
rect 11651 6356 11717 6357
rect 11651 6292 11652 6356
rect 11716 6292 11717 6356
rect 11651 6291 11717 6292
rect 11283 4316 11349 4317
rect 11283 4252 11284 4316
rect 11348 4252 11349 4316
rect 11283 4251 11349 4252
rect 11099 3772 11165 3773
rect 11099 3708 11100 3772
rect 11164 3708 11165 3772
rect 11099 3707 11165 3708
rect 10915 3228 10981 3229
rect 10915 3164 10916 3228
rect 10980 3164 10981 3228
rect 10915 3163 10981 3164
rect 11654 3093 11714 6291
rect 12022 4045 12082 12683
rect 12188 12000 12508 13024
rect 12188 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12508 12000
rect 12188 10912 12508 11936
rect 12188 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12508 10912
rect 12188 9824 12508 10848
rect 12188 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12508 9824
rect 12188 8736 12508 9760
rect 12574 9077 12634 16627
rect 12939 15060 13005 15061
rect 12939 14996 12940 15060
rect 13004 14996 13005 15060
rect 12939 14995 13005 14996
rect 12942 11933 13002 14995
rect 13123 12884 13189 12885
rect 13123 12820 13124 12884
rect 13188 12820 13189 12884
rect 13123 12819 13189 12820
rect 12939 11932 13005 11933
rect 12939 11868 12940 11932
rect 13004 11868 13005 11932
rect 12939 11867 13005 11868
rect 12571 9076 12637 9077
rect 12571 9012 12572 9076
rect 12636 9012 12637 9076
rect 12571 9011 12637 9012
rect 12188 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12508 8736
rect 12188 7648 12508 8672
rect 12188 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12508 7648
rect 12188 6560 12508 7584
rect 13126 6765 13186 12819
rect 13494 9757 13554 16627
rect 13675 14788 13741 14789
rect 13675 14724 13676 14788
rect 13740 14724 13741 14788
rect 13675 14723 13741 14724
rect 13678 12341 13738 14723
rect 13675 12340 13741 12341
rect 13675 12276 13676 12340
rect 13740 12276 13741 12340
rect 13675 12275 13741 12276
rect 13675 12068 13741 12069
rect 13675 12004 13676 12068
rect 13740 12004 13741 12068
rect 13675 12003 13741 12004
rect 13491 9756 13557 9757
rect 13491 9692 13492 9756
rect 13556 9692 13557 9756
rect 13491 9691 13557 9692
rect 13123 6764 13189 6765
rect 13123 6700 13124 6764
rect 13188 6700 13189 6764
rect 13123 6699 13189 6700
rect 12188 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12508 6560
rect 12188 5472 12508 6496
rect 12571 5812 12637 5813
rect 12571 5748 12572 5812
rect 12636 5748 12637 5812
rect 12571 5747 12637 5748
rect 12188 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12508 5472
rect 12188 4384 12508 5408
rect 12574 4997 12634 5747
rect 12571 4996 12637 4997
rect 12571 4932 12572 4996
rect 12636 4932 12637 4996
rect 12571 4931 12637 4932
rect 12188 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12508 4384
rect 12019 4044 12085 4045
rect 12019 3980 12020 4044
rect 12084 3980 12085 4044
rect 12019 3979 12085 3980
rect 12188 3296 12508 4320
rect 12188 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12508 3296
rect 11651 3092 11717 3093
rect 11651 3028 11652 3092
rect 11716 3028 11717 3092
rect 11651 3027 11717 3028
rect 10314 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10634 2752
rect 10314 2128 10634 2688
rect 12188 2208 12508 3232
rect 13678 2549 13738 12003
rect 13862 11933 13922 17035
rect 14062 16896 14382 17456
rect 14062 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14382 16896
rect 14062 15808 14382 16832
rect 14779 16692 14845 16693
rect 14779 16628 14780 16692
rect 14844 16628 14845 16692
rect 14779 16627 14845 16628
rect 14062 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14382 15808
rect 14062 14720 14382 15744
rect 14595 15332 14661 15333
rect 14595 15268 14596 15332
rect 14660 15268 14661 15332
rect 14595 15267 14661 15268
rect 14062 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14382 14720
rect 14062 13632 14382 14656
rect 14062 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14382 13632
rect 14062 12544 14382 13568
rect 14062 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14382 12544
rect 13859 11932 13925 11933
rect 13859 11868 13860 11932
rect 13924 11868 13925 11932
rect 13859 11867 13925 11868
rect 14062 11456 14382 12480
rect 14062 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14382 11456
rect 13859 11116 13925 11117
rect 13859 11052 13860 11116
rect 13924 11052 13925 11116
rect 13859 11051 13925 11052
rect 13862 9485 13922 11051
rect 14062 10368 14382 11392
rect 14062 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14382 10368
rect 13859 9484 13925 9485
rect 13859 9420 13860 9484
rect 13924 9420 13925 9484
rect 13859 9419 13925 9420
rect 14062 9280 14382 10304
rect 14062 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14382 9280
rect 14062 8192 14382 9216
rect 14062 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14382 8192
rect 14062 7104 14382 8128
rect 14062 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14382 7104
rect 13859 6220 13925 6221
rect 13859 6156 13860 6220
rect 13924 6156 13925 6220
rect 13859 6155 13925 6156
rect 13862 2957 13922 6155
rect 14062 6016 14382 7040
rect 14062 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14382 6016
rect 14062 4928 14382 5952
rect 14598 5541 14658 15267
rect 14782 13021 14842 16627
rect 15147 14244 15213 14245
rect 15147 14180 15148 14244
rect 15212 14180 15213 14244
rect 15147 14179 15213 14180
rect 14963 13156 15029 13157
rect 14963 13092 14964 13156
rect 15028 13092 15029 13156
rect 14963 13091 15029 13092
rect 14779 13020 14845 13021
rect 14779 12956 14780 13020
rect 14844 12956 14845 13020
rect 14779 12955 14845 12956
rect 14779 5812 14845 5813
rect 14779 5748 14780 5812
rect 14844 5748 14845 5812
rect 14779 5747 14845 5748
rect 14595 5540 14661 5541
rect 14595 5476 14596 5540
rect 14660 5476 14661 5540
rect 14595 5475 14661 5476
rect 14062 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14382 4928
rect 14062 3840 14382 4864
rect 14598 4453 14658 5475
rect 14595 4452 14661 4453
rect 14595 4388 14596 4452
rect 14660 4388 14661 4452
rect 14595 4387 14661 4388
rect 14782 4045 14842 5747
rect 14966 5405 15026 13091
rect 15150 11117 15210 14179
rect 15147 11116 15213 11117
rect 15147 11052 15148 11116
rect 15212 11052 15213 11116
rect 15147 11051 15213 11052
rect 14963 5404 15029 5405
rect 14963 5340 14964 5404
rect 15028 5340 15029 5404
rect 14963 5339 15029 5340
rect 14779 4044 14845 4045
rect 14779 3980 14780 4044
rect 14844 3980 14845 4044
rect 14779 3979 14845 3980
rect 14062 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14382 3840
rect 13859 2956 13925 2957
rect 13859 2892 13860 2956
rect 13924 2892 13925 2956
rect 13859 2891 13925 2892
rect 14062 2752 14382 3776
rect 14062 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14382 2752
rect 13675 2548 13741 2549
rect 13675 2484 13676 2548
rect 13740 2484 13741 2548
rect 13675 2483 13741 2484
rect 12188 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12508 2208
rect 12188 2128 12508 2144
rect 14062 2128 14382 2688
rect 1899 508 1965 509
rect 1899 444 1900 508
rect 1964 444 1965 508
rect 1899 443 1965 444
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 1656 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1649977179
transform -1 0 1840 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1649977179
transform -1 0 2392 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1649977179
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1649977179
transform -1 0 2208 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1649977179
transform -1 0 2024 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1649977179
transform -1 0 2576 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1649977179
transform -1 0 4416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1649977179
transform 1 0 6716 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1649977179
transform 1 0 8004 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1649977179
transform -1 0 1932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1649977179
transform 1 0 5796 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1649977179
transform 1 0 7636 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1649977179
transform 1 0 15272 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1649977179
transform -1 0 2576 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1649977179
transform 1 0 2576 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1649977179
transform 1 0 3956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1649977179
transform -1 0 2484 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1649977179
transform 1 0 2760 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1649977179
transform 1 0 3036 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1649977179
transform 1 0 3128 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1649977179
transform -1 0 9108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1649977179
transform -1 0 3036 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1649977179
transform 1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1649977179
transform -1 0 3404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1649977179
transform 1 0 3312 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1649977179
transform 1 0 9200 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1649977179
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1649977179
transform 1 0 2116 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 3772 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 2392 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 9384 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 13616 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 12880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 14260 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 15180 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 14904 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 14444 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 15548 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 15088 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 15732 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 13984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 8832 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 11408 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 10856 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 11040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 10764 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 12328 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 12512 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 7084 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 13984 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 15456 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 15088 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 14720 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 14904 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 15548 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 15732 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 15364 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 15272 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 9568 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 4600 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 9660 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 9476 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 11040 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 13984 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 15732 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 12880 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 13340 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 15732 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_A
timestamp 1649977179
transform 1 0 15088 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7912 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6992 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9752 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 5704 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5336 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5704 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 7084 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5980 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 4140 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11776 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 7268 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 7268 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 6532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7912 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9108 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10580 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 12052 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9844 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8740 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10396 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 12512 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9936 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9384 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5520 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5336 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5888 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 4508 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 5520 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5336 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 5060 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 9660 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12972 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9752 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 6532 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 5428 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 4508 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 6716 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 7176 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12788 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11040 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 9292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 5704 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 5704 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7820 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 7636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 10764 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 10948 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 10672 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3864 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 3680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 4048 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5612 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 3956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 2576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 2208 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 2576 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 4048 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 2668 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 2852 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 2484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 2576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 12696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 12144 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 14260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 14996 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 15364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 7728 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 3680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 7452 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 6256 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14352 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 15548 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 10856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14168 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 14536 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 15088 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 15088 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 2944 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4048 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4232 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 4324 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3864 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 2668 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 2392 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3128 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3312 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4324 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4140 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 2944 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 12144 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 10672 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 11408 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 10488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 10672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 13340 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4048 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 4048 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12696 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9936 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 7912 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 7544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8464 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 9108 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 5520 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output45_A
timestamp 1649977179
transform 1 0 14536 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_N_FTB01_A
timestamp 1649977179
transform 1 0 15272 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_S_FTB01_A
timestamp 1649977179
transform -1 0 15640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater108_A
timestamp 1649977179
transform 1 0 9568 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater112_A
timestamp 1649977179
transform -1 0 10212 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater118_A
timestamp 1649977179
transform -1 0 10580 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater122_A
timestamp 1649977179
transform -1 0 9568 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_151
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_158
timestamp 1649977179
transform 1 0 15640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_37
timestamp 1649977179
transform 1 0 4508 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_145
timestamp 1649977179
transform 1 0 14444 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_52
timestamp 1649977179
transform 1 0 5888 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_129
timestamp 1649977179
transform 1 0 12972 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_61
timestamp 1649977179
transform 1 0 6716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_80
timestamp 1649977179
transform 1 0 8464 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_99
timestamp 1649977179
transform 1 0 10212 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_144
timestamp 1649977179
transform 1 0 14352 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_7
timestamp 1649977179
transform 1 0 1748 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_48
timestamp 1649977179
transform 1 0 5520 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_158
timestamp 1649977179
transform 1 0 15640 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_16
timestamp 1649977179
transform 1 0 2576 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_35
timestamp 1649977179
transform 1 0 4324 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_115
timestamp 1649977179
transform 1 0 11684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_155
timestamp 1649977179
transform 1 0 15364 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_79
timestamp 1649977179
transform 1 0 8372 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1649977179
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_126
timestamp 1649977179
transform 1 0 12696 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_143
timestamp 1649977179
transform 1 0 14260 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_158
timestamp 1649977179
transform 1 0 15640 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_63
timestamp 1649977179
transform 1 0 6900 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_98
timestamp 1649977179
transform 1 0 10120 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_106 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10856 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_115
timestamp 1649977179
transform 1 0 11684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_32
timestamp 1649977179
transform 1 0 4048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_49
timestamp 1649977179
transform 1 0 5612 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_87 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9108 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_99
timestamp 1649977179
transform 1 0 10212 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_34
timestamp 1649977179
transform 1 0 4232 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_147
timestamp 1649977179
transform 1 0 14628 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_10
timestamp 1649977179
transform 1 0 2024 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_64
timestamp 1649977179
transform 1 0 6992 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_154
timestamp 1649977179
transform 1 0 15272 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_49
timestamp 1649977179
transform 1 0 5612 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_115 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_121
timestamp 1649977179
transform 1 0 12236 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_129
timestamp 1649977179
transform 1 0 12972 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_139
timestamp 1649977179
transform 1 0 13892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_143
timestamp 1649977179
transform 1 0 14260 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_153
timestamp 1649977179
transform 1 0 15180 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_158
timestamp 1649977179
transform 1 0 15640 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_35
timestamp 1649977179
transform 1 0 4324 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_68
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1649977179
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp 1649977179
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_92
timestamp 1649977179
transform 1 0 9568 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_10
timestamp 1649977179
transform 1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_22
timestamp 1649977179
transform 1 0 3128 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_52
timestamp 1649977179
transform 1 0 5888 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_108
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_129
timestamp 1649977179
transform 1 0 12972 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_140
timestamp 1649977179
transform 1 0 13984 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_157
timestamp 1649977179
transform 1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_19
timestamp 1649977179
transform 1 0 2852 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_22
timestamp 1649977179
transform 1 0 3128 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_93
timestamp 1649977179
transform 1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_114
timestamp 1649977179
transform 1 0 11592 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_122
timestamp 1649977179
transform 1 0 12328 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_134
timestamp 1649977179
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1649977179
transform 1 0 14444 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1649977179
transform 1 0 1748 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_76
timestamp 1649977179
transform 1 0 8096 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_82
timestamp 1649977179
transform 1 0 8648 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_103
timestamp 1649977179
transform 1 0 10580 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_126
timestamp 1649977179
transform 1 0 12696 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_136
timestamp 1649977179
transform 1 0 13616 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_148
timestamp 1649977179
transform 1 0 14720 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_156
timestamp 1649977179
transform 1 0 15456 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_7
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_135
timestamp 1649977179
transform 1 0 13524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_156
timestamp 1649977179
transform 1 0 15456 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_10
timestamp 1649977179
transform 1 0 2024 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_29
timestamp 1649977179
transform 1 0 3772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_65
timestamp 1649977179
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_68
timestamp 1649977179
transform 1 0 7360 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_80
timestamp 1649977179
transform 1 0 8464 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_88
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1649977179
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_128
timestamp 1649977179
transform 1 0 12880 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_156
timestamp 1649977179
transform 1 0 15456 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_14
timestamp 1649977179
transform 1 0 2392 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_45
timestamp 1649977179
transform 1 0 5244 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_48
timestamp 1649977179
transform 1 0 5520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_56
timestamp 1649977179
transform 1 0 6256 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_81
timestamp 1649977179
transform 1 0 8556 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_101
timestamp 1649977179
transform 1 0 10396 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_105
timestamp 1649977179
transform 1 0 10764 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_126
timestamp 1649977179
transform 1 0 12696 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_11
timestamp 1649977179
transform 1 0 2116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_23
timestamp 1649977179
transform 1 0 3220 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_65
timestamp 1649977179
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_133
timestamp 1649977179
transform 1 0 13340 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_152
timestamp 1649977179
transform 1 0 15088 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_46
timestamp 1649977179
transform 1 0 5336 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_7
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_26
timestamp 1649977179
transform 1 0 3496 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_29
timestamp 1649977179
transform 1 0 3772 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_73
timestamp 1649977179
transform 1 0 7820 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_10
timestamp 1649977179
transform 1 0 2024 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_100
timestamp 1649977179
transform 1 0 10304 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_142
timestamp 1649977179
transform 1 0 14168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_18
timestamp 1649977179
transform 1 0 2760 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_32
timestamp 1649977179
transform 1 0 4048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_45
timestamp 1649977179
transform 1 0 5244 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_17
timestamp 1649977179
transform 1 0 2668 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_21
timestamp 1649977179
transform 1 0 3036 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_29
timestamp 1649977179
transform 1 0 3772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_92
timestamp 1649977179
transform 1 0 9568 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_158
timestamp 1649977179
transform 1 0 15640 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_79
timestamp 1649977179
transform 1 0 8372 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_151
timestamp 1649977179
transform 1 0 14996 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_158
timestamp 1649977179
transform 1 0 15640 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 16008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 16008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 16008 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 16008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 16008 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 16008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 16008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 16008 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 16008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 16008 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 16008 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 16008 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 16008 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 16008 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 16008 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _34_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1649977179
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1649977179
transform 1 0 1932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1649977179
transform 1 0 2208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1649977179
transform 1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1649977179
transform 1 0 3864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1649977179
transform -1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1649977179
transform -1 0 3128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1649977179
transform -1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1649977179
transform 1 0 4600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1649977179
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1649977179
transform 1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1649977179
transform -1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1649977179
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1649977179
transform 1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1649977179
transform -1 0 5704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1649977179
transform -1 0 6716 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1649977179
transform 1 0 11224 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1649977179
transform 1 0 7360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1649977179
transform 1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1649977179
transform 1 0 4140 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1649977179
transform 1 0 2576 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1649977179
transform 1 0 2852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1649977179
transform 1 0 4968 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1649977179
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1649977179
transform -1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1649977179
transform -1 0 3772 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1649977179
transform 1 0 4232 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1649977179
transform -1 0 4048 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1649977179
transform 1 0 13524 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1649977179
transform -1 0 4876 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1649977179
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1649977179
transform 1 0 5796 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1649977179
transform -1 0 5152 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1649977179
transform 1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1649977179
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1649977179
transform 1 0 2392 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 4048 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12880 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform 1 0 14904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1649977179
transform -1 0 14444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1649977179
transform 1 0 14444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1649977179
transform 1 0 14536 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1649977179
transform 1 0 14812 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1649977179
transform -1 0 15640 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1649977179
transform -1 0 15732 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1649977179
transform -1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1649977179
transform -1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1649977179
transform -1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1649977179
transform 1 0 10488 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform -1 0 11408 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1649977179
transform -1 0 10488 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1649977179
transform -1 0 12696 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1649977179
transform 1 0 11960 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 7452 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1649977179
transform -1 0 13708 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1649977179
transform -1 0 13524 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1649977179
transform -1 0 14996 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1649977179
transform -1 0 14444 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1649977179
transform -1 0 14812 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1649977179
transform -1 0 14628 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1649977179
transform 1 0 14812 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1649977179
transform -1 0 14536 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1649977179
transform -1 0 13984 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1649977179
transform -1 0 9568 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform -1 0 8832 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1649977179
transform -1 0 9476 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input37
timestamp 1649977179
transform 1 0 10304 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input38
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1649977179
transform 1 0 11040 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1649977179
transform -1 0 11040 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1649977179
transform 1 0 12420 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1649977179
transform -1 0 13064 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform -1 0 15732 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform -1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15732 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15732 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_2  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14996 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 13800 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7360 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4324 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8372 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7176 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 8648 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9752 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9936 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11960 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 5888 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 9660 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5336 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5704 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4140 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4416 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 5888 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8740 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 6992 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 5796 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4784 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4140 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4784 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13432 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 12696 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8832 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8924 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7268 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6716 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8096 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9292 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10764 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13708 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11500 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8924 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10580 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13524 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10120 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11040 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7360 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5336 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4416 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 6164 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 5520 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4784 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 3864 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4784 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7360 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10488 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7360 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9108 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9844 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13248 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8188 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7084 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 6164 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7360 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12788 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12696 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10948 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10396 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7912 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7912 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 5888 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8556 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform -1 0 7820 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8464 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9384 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_ipin_0.mux_l2_in_3__129 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10212 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 9844 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 9936 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15364 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11316 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform -1 0 10488 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10304 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10488 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 12880 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_0.mux_l2_in_3__130
timestamp 1649977179
transform -1 0 12052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12328 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10396 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 11500 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 9844 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3312 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2484 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_1.mux_l2_in_3__131
timestamp 1649977179
transform -1 0 2852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2760 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2300 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2484 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2024 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3496 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2668 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1649977179
transform -1 0 3404 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_2.mux_l2_in_3__138
timestamp 1649977179
transform -1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5152 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 3496 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1649977179
transform -1 0 3496 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2760 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3680 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3404 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5060 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2668 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4416 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_3.mux_l2_in_3__139
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 1840 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 1656 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2300 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12696 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12788 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1649977179
transform -1 0 12328 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12328 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 13524 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_4.mux_l2_in_3__123
timestamp 1649977179
transform 1 0 14536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12144 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 13156 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12052 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2300 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7360 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6532 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7820 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_5.mux_l2_in_3__124
timestamp 1649977179
transform -1 0 7360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 6808 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6164 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5428 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13800 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14904 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14536 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14720 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_6.mux_l2_in_3__125
timestamp 1649977179
transform 1 0 15088 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13708 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12972 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8924 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1649977179
transform -1 0 9752 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1649977179
transform -1 0 11408 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10580 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12788 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13340 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_7.mux_l2_in_3__126
timestamp 1649977179
transform -1 0 13984 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1649977179
transform -1 0 12512 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12788 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1649977179
transform 1 0 11868 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1472 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14352 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14444 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13800 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 13892 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14536 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_8.mux_l2_in_3__127
timestamp 1649977179
transform 1 0 15272 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14904 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14260 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12604 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3496 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2668 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2116 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2944 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_9.mux_l2_in_3__128
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2852 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 1840 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2024 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2392 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2392 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2300 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_10.mux_l2_in_3__132
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1649977179
transform 1 0 3128 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2852 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1649977179
transform -1 0 3588 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8648 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1649977179
transform 1 0 10212 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9108 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9936 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1649977179
transform -1 0 10304 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_11.mux_l2_in_3__133
timestamp 1649977179
transform -1 0 11040 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1649977179
transform -1 0 9936 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1649977179
transform 1 0 9660 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1649977179
transform 1 0 9476 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14904 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13156 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1649977179
transform -1 0 12328 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13800 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1649977179
transform -1 0 13708 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14260 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_12.mux_l2_in_3__134
timestamp 1649977179
transform 1 0 14904 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1649977179
transform -1 0 14168 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1649977179
transform -1 0 14260 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1472 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5888 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5060 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5336 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_13.mux_l2_in_3__135
timestamp 1649977179
transform -1 0 5796 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4416 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4508 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4140 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12328 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1649977179
transform -1 0 12696 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1649977179
transform -1 0 11408 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1649977179
transform -1 0 10948 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1649977179
transform -1 0 8280 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_14.mux_l2_in_3__136
timestamp 1649977179
transform 1 0 13248 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12328 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1649977179
transform -1 0 11776 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1649977179
transform 1 0 11040 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7360 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7268 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1649977179
transform -1 0 8004 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6532 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8004 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1649977179
transform 1 0 7728 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7544 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_15.mux_l2_in_3__137
timestamp 1649977179
transform -1 0 6348 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6348 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6716 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5888 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output45 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1649977179
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1649977179
transform -1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1649977179
transform 1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1649977179
transform 1 0 5704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1649977179
transform -1 0 6256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1649977179
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform 1 0 7176 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform -1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform -1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform -1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform 1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform -1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform 1 0 2944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform 1 0 4048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform -1 0 1840 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform 1 0 5152 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform -1 0 5152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform 1 0 5520 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform -1 0 5520 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 6808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 7176 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 7544 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform -1 0 8832 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 1840 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform -1 0 2208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform -1 0 2576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform -1 0 2944 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform -1 0 3312 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform 1 0 3312 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform 1 0 4048 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform 1 0 4048 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 4784 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform 1 0 15364 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform -1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform -1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform -1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform -1 0 2208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform 1 0 2208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform -1 0 2116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output104
timestamp 1649977179
transform -1 0 15456 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output105
timestamp 1649977179
transform -1 0 15732 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform 1 0 15364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15088 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1649977179
transform 1 0 15088 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater107
timestamp 1649977179
transform 1 0 14628 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater108
timestamp 1649977179
transform -1 0 11316 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater109
timestamp 1649977179
transform -1 0 3404 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater110
timestamp 1649977179
transform 1 0 8096 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater111
timestamp 1649977179
transform 1 0 14536 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater112
timestamp 1649977179
transform -1 0 10028 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater113
timestamp 1649977179
transform -1 0 4876 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater114
timestamp 1649977179
transform -1 0 5060 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater115
timestamp 1649977179
transform -1 0 4232 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater116
timestamp 1649977179
transform 1 0 8188 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater117
timestamp 1649977179
transform 1 0 13156 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater118
timestamp 1649977179
transform -1 0 10212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater119
timestamp 1649977179
transform -1 0 3036 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater120
timestamp 1649977179
transform 1 0 4232 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater121
timestamp 1649977179
transform 1 0 13064 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater122
timestamp 1649977179
transform -1 0 9108 0 -1 4352
box -38 -48 314 592
<< labels >>
flabel metal2 s 1030 19200 1086 20000 0 FreeSans 224 90 0 0 IO_ISOL_N
port 0 nsew signal input
flabel metal4 s 4692 2128 5012 17456 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 8440 2128 8760 17456 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 12188 2128 12508 17456 0 FreeSans 1920 90 0 0 VGND
port 1 nsew ground bidirectional
flabel metal4 s 2818 2128 3138 17456 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 6566 2128 6886 17456 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 10314 2128 10634 17456 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal4 s 14062 2128 14382 17456 0 FreeSans 1920 90 0 0 VPWR
port 2 nsew power bidirectional
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 ccff_head
port 3 nsew signal input
flabel metal3 s 16400 2048 17200 2168 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 5 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 6 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 7 nsew signal input
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 8 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 9 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 10 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 11 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 12 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 13 nsew signal input
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 14 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 15 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 16 nsew signal input
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 17 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 18 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 19 nsew signal input
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 20 nsew signal input
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 21 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 22 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 23 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 24 nsew signal input
flabel metal2 s 1214 0 1270 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 25 nsew signal tristate
flabel metal2 s 4894 0 4950 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 26 nsew signal tristate
flabel metal2 s 5262 0 5318 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 27 nsew signal tristate
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 28 nsew signal tristate
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 29 nsew signal tristate
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 30 nsew signal tristate
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 31 nsew signal tristate
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 32 nsew signal tristate
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 33 nsew signal tristate
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 34 nsew signal tristate
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 35 nsew signal tristate
flabel metal2 s 1582 0 1638 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 36 nsew signal tristate
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 37 nsew signal tristate
flabel metal2 s 2318 0 2374 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 38 nsew signal tristate
flabel metal2 s 2686 0 2742 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 39 nsew signal tristate
flabel metal2 s 3054 0 3110 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 40 nsew signal tristate
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 41 nsew signal tristate
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 42 nsew signal tristate
flabel metal2 s 4158 0 4214 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 43 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 44 nsew signal tristate
flabel metal2 s 8758 19200 8814 20000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 45 nsew signal input
flabel metal2 s 12438 19200 12494 20000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 46 nsew signal input
flabel metal2 s 12806 19200 12862 20000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 47 nsew signal input
flabel metal2 s 13174 19200 13230 20000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 48 nsew signal input
flabel metal2 s 13542 19200 13598 20000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 49 nsew signal input
flabel metal2 s 13910 19200 13966 20000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 50 nsew signal input
flabel metal2 s 14278 19200 14334 20000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 51 nsew signal input
flabel metal2 s 14646 19200 14702 20000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 52 nsew signal input
flabel metal2 s 15014 19200 15070 20000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 53 nsew signal input
flabel metal2 s 15382 19200 15438 20000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 54 nsew signal input
flabel metal2 s 15750 19200 15806 20000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 55 nsew signal input
flabel metal2 s 9126 19200 9182 20000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 56 nsew signal input
flabel metal2 s 9494 19200 9550 20000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 57 nsew signal input
flabel metal2 s 9862 19200 9918 20000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 58 nsew signal input
flabel metal2 s 10230 19200 10286 20000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 59 nsew signal input
flabel metal2 s 10598 19200 10654 20000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 60 nsew signal input
flabel metal2 s 10966 19200 11022 20000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 61 nsew signal input
flabel metal2 s 11334 19200 11390 20000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 62 nsew signal input
flabel metal2 s 11702 19200 11758 20000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 63 nsew signal input
flabel metal2 s 12070 19200 12126 20000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 64 nsew signal input
flabel metal2 s 1398 19200 1454 20000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 65 nsew signal tristate
flabel metal2 s 5078 19200 5134 20000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 66 nsew signal tristate
flabel metal2 s 5446 19200 5502 20000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 67 nsew signal tristate
flabel metal2 s 5814 19200 5870 20000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 68 nsew signal tristate
flabel metal2 s 6182 19200 6238 20000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 69 nsew signal tristate
flabel metal2 s 6550 19200 6606 20000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 70 nsew signal tristate
flabel metal2 s 6918 19200 6974 20000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 71 nsew signal tristate
flabel metal2 s 7286 19200 7342 20000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 72 nsew signal tristate
flabel metal2 s 7654 19200 7710 20000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 73 nsew signal tristate
flabel metal2 s 8022 19200 8078 20000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 74 nsew signal tristate
flabel metal2 s 8390 19200 8446 20000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 75 nsew signal tristate
flabel metal2 s 1766 19200 1822 20000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 76 nsew signal tristate
flabel metal2 s 2134 19200 2190 20000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 77 nsew signal tristate
flabel metal2 s 2502 19200 2558 20000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 78 nsew signal tristate
flabel metal2 s 2870 19200 2926 20000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 79 nsew signal tristate
flabel metal2 s 3238 19200 3294 20000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 80 nsew signal tristate
flabel metal2 s 3606 19200 3662 20000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 81 nsew signal tristate
flabel metal2 s 3974 19200 4030 20000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 82 nsew signal tristate
flabel metal2 s 4342 19200 4398 20000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 83 nsew signal tristate
flabel metal2 s 4710 19200 4766 20000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 84 nsew signal tristate
flabel metal3 s 16400 9936 17200 10056 0 FreeSans 480 0 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 85 nsew signal tristate
flabel metal3 s 16400 13880 17200 14000 0 FreeSans 480 0 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 86 nsew signal input
flabel metal3 s 16400 17824 17200 17944 0 FreeSans 480 0 0 0 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 87 nsew signal tristate
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 left_grid_pin_16_
port 88 nsew signal tristate
flabel metal3 s 0 4224 800 4344 0 FreeSans 480 0 0 0 left_grid_pin_17_
port 89 nsew signal tristate
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 left_grid_pin_18_
port 90 nsew signal tristate
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 left_grid_pin_19_
port 91 nsew signal tristate
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 left_grid_pin_20_
port 92 nsew signal tristate
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 left_grid_pin_21_
port 93 nsew signal tristate
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 left_grid_pin_22_
port 94 nsew signal tristate
flabel metal3 s 0 9936 800 10056 0 FreeSans 480 0 0 0 left_grid_pin_23_
port 95 nsew signal tristate
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 left_grid_pin_24_
port 96 nsew signal tristate
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 left_grid_pin_25_
port 97 nsew signal tristate
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 left_grid_pin_26_
port 98 nsew signal tristate
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 left_grid_pin_27_
port 99 nsew signal tristate
flabel metal3 s 0 14696 800 14816 0 FreeSans 480 0 0 0 left_grid_pin_28_
port 100 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 left_grid_pin_29_
port 101 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 left_grid_pin_30_
port 102 nsew signal tristate
flabel metal3 s 0 17552 800 17672 0 FreeSans 480 0 0 0 left_grid_pin_31_
port 103 nsew signal tristate
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 left_width_0_height_0__pin_0_
port 104 nsew signal input
flabel metal3 s 0 416 800 536 0 FreeSans 480 0 0 0 left_width_0_height_0__pin_1_lower
port 105 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 left_width_0_height_0__pin_1_upper
port 106 nsew signal tristate
flabel metal2 s 16118 19200 16174 20000 0 FreeSans 224 90 0 0 prog_clk_0_N_out
port 107 nsew signal tristate
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 prog_clk_0_S_out
port 108 nsew signal tristate
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 prog_clk_0_W_in
port 109 nsew signal input
flabel metal3 s 16400 5992 17200 6112 0 FreeSans 480 0 0 0 right_grid_pin_0_
port 110 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 17200 20000
<< end >>
